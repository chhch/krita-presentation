<!DOCTYPE html><html><head><meta charset="UTF-8"><title>Spice-Up - WebViewer</title><meta name="viewport" content="width=device-width, initial-scale=1"/></head><style>.slides{background-color: #363B3E;}html, body{background-color: #363B3E;}#content{display: none;}.slide{ background-color: lightgray; position: relative; overflow: hidden; margin-bottom: 16px; margin-left: auto; margin-right: auto; border: solid 1px #0E0F10; border-radius: 12px;}.slide-16-9{min-width: 1920px; max-width: 1920px; min-height: 1080px; max-height: 1080px;}.slide-16-10{min-width: 1920px; max-width: 1920px; min-height: 1200px; max-height: 1200px;}.slide-4-3{min-width: 1920px; max-width: 1920px; min-height: 1440px; max-height: 1440px;}.slide-3-2{min-width: 1920px; max-width: 1920px; min-height: 1280px; max-height: 1280px;}.slide-5-4{min-width: 1920px; max-width: 1920px; min-height: 1536px; max-height: 1536px;}.canvas-item{position: absolute; display: flex;}text-item{white-space: pre-wrap;}text-item span{align-self: center;}</style><script>if (!String.build){String.build=function (format){var args=Array.prototype.slice.call (arguments, 1); return format.replace (/{(\d+)}/g, function (match, number){return typeof args[number] !='undefined' ? args[number] : match;});};}function base64Decode(str){return decodeURIComponent(Array.prototype.map.call(atob(str), function(c){return '%' + ('00' + c.charCodeAt(0).toString(16)).slice(-2);}).join(''));}function makeIdEditable (id){get (id).contentEditable="true";}function get (id){return document.getElementById(id);}function downloadString (element, fileName, mime){var dlAnchorElem=document.getElementById ('download-anchor'); if (dlAnchorElem===null){document.getElementById ("body").innerHTML +='<a id="download-anchor" style="display:none"></a>'; dlAnchorElem=document.getElementById ('download-anchor');}var dataStr="data:" + mime + ";charset=utf-8," + encodeURIComponent(element); var dlAnchorElem=document.getElementById ('download-anchor'); dlAnchorElem.setAttribute ("href", dataStr); dlAnchorElem.setAttribute ("download", fileName); dlAnchorElem.click ();}</script><body id="body"> <h1 style="color: #dfdfdf; font-family: sans-serif; text-align: center; width: 100%; margin-top: 200px; font-size: 3em"> Loading presentation... </h1> <content id="content">
{"current-slide":8, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(to right, #3ab5b0 0%, #3D99BE 31%, #56317a 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/45-degree-fabric-dark.png" , "items": [{"x": -622,"y": 444,"w": 2791,"h": 472,"type":"text","text": "","text-data": "V2FydW0gaXN0IGRlciBIaW1tZWwgYmxhdT8=","font": "sacramento","color": "rgb(207, 227, 242)","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -615,"y": 771,"w": 2768,"h": 315,"type":"text","text": "","text-data": "IHZvbiBDaHJpc3RvcGggSGVsbG1pY2g=","font": "bad script","color": "rgb(49, 58, 89)","font-size": 16, "font-style":"regular", "justification": 1, "align": 1 }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nGy9Z7Bt13Em9vXa+9yXE4BHpAciEYEACZIASAiCmKNESh4FSiPJGiuMPfPHY1fZ/jfl8lT5h1OVPR5VuVxyacqasa0pqayRNBIlykoMIphBgCQCkTMIPDy8fO85e6/2j+6vu/fFXPLhhnPO3it0+PrrXr3lzv/8P/3D8dixj0EhECi6AtIAAaAq8C+dOkREAQAiEAUgDdo7oGp/E4H2DmkD0LtAGqB+ARHoPCsgkNbsuqr2+jAAEKDP0K4q0gSt2efmGTEYaaIKBSDSmqoqBCLaZxWIAAJVhQwjACh6R4xBBDptIOMoOs1AV417AEDvfh+BNBH7nWNUQBrvbP9UofMMkWb36B0QsWH0Of4m0uy9atcXaQAUvL4MI9C7raO9I64f/wC1xYXa2qvdq8+AjwoKoDUIAGiHqqiIL/M82a1VFH0WiNinoAKFqto47bMqqpprIqJQu719RqB9zrHaGyFogHaJscPerzpDFGqL6sNV9XXwtdKukEHsehprAeWed7XhNxsLINpnbZyIAiIDgK5dAe6qAJj7jCaDoM/otpH2eq4t5yK2R/4aFFBRlGvFfFxOqB8iAtUOUYHGWqhtF2VGbZ1yrC4T6lcTMTnw+djmQFRh+0hZtzHGnue+KGUBokDXDkEsKHUIUFcmW0dTelVTaIWN3+fNOQPATr/wl+N49OjHcMmx/dxcAKagrSi6+gdFgK7xN+UkhtFem2f7ORQcgBkOe59qKBHlHc0VTReKaZ/zn4UbKA1CQUIDlUGo6DRiscODjWva+LLY8sk053qXBVft9h6OwddCWjO5iEX3NRGBjFvQaYK05mujZrCoDNrNaJg2A/PG5uFGJK45T244x90CUATYxTrW0T8jza7jAie8fu/QeUJrA7SbkOu88XtzkVyg+xxjcmkCjYR29fGbCIt2SBt9ejOaDGFAbF2aK4LtuXAd/GeRlgZHe1kvM6TcA/E1jmtTSaFA1zBVdX0Gn5v2CYBgpdznGY1rGGOCr7/pWaOKaJHf+AzXSiBthPYJAp9nuaYpX4/r8t58re6rYjZ5RLPXWtxo8T4aUffmddIu126g3GgpOgb6FgUUE01kXh8KRUdDSwPlc+UcqrHQph8bZbXycdEbqCmwC154f/GNav69u7fh+4YhFd9QhAlUE7ORfg+dZxcov+esIQTaO2RwQZ5nu6a68gEAehoxBXSzNiWVIccwT65IMyD+/nl24+O/Q+13Ecg0xfxiM/l5n7s5viGBVuc4DCGYMfFB+e+8XoIzNwgUwlAu3w0RR2TFUAuVDHE/gwKzKXcojhs/dzrqxlMoFJyL/1XaaGhDU3Ag8e4werEu3HtHkHBjYGiEc3eUwHUNRequPFiOJxSJhgKmpOJOgm6ShtHHqn0DuHJxDGmoOpRORDvgihBC745Hdc650DBREWnUBBAMWHhcN2bgfcOQ9HQOoWycXyo3nVF8rhjOQJxcZ14HXIvOVxdyk6/PyzXmvnLPpdm8y1caEH4m1ypRo4LmbNR5RkBrwBScytD8li4MogAGX5S5mxISHewKG2Rc2SZPkxsRv0bLe5mAdWAYQxHS+Iyu8IN77erVuxmruKffA5KCNQw2RpUMc4bBjdAYBscM4OArZIZHoID6OtBwrLbMsEiDYuOWHPFZccOBcYwNT6WAzWsYct4KUw4PQ0RTSMK7yeiKOYPoSsM7uSARzYU3EBfw2HozQmpGRcaVjUsQa2VGiqGG2r4vIboJbu8+J+5jM2/YZ0eJPt6+CahtCsE917hOGAgwHOmADD5XKl5Vj0SdQkTGaxDh+udVW1xf4KjKnYXGntMx0BjCMH+gyw6R0RWsYpiUMfFfIQyj1Y2KxLiokMKpaEfjdaXOsYQwgghbQTEtK2JjG1ypK9LId4VhQ/d1WZiagiLNJFUDY8OKoJCGSkcREQwDdHaP6B8ShfMPtNQG4W2jczESSpcvKrZa7K7rNaT5PcYxPRfElGWe82+9l9ClzI/eYqZ3K8rFn+lhxzHRBJBexFFP8AptCEOVvAPSSPDa4ugkNko8lHJF83spDQaHPU+mQB6b8vNwyIg2mDH1EI5/S07AN6+5waL3Fsqd3Z8CLuSNZu5HQQ7a/doM2Sx0kV3hZq4Rvbkmaqr7oFjse/IMDHfWNk8aPcJ9X7NAOxHutLwuxcuEyQyfwte9GlSOKw2FEJn4nqumvBrl01LZJb18GAnQo1dU0FNtKUturGzeGp8y4zLkmrv8aVy9QXXKtfB9qwjEjEBbGK76IsM8cidLBFI304yGxvj5czV+METl1+E6pVDwTYpRoSq+uBpKC4d75gWIEGRrC5hnmzgVjBuxWTukKh6f3sQJU2n0XCb8OtNjIj1dL0JJIpHQvhEWJkQOgSE/Uf8RvtNzlYnHV0B0v9e8k8ZDGjCtfTzNCCxCRIewutmx920sxJDWcs2CS6CV9+80ZH3OOXCcjq6EhgGwuXHtnEPlXoYCgOvnyiEAQMMjvsRF0H0dyC3YOnNusHfPhkSgsy9z4WIA6LxJr55Wne7GX/M5O0Izg6rF9nBt4PN2geCeGHEJciZEP3XeoTQ0yDJAAl1V5Sn7r929tJGBodAi6H0yueWclDOiw5xSdgDbVxLYKPMNb64ZMmGOOSQ3xZUTIJCCJLe04OLIs5sDr9jDwkJB93CDe57iwv+6UQaRFsMwuDFxApbXtfvJCBUJS9waMLQSR7mXag1Ybdmgh8GEyoWHQkFWX0YnO3tBANUz9w6MLa5VMi/+Xl/oeQLGlVtZgLFkoAV6YnrCEupg2qQ34j1DETP+jayFzqaMMkD6Lk/XPKwAAqpTAU0uCetLKOaKb5C/O3np60voLoKA4BVKdhfSui7OtZiwFYEXQcJ5APNkGxzobDKlEL+GmlJlvM79a2bPKJFu7GR04o3sPXqgDJEGGcaA+AwvwtANNFQ07MnjRBhKUjaQn3MWVAoPTTN7QOjugRH3CK7AHFugIYQRyGWrnpXrR6jmisN9LAilendDMSV7BZ+fIkJm8gMCgYYRpDEpe24QMdE7EA4xQxKOlwaMBgnoQZ4rVJuHDBnC1GAmEQgdTnIylIUgYnMXDHACGDE0RWsGp6mktEC0arEA7hXIaUyuNK0Z9J+mICVD0Cm4laewFU9ewY2N0qPXEILvhbPl4QnzZSMv/drFS9PjRFjDa5E/8XvKOAbxml8FOSmSmHXy0tKRgzs/hjKDE4/wNBgMclMYKTDxfvFrrtLDB4lbvDNRDzeFHBINMREKSdCB6+1oRhWQ0W7fu98fzj/BQ4IydUHOm17euQRTAs11VQ2ei7DeQo2KLj3+FYlwwWzUCtI7tEkY7rQdkmIea1NFouVgNdFr/o40bJQL7sfusIf77WtqKVCiD1Na8XUKNLO4P0ORDtVqxOiZJZxUoAlyOlr9dyqshmIDi80J4tzTroE6Wux5zpe8AzkOM7w2vyXZGeMEsUuunb1XMWKzCSEKTkQ4KJeTacqFEXHewck8IgjVEv8XS0zvD5hwzbOhk2lapGh1vZOemYOYnfMggSbixsXGJMOYihV8gSOMWPsWApSGwjfJiVGdpgwL2oAIy0o9gbS8jkiDilpYRfK1jcGZGOREbmorghLK58aob6Boi0wCGAfTABavRygvwyquYzl+hEIwexMKpi4wQMxb2hjQOJx/lZzOzA0RjBuEll4V5GzU96SEkBmu+X4M9t14heZk6Xr3XYNTSbI2ZUn75Cij5R4uMgyKJOZyPRYK4EaJ6UxTpMxmqbIagzpAw90QLKUUOShcDACaFX8PjQSNnV1HI0wgUvA0ZyAE5NorjSVc4c2AEXVlZsXDB82sSVX6JI7zr8uVxy4DYiYyjaVoAwDdTAbDO9NcpnhKpaPxGIYQOHvPDNYRGElZQoMK5YYh/40rX/uWKULCeN+g4B+GMScyz0lAAmawoIaEyBEwqwEgOINdEJJEH7qPm8ZuZhza7V4EjrxGURIaEeWcuRb0EW5YFFaDIm0wpSJ64/i052YzXc15+H0tTVoISxqUMGbpxZXXbcbOa1GWQCrOfei8MWXxPRSuTcTZPv82xucVyXEo58xUOcnSokicsxfJmRdc1JcU7+xGXcoeLlOcPhYFVCcbh9eThGGK2pswF2GwJdY7DXEqel/ISAQNizRuEriINSjowfmCVC5mZMrchHUQObYkKQsXFPfbJYNlHIuQND5PI5BhS+5lvSbRKd+jcZ28lu76H2TEapXGYS6Lx8+6MjFTgkbvnvFihBRAcgj8GjKFZtmBoqiqhk5kTCEtwhFerY1GMBd4BUgxThrvjTRpHQsNBzSRyMh5Z5YjY8EyjkjbUvDMAJhBoafxNQhzLYC4Je9zTolCVmsxvLjJ5lZtvaO4QXJcXa0OhZsqS2UTVnCSH4q5I1KzIg06CDC5wtHw0WAED4S4rzivk56UNTYuoIyvXQgz5geydsKrVB2NSM1Ula8IRQUQHRzduhwAhuiYuaJqxLV8jUn+7SKWzdgQjeib7p2K73US5XXjDxi2SNkzwOJ+KlqqWc1kGKmYHAkpZygQBW8xbr88EV/RtUyJ0ji6+i8yJm5kfDTknSytzHXTFNeFcS3z9cwJjZuFIUMh3jQ9o33KNopZDiu2Eoexml59noBhBaiHF6stYCjKze9zd0iKpVHhRjexzytScBneNEcTg6cc22BkZsB3zXACjloCeu4yAt29SaCPVLzIQYewVDhuiMgQ6VjmBvPWzYvTPLcdvqIXWA2E0qjQ01WYTAPoayD+/soHVaNMpSjViIxbDfbnGAPJkTBlBT+NE2wpkrBsETqIDKYwUc6eWR0LfUbPeBUkBFYwVg6DS8CqXknnEcbKjTp5ERksDGnN+SJ6TDfyu9KLFY7TYBhKK8WEyLHkGrniSw0HmOWCza8YmqjOjHC3SEzsfxXyf1+Y1EOOzEjY+DLjo4vP5345wtP6SjH8dQW8XiQMvnMdkeFRGknnptxQECU1iI5og1iGgxa5QzcbYCgMt3txdQ+mfQZGAHO3eN+9GnTjpc8DsMm0mnlTNza0pCzqoSdpAKZctEAgcQ3PKogAOzu2KnQo5C8C3rqCLYqwfMHDEPZSnOWfY0jSEF4QgYiyWE20QTdMqQ5poNTSzyyfNkXx6zYzuAbLh9h/llODwhMeewrPzRJxnTbu4T074NwDIkvAazpqCdIzhRquKMISbVdOU8TRhuV7rX12OW6WbWge+rBKlk5inkwI5w3VxObiYSwdb6CRQApizoWfKRXAJuqJ/Pq8Lv7PjS8NcuQV/fp9CiJTqRB8R8vQYlEnUslzIJVGO1ilqn1T1L352BFhUNQglXCOSijiDoayuQgDSGqWLAY5FUcDLcIMKnM1DxyT5P572NgW72h5X2VYQqdq5CwzXjkeu2fXWUZx4iksHucwd0NWDDmG0eG3Kw4rNcm8DwN07ecO6AGJDlqDwLiCRYl4KXSKrEl4F0cXXkgUVZzjHgDzYtJmqHzje7kW/P4U3shbo3Aqzq+QpgiuxqC6rLaAccvmt5kQqVN6vJFxtEZ2hWy7WWozTBZ2IOcOmPITUkcZO8koeikTi8biq1rpGYgCyIyBzSs8NvklrgVDkZK9oDAR1ZD1lzYmmozQC8GJSBug09rf69wBc//SoK16XVtrJaLzvQoOAxKcGYk8GhERhmphKiL+j+tqqYsgj1H/FhJuV2BKk2EJoJ6xnCCysn8QAGbMgiPRTOWaDxgY05tRgJiKSq2ilEA6ZmDSCHE8ywpLor0BJGADJfM95FLqHONnhkEoa9iWSIdq4Qiie/WoYAj0QYTBD4zauwp5CE9livMY2jsWnIZu0jITbkdJdIc0q8uQCpFVk7zTDnRJZfXDp8aWD2EcFkw8YTe5Bj8UZhB4zNfpVcIoGAcjqz3JSxCv8YvvjSIqpEK15iUoHTzvwVg80sw0iGXjQGGvNQOSCK2K7gLxSANaBwnp2Gxn5FnxqMh7xinfYbTVmj3cmmeocNPLGRJl9JnKZkSZp1NhaEDGrQjTtBjxmDfrTNwgmQGgorBgyvhzng9BKBMAGZbXld3nFlxZZAB0KvUaHXF2hAiJ4/A1s/Ufl4pVN933PCtZJXYl0poRvo0I44uWCRFNOcr0LM/L1DCLPIPvo6rNXSlqEtuf4/QxLdKbWl5lBsf1Rbywyjm3eB1Z1SkuM/ka5YLlCR0No69gj/nQqAoamjRtUPVQQvw7wiqn50eB7+VrmtJz+alJWa0y3iZTvt5AN5vMHtD751ImYcWU7FAO6nCTKRjh2d1a81p+bXr+QBydxGJmLOr742fuonY7zu7jY8EZgAjXdNr4704aheFyCEiPNa3NwM1TKl8VjHp/aZBxa/cqx/sjlUuYzrH0uRwMkzB8LFSK/VyEhR4mMRQhQqlrxCxEjBflPgpWMjKNq2WfdJ7Q542tv/Zdc+eUbM8tk1IyRblBfnfPGgUKQXjJIO2Y8fD312vnjns2oiASGk5bkzzoRyNKebD1dIOtPT0+6M2TL7Ix2b9ELmEC873KMv3M+iHW0LdEl3rCUIVjqKjRdrE4FWT1pvpnI7wIpFYyPXCjuDBggg5L14/CEIKwdLZqRgUKsdiSdGwOU9UnsDu7IM2ITUJraZCmecDKPbTurBGnQhmasArTi7Jka8stInIctbhKseusCZxrGcpYhoD4wqpPxtycX1VgpgCjfsTDEsJpohSijKFkcuDGA4ZMLPNg3qkex9d5AomlmDthuPMJMo5maIh4CpMeShzVtC64zIYQifH9TInTIHIPyHXMc1QZCgvcIlzSNMgRsbiSDCu7N1pWiYoXVklD80yYeCpcp3WgmdhDZCggIlYRq+r2i3tQsgdgVqOkIFsDvIVAHM9nOplH8z3Dk5xF4SuYQYHEPSpktx4PbCtQwyoO3wv2iFL89TyV2xGHAXkPcU+v6tw738sjAICFMhwTVXcAayotQ2Ohkfq+iGdTVFm5QaMhQDkn0pU4BagZlqWR6TFeEUFLb+XCtrXHRhVpriSk0ATeOCZTpTQiDD2mCVGcZE1XMtxg6nDuUdeBGgfHYSQXFAUwOSLhv5LLB6FrNSD1Xxx37+FRAyHMxYM2q/9IVEBv5CGJC72RfL5ZHnJEzUWfo2YhyE3OhRAajLMl0ZWU+fC6AmDa8bFPebQ9EMVc+AbNfiJc40oeF9KuIjPLnJsRk3GVn0VBIGHEppQF95yJQsQRDPduyr3gF9c9PPgcpF9+rmT0+4w44VrXCMVLU9hrVsMJVBOf3PMkIEstjHMytiZYGnyGRqD3b7HnWWtiylQPm8V258T9kpVbyQNgUQjmn+o6xfpqkGg+74oKaIDLfbJmo6xjQWEZXpjRaI5mlsYkTAM6WJDIPe8YAREryvINYTzqsXxkBZrnvBuszJuFS7XblCri6K9X+6EMIapE6fkUKQgLxUEQaxhXvt693MM9/zAG2RbWuOTfAfFMguR7UIY0ew1Ea0boevoP4dmSewmCLzgSxDh5XD67hqUBICmsItY0RuwwUdSDUKh3ZyiEiKiH8SUyCUFnpoVewbMAtg5TCeN8HNGkx7MfLOypvEknx6A2Bp4d6BMWjgUI4Uzj7ZwCX5NSUwIYhyF5NmPRJAjkYLwPCrQ4f4Yg1nSHBiIQZxhaLmmPLUovjUQYFIAo+ipZAs4n5ulOkzLDMavzFBEKpGIzzathdBsyi1WqWwNlkPNhURmdi48ZXugV6KPseUlLdy/FZ3KI8kSj3OP0qcR8K7fBhRJHsohzJoCIHayPUlwAGVb4QosINLyUugx5SpK8Rpwr8bCie7qSSsrr1zCCBkncMMAzKwB09hiV2RN+Vg2CBqQcRkvzOj+hM2MxXwzWYHBxKznnyic86wJkZofzH0YLXfh6G/IMiXaoQ8CQSwi0ZeVeeH9mLYLtr96wQQoSEBqjVrJTnqYMgS3Ea6Qw/UBX8BOFZK7ZjxASlmnz+rFGCaMDaWidO8m/XUYe7J5F5TRDmF2zEGPJ1ULwLzRS4THLukUjnSB7p1AsnjMxL9Yj7AgEEd64GIBCuqIYqze9HmtTC9eWvIrplcTfefLVDLHGGi5Tm4JaNGZGU5bXhF9T4BkYR72RHdldqg6Q49GYdzliECue+yzFYNj7aSCKPIdR6jpiGPKsBye04Clc6LsrR5OsJYi+ERJnNmp2JJXEDQqtPw+QQYFZrTBJPWwJRGCka+9A430g6JuLiPMMNDzzBNUh0Q6hYTV8RalpBOPIe3h4SQOlkiELXFl6GqMkpVwYOzMAvj7Rl0Li/lZr4GsTkDgOX/t+kxCkZ7exaZ8M+RB5RdrUsz4U5vo5zovH+imQjmJM4FyI1AW6OxcgSCMNJKoYVhZ2RKYFQc6aUfATBaU+wYzCEHwOQ7JFeMTrADZPrx8xkbLuWOn9GArV9GkW8pEH0Ng9INLYbuSs9qPnISxwm0rKUZZjtENY/j6H+TzIVesywvgk2LHpBW/Bl7N0gMVVefpULSxxlJu9LRDhj3EeBS1UyOsyl4aQJ4hjYbjzoIEgM5RmhYbO1meUYbDR0DO7TYteE34yEV2QhVli61s5BNZWbDZWyQlk7BwuEW/OqhQCMg9QqZ0hmSbzuvFxQZy76D29usILlIYkJqmUCuMj5skJTZ8Pqz6lOQLhPLmBGhkX6d3XwzZEPXZlhypBs/Jp997C1nI8vg560CJ8IoBDaqXxkGaIQj0EI0pzyx88j8fhrGbM8mrJcCjCuQERLtFnxSldBH8hoPF1QwKFNs37S/HcVDj2PegbqzegEUaDdIpwet0QUamp5znHUmFz9W/SHPiU+oHiZaPcXIoSNz8+Hx27EByFhSNTePPgB9yDi2dfloroghYh2ADr80FjmMf531yta/8R8c/Rg1PhmZP19GclXwMNKms53HBE7UVFAL6//poEesjOYfU8i62Wjz/G4M4p0AZinUcAots7fjALwOTMODkDhSmgainVpkL6P3Zm6j2ITxlZDl6Uj0Im4kjPPQWb7pAA4tFvRzcKWLgAIhSULISCdRDQnhkOepyhlIRPVpka8+GCi1g3r9WWoRQuNrAonNLIFLjgzcWjUgmL0alnIepXlPHS+LLxrnJ+LsRe8BSpRe0ZVqmWsMCFvKWSmdeZoYEMnQsgMbtZl7XSHFPM30k8ZaVkOTvi86Pw2dgkMw0hkAxp5E3zj0OIjqKCB6EBRIHdfgaCNRZZz9IK7wEwVWmobvJx+0lVtrwjmhJB7xs0WS1CNnUUl6islblk42M4CR4ZEPgap5YHQjA7VMIpKi0NQCimQlnRWkKPHEMlV8ljZJjNkIuRLN9jCIEZGVZ/8jMNHTPqWRmNa1WcARl1mhRDaQ8W6b05lCGQwejcwMa96LjKJjT0msyaMHUKrrX4DNTGFO3RaER82VhsQsXwgiO0tOpxBL3VxXSvO238tKpkKAU4mVk8RRV6cb5kntwwMXxw4+ZpyDB+PA9BRdndvJjTcr5HAQi9RnANFCgtawywb4gMqxxbqJmTfIX1D7KQ7w3F0RB4VRp1hg+9ZJ80x+21AQvSsQ123z75fMeExHaj3FuGngFzke/holRZCNShMeY4rcr7xzV67gfUOR03iG4YxPecSqt+QtRuz7QmInyNnp28viLmbqjDkVN48iSjOQ0gsxr8yqrUsueqYFUnlTGRB1s0lhaM4uu1WAeX/7hveSwBgHqqNIAjaNzUP5OoxT4zu0Ee4y+1QY/G74pRhiH6Uug026nGZp4dXsoMscpMdIV2BcZxCc84J3a+opFhf8nWLDzhArXBPXyPhrXwjYxKTnbd5tJSaqQB0tMI8DqRXvOxBJFGwbNsRBKekrUIUTthjUEIc+2w1ZajhNnCihAk9xo0GEXgUD4PJ0jtUGK9r68xURkNMmWoZGKW3sUKnpJZZ22Bx5vS7KSqeopy3GMFZjzlSikZEPOyz9Czj7mfbkDSaGTFaXjE6JLlQkmvLH7gi+8U84JZfUgizUMGKKQ0XqqGgmFIIIeo4rQxaFm7vBcv5XscZF4D2rwIr8T3JUjgZqQmx2pLX2SrQP0aMtDx1ZL26pyyPmPhsVOmdHmt5BBQjHh6/kh30rA5EmsyxtmSWAch68Pwp8U9qqGLsMPXiq8roCNUoRsv4ybM6RRWxpXcNZJqnHDxpjxoRXRCVj7CA0L4BhmHqBrNKsqWnhaSSt3NQrPZx+7O09kar4wXUprlOixmbQjDCn62nu707leLClZJpeBSEp7HLkQ8mcw55yLSgiZJtNByTIV4DIXntvWsERC2G6xkYoHOEWHW1LEiQxnnoJRKNc/Itvu+vhX98CuUIitBSawRnah79RATR5CLCsc2JIEdR6VNJIMzqc124Y4pUokph8woZes8Djs7QgV34dmT8L6e6aAhiu7dDAtI9Lqy5HiQsr8gPmtDXMn1iT1lwSMJ4FilBTKsRpI9MpkR4cnhXDPOw11W1QcYMRpZIE2Q0hdN9jTuJYv71zFh8Z6m0ywG0QlHXSFo6WhpiyIHQiI5OY7ZZzLKlzVTpYnZ7OabTS6aSDa52V3yK2IoxrkCFSwzHCQ7nVwM48R7dvcghdvY/Y/dsiKcokLsImbrhlgrvq1SrFWyAtCAuUE08mvelOPVPl+fc6ATvp0hGPchEBFyf6LxDqsZWSDFMZihZDFSNHmZ53x9F+Mff3NFfpO38+5kfPaI2ZEe8lKLxcKYAX4ilbdpED/eT2SS9wbeXPrtcbaYQTbg5ZwHNNfICdMsyALiWSC+FvC6lTTs9Kw576WfTZgvMmJJFCKurY50tK6fWvPfPONB8tiL4Wr46fOsj0FIY8uPCxLJVKNjJHUGH/yZf+3+b2lUuOO592UfypUaBsDKuLjRRQFDyCkshRvwt9rDgDT/kW2fXQmpQM5hJAmaQgRg+QCgaPNfBMVJwGj6Ei3+kGOUejSYlZNEJWkAMu/llr73fIIaiU8gyF2epGTMC4etYJ7qoLAAACAASURBVM9IXtYVnUKaMLnGiH6dYpAA1mz4NrrR0M3az6PMYGl2HoYjgkESkSRghUz/nPtZQ7zixRY9LgpiCSTGvQ9k4VCZRVvq4/C/MSUaoi0tjJQQ7YVBS3QV3jL2vHjQZs9wWTx/hXPhfHSXktBQE4lwihE+da9HIbJiGFjXYBnXVwSX68dOVerylBmmQJ1h/8Rfc/4o3mPIQYQ8C1GWAIVUdirT5kd5hsT1hD/nAJBGhgawl9dyPAtjCdZuSK4bSHR2HSHWsDc/oyEYyn6ZFPKaRZA0KtFPgpyFQ7FFI1zVPD+ivshMoUVthqcLqYXDCGw2iKIlegOPh8W9I+9DpZVSxLV4jACVY7I2glEIU0va4bGrhx1RjETPVGEjkZSXigfiAsA6CynXXYZZUq7JdffNr6dRueE0asxSUXnFU4TeaRueujT56XaCFCicAhl+lPHQSGP5eoXhNOJuQKLRjwyQxuIzuPFN7kFkiLDE6liaGXTKTnh5F/BSxSpuRERmwMOJqChsI+BVqLZ8XgEKIkNB9As1aGPXim5kJcthCxTz9ue2umpSAYtSabd5Iw1c7Me/z9D4+vGUZ63F0Gp4FwgPaI7S7LIMOyScEI+wI14xo8FTt8tajJb7zP2k4UKSmMmjJC/CvheGBVmy7LwCezJgzN6JFj8WTx2lz5IdnDYbX39Xup2duEYQkUyvzvSsDFNKqDNtwJLdqNashCk9Ixe27z6c5AulyPoCop94QlovNR9SUp6anwnlkEQigqy5EPEyajb68SGFggFJeM3g085Mcd3whSE2iBzP7qCxGfzQ1Fxy6/SqQqXj3FvwLPTMeXDLhWZhGN1g28R9jZIVt3vR46jVm2j35306N9BreIHgSGwriB7cCLC8umQVyNSr+pmioRYasVozFS+U3XkupQIxFAgZoAHh8fdESrF8bCizMBSE+hJGw1YjeY6cC/khhCOJLIfqQknDQBRjEuc3ymdpBAD1hxtTybnA7v0DNyx/Tw6luVEphXxRJNdiBHaNhjQSCGcf1ZuGLDCiNVv+lacbOwtFYB7dUYEMDbopqdSwTPRORfnoPWu4QaVYKG9RVAXiqWfc8CJUCwVnQ54gV/3zBT2Io5JAKIo0NiJgByjQA9GQwf/OxXe2nA1gTL/88/Q0PA7fWYlXPIQ4Iy00xGVBqoHkvcB0X8m6iMAITl416zYkEJcLM42eZ6REkp2X6D5GZXbSluGapPipoqSeWXBEBRMwmxGGIWC+5NpxH+P3JP9CuCkjvSpTQWPqa1eKwaI5zwIZ0MA6d+ZGUEt2hkpgRorooXjs+GpAFKANMW4fqP/u4WjUPbz5K410eBFT2LIW/IneuxqbvKeUEZa0K7ctWkLyXJeXwSv3KxFxi0cZ5trVmctiLPyLzWMk2SUQxHNPXRGUpzXbUAbi9/FCKj5LJLptI8eRDLtPbPbXeWR9s07v1VoYhCjFVkc7XYHZ2sarP7qAXIN93Et/SXICEBrwelTZBcbsjyQvMZUHFkuDTv7oPfENInoq5cjZFJfKmlac1hnqKdPerfXcuCprRENYUIHS4LbypHRPb7qBXZz/4ELzyD3rHyJs8PifoUMgGhfwhkQindwCy72XsbsVUvWYV6KQgjzCw7unZBgI+FGB0YhO9dhb8mnvRG9Acj6q7BmyKZ6RhGIp9nOZiydtRWhS+o9SJjvLsp37cqTSdTLUIigHsVzRFLmOrkAAvLkPf/N1IB8GO4TZFr0qyK9UI5AcBfm8RC1mjOoZkrxUeb06aP/ZDHlFaY4TioGks0vXVs0G32HkadfZ8Egw8ez7MLT05sMQkF+GlidOawhCspP5ZU+HisPwOL06kuUW73iF9Kz8LFELX+PrfozaWGQ3PoO1fQMZeo41yNpMxUkssMeh5DLghgka33nkW4Yh0I+qFarFeZTBMxmxd3M+loBjBzJjsdoyBWHYFVkjTx233OjwoITNw8qdI5XJswheLi7DWEAcERvnm8IlxXNHJ3BCVJa/02hT8HjGpZdrRbaiZFh6HtfO8KPHU+cE9PJcGxodenZ+SbwubbXrb3AOJB+KVQu47A1t156nVw8iMpAGsDBQgnydhq/PqVwLngIers957/i77XGLkK6QrrEvhf8SBFrIhjjMjqVBYa8O/hwfjveVdahzD8Iz0SONrzhyaJGFsTVksVbcQZqMaCwnblg0lo0wAKFEOtvrIVhTOTegai34SMSsvIkJ3KtEalMy28IJu+LH/caWk/TGv5EhEEMCtoa0rhwvcVlLYZ7mkJ84LSvIYjBKKZvuBsSbgV5jPkdPRCdx/qJnKABx4+oICX5CNtJ8RBHw8ypzIX17lshDDIX5/KK6j8gmtlVjPPFVm7sEmSyIMmoR5LmJJL3iNOwC8WggvUhf8wAclWzwPW9Aa6uAuFKQXpx/AZBt8YggSFgmYrJxwknUDD1QZ6+mYJGhCEJU0VnXACRycTkNHsHnWCsa1deN4Y3C1z2UMOVNFsizoQX5Ts/OMzeSdsznm5WaXA9yFj19feV56p4rYjxpGigNffEXKfOLfp7FuGRjXqJU6h3rdhyhYYYAOtK666T5flZWFmEFrZKqwXYqH5DpUMb9JAPJ3M89FjG81q4nZuUDa1rcJypBWworunurMBJ+fwowPTArE1db9p11INFZW0MZIs2n8Ka7ZdHduLGwCSjl7bHItsAKeI9GX7d5k0LLTZGWXqP5fbz2Ioh6Ny7BkXhBUyDAepq1eHwpZz3M67qw9FRIm6vtXxCOPv5FKjEuKqHAcV0wrqVxSdY9Qqfq0XnUWmqWx8uVw4gyXGA5u2RShmiLl/MfFEuimwa8secFDQzDEldCRXbOtk+Sz4hJw5SxRewfhqF8xdkJRfTpqP0lFnvO5Kcb00yd0jl59iVIbBo2FgNynYrMAemoiT7i7EeeJI2j/HF/XqJes86OxqfUhziesxdr5yg+GCi8v/8ML/sdBsTzIchzCApJZUpoXbV6nlyN4icUok2W8T+Vp3vtA+E5UQDDDhqwWhMiJJ12QVKe54hWc5qfgXMX4oaBf2XJu+YCy8Cna7nX7z1CkQrHMwzz8yT8XgQ9vhb9QKalgBPVRfq3LbY0vCOwCLm4rnmQzcqps+M5Xy/1CyQ7g4PhGiFrPSL0SGMVncJiTeaI23mvRSaAXEo9f6OspehZABhOCqaotTOUhhr4vud7Sc6zahJEvkg0ABS4H54216XukZV7J2dQMyepuO5wS6gndfyL96Jcw8+2hOHgXpRwsyYJ4hpEKzmOpD8ZatPI8D1+v4I+UIxanTPir1wPy8yMKWCCZQ9MV5yhMLrclMVZDApJ2UgaDyolO4dzLPPsIUtyH+Hta9GWNwGOdCvHWpnz2tzG0UH19kHuOQRflJH75kc6URWAC/uwCo9CRGJpwSHi2zz12XOtIyZkNsLmFkSnvxwVr7GGZaNCeWDd1rnhcwpWHm7S+Md0MRiiqRmIqImoxVqBFmncJ/ApE1Fsxffw2hRwfl5RroXs40kPG0rVA60uKkdD+Itn67NvZwmT1NOIEXH6mvoeL9VJc89r1zf3/uGFI71pM4rTzj426x3ip1epOFLWOgcAOp0IU0LBNdeJHBRyTZdfJDATJdgtkt8IJKU2T1fjwLixISJOSBpBW4vWwkEGWqGDLKglQqk0Qk3IarRWumX5P4UVAHFBGWawXDnCkcIWc7MCMu5SgvpYvWqgKqEJ9axMQ8S3Aa9R3gcfw7qw9JoeYtFmX0LQ4299BoZ6zl99w8wARfms30v5CALYXOMZGgvvzPnbLyztjuxFgeCBdBbyQgX3eLh6ld1oiaFBbLrvUWuhCJFdIrIIgfU1qWjEBX93Lwlo9rBQuBHj+xd77rkQ3dVNmwacvI/Pa5k6JVpJVLO7SClrBdSJ0iRHOfdsxss/tlx/rm8QmKlgCySEDEeCkC3vg88xJ1nLw6kH/749dyO8q7dH8gXidkZ2vQZEqKCVUFWuTPyPf4EqWoQjtYq4hillmYq58UkgHzCksIZ8GudSTRgGCeWnMNETBOlJ5RYjzVhVyKrJ8Gw0LtyVOCLuizFNptveNSuIp9YKymMM7IU9Y0vD4P0k6rMzIC2e4cmH8UKaHZRzLkK8uYfBXwSHIr5IwiyIOuyMMKtFTYcoD+lwk1vaP28iJFTOyRVac06GUOhJXRnbmGiN6WPOVQwhgE8/B0lGyc8CHk75ISYe4KPHcuO82B8AwBAeM2s2CgIJQ0tj5MViTaC9svIuqLEuyHHG1L1ZTBvAxjH2KT8l6qigNnyBvxeAV6+6Ae4dzTMhWVvB0Mf+Vvtw0BOnQRRLuYv78VJ/EGEBjasI8uFJtYzat2FxmAxYcEG2yei9Gwka++GnhYunz9CFqU8L4VhRwjWu7f2WhoAzpcNX6C7jBIHVZXijmzQ0ungPNA16HFG3OL/FYwihKKx/lj3btSTZfW9xj8G3gJ21IrZFFlK58kUXaRoYevrWYvKhwAH/R8v/13Cpe/MWZ5ZlcKXxcy7ic6Iy875S2qqZYo3FoBUEQy/G8xluCCOF2PLgl3bnbcYtJ0NnxNPT3KCaMZOsW6m4WQAZhxKiDFBsDBI3FxNvDGTj3mD5ACMPM9jz1NNrjNLC408boI1OxNnfEyX6XCNLkAbEvD15iMHnRImiEkvuJXtutGZQ3o/927NcxCswNQysBEynIqEgnjTI6qESjYL4IynIQdj/XQkAd8YBoiFiqKiJVzyGLRyAcj7KSqW7yVJUcNIQkaR0AppPStOsMbH1ttRjNp6p5GmDSEc+DLxmi/y4PFGbPwqgx/2S/LQwY8hr+hpohB9Ax7wwNHYt3383cjQU+eR0uk6WuwvgqdVR1zsqO2urgegJoYReqU+ZleAXu1aJCzLhEze4+XtYXRlQ1BbCzpJkaXm0w3Ory/4CYRhQrDlb1ukM9WPxjqARB5QACOacTzF2Ug7U6HoHkQYGkmzsHlqtt9NodY8Vd3sNej96zRIiQbsVPmk3mavt++KsAcIYMJWV9RDAojWckPD1j7rCq3bv/9Fd33VhBLXyA8pTqHw+bUf24vTPsH9HFbSAwBKGi8RtKIL2kIc89cql4DkOfr75nO1zgez4el3jNnipOQ15ObDmzXttSZacTAYbNHyK3o13CvTj4Q/5hN7XadBCBzRkN77E+YAwFGUN6OGVXdQdPShyRX2/wxFL2XPUsIjkLo2xhAyqMD1r60EUxaZ4OWCNJjgVRdSfmer1pfOvzJaodh1l5VWF3eM5gVdG+s16gXeE9vFMA2S2omkiCW7qyIcUDfn0MoghF2+4E4e+aIFJsnI8cE/Ti4BNs3ssLrhkZ+6I70pzFRoem7bB9rlbCbvuep0KXe4XIYKHJTyGLVwTD9GkFmQ5cjJ5cOM3rtzziBsm1noogAEsFgtPFugmJLHspESWRzCU9RLkg5IDXsT4DbEgH2sQh87KnnP/UHiAqCIFkuhkfU4Sd0zXsq6D3skKxxjeUWjdHPHUcSgNFujMFGsOtMK1MLlAymJA8iQC8/d6TkbzM5AwZBkmZ2GcQfldHcN31UbEfvhrtAEmu2MxJvbIwEXx2mLceY3wgGG0EGux5FdcbsNIAcFhBWnZAjcEWhAkylhYQSSCWYQmghHTJKiwvSMWifDO0pFJYNlJy9GUNgg8RGWneC+GNBw+D25u3MtDFN7TZm2CPXis6ogA4yoMjqURBehSai5gMJsNbJmJ6F5yLB4iAHEqMk6k1hiZm7ZIJfqS1jRhtyPh2KxDEUO5WwPWO1CfJ9Ot0S8ylJGe0jeGn2cam/ceZFHxyoYqYCs5aAIVAaRtJbEYSMmQgQBu8MhPFMLT19p01sfFdXFeyCoaUTxzD8MaHBcJMofkYWCInoK8FCzCnbZUHCsemxYGylCnIxTUg2JGiNtWlkcuOHqF8ydu0vhxX2fecbchAbIoyhTXwPQmjYcbYOvp6aE8jU0uk38lWqiOv9ZKgMhSUt4gfOoYwwVbt5qatad6MORZ9tkE3DBUYrmGTlzLipBcXhusRydU0TAMinGo182NhGbKknGVW3Y2sIkCLWfhWX6t0yavRy/HbEt9bXYORJDviadwFf5js/ZeFhLoBwURoEI+FocFkeTv8xJt9TEZqnLv4f+i6a34JolxDqF85C1Y3l1INYwWwyoNCAg/GSppNurhF+NuEsk0CiCBPAHTGvFYO9/I6EytXkpPi6yI8xc0OFEbQ+/ZBuS5Du43r4xEE9WISl7XsgSJOK30nJ2wuBxSrqjI06lalLnIm86JXvyFzgcbxft2pSaVZGSLa2T1I5WKGS9XRMlnmygNeK2sBYnN3dkPM7Zx3oQGxis8zVAUtFIAftZSIPaFvABf516wgKoex4/X3JAvn4TGdyyvwT4ZzgnAyNQWV9P4ydFMHHDzdXUd4JPJFN3KvcP7s1+FH3iKqkUpCgTJ8yJ8qFAQhmnxAXg6tsSfvEcIiGYYM03LYjDOY7aDL2FZo5GOxuMRjdAcCmTu+d1fy4c8uyCxeGvBV/h1KEws5iL5KzAik2iKhiJCFoRH5UlJSPMsBgu0kAYtMiIcG4fo6c7N2taWaA1wo9hzTxRG4NIA+TxlGBYhE/eYmZPYExpJVotCjEisKVQRAN63gsQwJA1dEVlLsdYKzpxYVWQFCo9RnJOIh8Ganh+Mx1OBhQ/pcYTGZ75yT5dt7AyN2K3KnGIPGDIqjOxsgLemI8IhdEvPXLgJH7eU9yyfZE5o3eOBXYsKV4U/U8YzO6iko69cdeAoSEJcJhR+onSOewV6KI15cj/y+knI5vVJbOZcmo4ULED8ORGahVgkImu8PpTj3Hxtsy4xnm1IZD6ANDLFIttYyO56+rNuYgkP4vF35Af8uxHZbhSaJNdQznAsnqVauQggP6eAjP6e8FLeOIaNZVxhlSddV9YI18ZRnw/CDe7pBFlCTk9NpBNCR3k2ZBVt//199TGQi5ZzqvZAYvegACyz4q9ROaL3pwsBvbVA/EE7jNEBPtkMVB7137ufTm6OntjLNNC43wdAphllIaQCeLdz9W0mkZ5nU6h+EF7DEBAdgdkGLSijxVytQ7V6ihZFJrnnNCaeI2hUCkmP7+c2ggQtXcqkrSIjQw4kzQeRgg8ruAk3IJ5+ta1JQ2EPle7GKgSaK3LkjzWs6CoBewnxBIGSFGrGpGR9cmzcE0dagBsDViwrjQMQ51sMpYzoXbR23oZA1+uo5jRvuDv86KUrt5r3F4dvbB7jzVmjBoKl0fRytJTd+mDayUofQ0O8RpSTBJvGxi4fudidM/H7sKCGGw5YKMOj5hHHa4QaAliRlz9+gPUQ6mSkeXoTYJ02btQ9hu8zMPKRCrJo4xaHPnzscYBns2Pv5aMLADtER0RSD7u5wEdn7xi7lLnSOxfBk0y3CisoeTakqLHO64idI9Pgc+jTGgJLK9p5DgDkCWgo/HBaIA4/GJbeSn3LbV97ZHnce0fGoBSRFWWLPSc/FilQoqblobBEh0leQvl8FnPlLCDUmlHRyWkURwZ9Qj6Vb3J9YvhQy7qJmhBA3RcRRAZxPZgxSb9pit3coETNg+sI07AInMI6H8T7KhcmmulWa+POTIcW4yElteq6qDQcgg4LNZsfQFMoRlmN0JEQFKbsPP04ECnA/rbZZIaDYUifgdVoWQ1xdliahSDzbJkPcg1UXHrKyest2laSntOUz0kNohXpeQM+ugFYpHXTAMHJzXh/jX2BrJLkuGnRI+PjKKg5iiEnAXoHT9+Nq/hbtrnj/V155snWIdCNe+xxy+85OMejWVyWrsTnbqFUnFjkxlABg6NIg8rin7QKDRB/pEGtLyEqKClNu+cIdDvtG0LmioTm73fhFQ+92JJwQc6hxRPt49EDzWNq5d54h/Bg4uEIhL8n27/sDIWUrZgPjXQ1h7Au5EQmAtv7XV4cIGpwtYxaitwLnlMR7jkYNiANrM5oNIaRomYdhyMANqgRtvsT1BRtZmi8FiRkvH65QdE0SokcQjIR55TSwnidxjLN2jB4mtWzc7HmKk03G59dj/bl6r8DEoRfxMl9Tr6iwmmeJh1XqZhUfh7KYvhCAtNW2xSEh85qpsS/R1kzrweJzMiilVooDHIMnllQtTkECcd70LgslA6ZRfBFrIeuwhhQ4IGI+W3xnQQs1l67kVLaZ0MvrjBoEoaC7wshmAsZ6idR1Q9qVR4i3h/8hBNgJZVo8zXjlS35kzdZdPgKPoToofvb83xI7LlzQkngWZoTEcp4Z+k+F68qyK5WHIOGgisNiE08EEsQgapxnaoAeeSgx/uU4/E9j9h/t3GlwdMFNYn8Ioznk86BWq8RfIrPhWNTX8c4YxJ8CkniMm6OFzkP9XVh2nNpLIg83FDE6/k7TwfHGoQlQnlv/KEY4r7rdybZiRRCQdWF2W2Le1tpzTxkECv2PpAwZL/NNkDX3peSx9jHlf0ctRctBZUKLBaDKjt49x4WGWq/Rwt4v7+wt6cilYNt90hauscWaRlXhwdOIY+NH4wz4JFvGUaD8GWxs2FQqfHwas0kJDVOqsYaQiDjyobPw2T0Pl1LtqWDhseGN2MJd90T0dPDDU1NT0IcNTmiqWR2RWEBH6vxT6/Ixx7akiUSE2Qlq5Hhm5QH+LqReIZGxozziX2gAQskVFCT0mgVlBCl7Lkfy+a0jhKdrLaHGxEFKNJLw40DvbiCKXMb6xD3sPcU7qhkWxQsGPN5i312UVjFkvzFM1OYMuVhr2KwaXyKQge/AoTRy/Lwyp7YtVlOnkaPSIHoSxdXjZ8oM0uJxxgKTsISrsjQKE8OBhewpize7j+qH7VDpw7rwszFKSQi4HVcBTqy8Uvvqdwc6GqVgkJiinn2tpVzhvjTtkjO+O+DN5SpxT7al9kWoNQglMyEKxS9mfh9oLAiMLLubWUbMU+7xopiiBRJfI6OHCYnCX1jakjlRip7YvIBMy3n5KnPOMhGb8iaFDYqCkNYNj94jDH5HRKEREE1ewXKr+Y6+TkOqzVZZnGiBD1Iy2xsTKNmSjOXTISFe4uO5iQDw+isfNua7TF5CA6x2wOlskFvZk4iZHD5yFqKNDZ5ereHHIXiEsUh93eZZREsUKmmh89u3s7PBMlpxt70vZVrleuAewbACcfaXwKBGvh7qnY1AfFzELI91iB5kN1oBdhthBqAMb0YimDBDQWcZGy5ORHjJ9Ncy1bNOLdUBLVSZ2tym6gFgqzq5BkM8gVxeMs9m0oKF5vucoME/qQxC3dES/k2qkxouS7j4ALBaqrQU8jxBPeQtgHA5LB7TgMR0DaVLzycl5BbjQLCQJHxp8IsCogircvzMyWk6N0yIIEu6DGbbx+9Tc6bip18R5l7YekptFGLEV6IaGRXyELjQ0WiUQ7h97MRbowFrtiOvKIoDm5IRMI4KscjNWzKOVtI7EZDqBxlr32OtclM+smsYqQcFNyC5Y+WFbCScF/3/CDC+ZQwLubARz8uyFeJ71y6RAWpwLHuvjb5e+552P5CijregLrcxOnThbwvv/hJcbNQwx2u6+LUKUQ87CCjjyyHdsMgXIiR1ZkCPtVJ2L8zBB0+bEE8kIghBuEosyPzVCo+k8iK71QqchpMoapnXqYNwGwK+zY0J1Y5VoZbwYt4sQlThf5g5BAdIp3WzGPOUx6I43s41nhI765FpiF0vkC7QpAe0BTLPh/NhovgSRugmEJgLGNkZe72MOuNy3Nt0+Zq4XxCeuHkXKo3tFOq6Y0tJneHEN6pGJoOv5YEcVfb46FAWVsKHvIT58TIgdm6p5cuew2mGh1JMbSp69Kn6HEpXs8Tj0/YbRTNW8WeJ0KqdQlV7FxptJyA3aVaZshpOMu6EqnA10kViEY0ggVRy7C33qMgC6Y0W6RYaIBQjIovN51LeVRAYdzinmEQJB8JGuGLOw7KdzbQsTm22IBhiMGHRevdH+AzmZLPPR9956giblLkJOAlWJrdrNmNWHwfIUrdoeAnkFY6+ApXImZD+BqNUIWw5C+i74Lu+kwRJKZ5F2dPXEAdVehmjeiwzQY6LnAxD1VTBKIWGi0gsxvSrPZk8Tn/Ty8xuWqEGFGZSRI4zo1IUaIh54o63yx5juIyrjc9FfteFk+CSD3PzpPMqM8mzea1xaAv9hwg8oyGwsFjLL+WcF7jd4rA4ppcsKirSHKR+2kwuyAHyrbsfm9Lbx/u3f5ub7EzLcEvBPGvOY8wcJn2TaRnWTMjNDP7Ueexu/dnJTlzGQfeFaihQyCVikDE145H8nkk3vcIyc0U6xbjId9TH4VYe1qI8JG9UR0I88be5h/O4AdzLzByjl6jEpYUmNhpZH1DNMqV/Jt721Tcotx1M3r34qcev9978+2479qrsuAKSOje5yRPqzLXZjU8mh3K7X+fvLy49zCIPNchTJH652S1J4xQFFG54EcBUWnGmy3tpBzi8vESNQGIXhZQq4cIXkBz/L00mHEDuniuqlQBoCLo8nmjYbB1UXeSBpYKLkDLZ3xaSwAvXAJ1rRip+AwfEVjWuIzFbk14jVwP/7v2DYLEQxmX8woCxPrHaVQQDcGVvRiR8sDqavC1T2D5Ob0+jcuyjb84kknkU7MQbA5E42CGbYhPp3Eo44oYOY2WYndpuL9eORaXQ7v/0giR0Mz/pY7sXpulYVB/hyGmhiwPF//ZKjjHAXHUnI8C5AGtloVGlK3F6VISo6HoLhwszGpDHrZibwi+TuvvIYutiz/bdLcFLwr1zacex3/xkQ/i28+9iPNrHneX4omkeFsXoghHgOh5KY40GAbB0sKCEiIFKsHS+EwbsFGOMl9fTmCyQYmlUFHOkUg+nY1jqVmf+kWlJaKg8lDYnG9a1hyov5XxvWeqPLsjBJ5SKgzZOTwaAfk9lPuyRGdBVCqLjYC3Xncdfv4n7sU37v8a/vZbT7ph8hCE01rsae55lHCHjBVuIprKEH3QYJB3f9wZOwAAIABJREFUQl4rUqu8XT3N2hDP0RCGK+XUqgBJ/An2HdiLzfYONhPiqEGS3haej1tbuPGmE3j2sWewveZ9qpGasWfvXgyi2L6wQRqjFvudjy90BKGVtwCybJw6aOHDamsPrrr+alz51stx8PB+tCbY7Ozg3Kmz+OFzr+ClZ17GZsN6CUcHnn0R6qgG/knZAXUmDY+NQmW4+iMf/qfYu4cP5XDBAJLA1HxeJ4V1nq2ghV4x7pXv27+1BzdcdjmuOXIU+8YR59c7mFncJM0QyTTHwPJZngPedeKtOHXujHfDt5BAKHitYd7s4OCh4zgs23jh7EXEUW8gjRgNUMR7NYRBLkr1yIz7AERaixsrAnRHKFQsLjw9TU2/UvhdsPMAl28Nx0uWHAjFY0UptLD7HCPX3I2TFEgqbiSjDNgFIAzgbu4mvnzMNC4+j2EYcfjgPhzYuwcDFNNmk4irfG5Y7cWv/tyH8fSLJ3H+9dfwzCun3yR0xokN2Nrawj13vwM3XXcFXn7lJDYTz4ek0ds9X1uPuexlKejivsVe0Gmko1giGSGsXsoBcr2uufkm/NKvfALvftd1+PbXHsbsBHOEGb5qP/MPfx7XXH0p3vmOE3jwgcfrpQAA+w4fwa/9k1/AvR++E49963u4uJ1H9kPdXBnrfDIFzO3JdPDWvgP40M99HJ/4uQ/i0KG9OP/GWZx8+TWcOXkG09Rx5PgleMd978GHfvoDuOyyQ3j56Rexs8MDfhrX52CzBfTSUREz8acu0zTGAFvLsx+byc4MDCU/7cqCoT4DxGFWeRL5ntVe/OTtd+HaQ/vwxGuv4uLccesV1+AXL70Ef/39b+Erz71kA+DBMTaccW9+eN9h/NJdd+Gfvfyie0M/0bjJp4QBwJMnT+LO42/BV188addjyhNwQhVpIMJJEQIXAxI5+6KMrCAti2rzJanl203iV3luwSsXaSD8tmnJy338HEjG/s6f0BCIGGkbCIn3y59Xe/bgVz/9IbTts/itP/miNT1ppcIWMMLLBS8bC5WQoU9msPoGTIvu278fn3z/3bjuLYdx7sIOuiq2ViP2bo1Yrzc4eeoMXj11Fm+cPoepd1x14gSO7t+DJ8+8hi899GxdNQcntn7D1gq//iufwePffxivn9tgYC1DkJIaBtIO8K3ftIeV76lZhmzuy/X0QuYIdVKLyWdEhiRSrLbnH/nke/Gv/7ffxSd+6Wdw5fGDeP6HZ2PfeJWDx6/AVYc7fvN/+iP8xn/1D7B/q+HCTi9zF9zz8ftw/7/7PIYrbsTtd1yPL37xYXv+rvC+6eUFxnu10u+CaICsxdbBQ/iV//KX8cgXvoLf+r0/N0MLWVTX8mtr317c8cG78Wv/7D/GH/2L38XTT/zQ18kPJqJBYU2auQ5mQOshtrkEJ8ju3uopSd3e8QNigK537G9okNEhiZ8bkRBgsY5TIhhlC//o3g/jW09+F//vA88bgPTr79tzAL/6vvdjzzDgb555wWbGzIQvHFTx43fciZ3tc7g4zXFQTdmGjynU1nD6/FkcOnEiFFx90aTyI0QHxaPGw4a7Auhu5MY4Gi7iR6398Xa1fZ4tJuGjLLw8IF4ENICdwkQEypoI7YaAnLMQYFkkpYp33vw27NMdfP3xF8xQEKVUfgEpGXe/4zY8+8RjOHb1DThxdB+efWPbW+yZkakpVAsle64JEHOsPUGH1vDrP/NRfOnLX8Ufff5VzPOcPIoq9qxWOHbsCI4fPYijhw9iaIoTlx/Dn/353+KrD78AEnGGppCoTAQ/cu9d+MEDD+Avv/F4QGBblyIDJVzIsKUH9I/wimTmbqNRZIlAPuotfN5sgtOdwzFPbkZ577Hj2D+fw6mza7x+6hyOHN6H5185GyEbU+Inrr8azz72NFQVZy9scPjAXlzYuRDmRKG49dYr8X/+4Z/jytVxXHXVQd8JKivQg3y1sTc2zgmlxuLrx37643jkr/4GX/7CowUlAfCsSbb5F+xcuICv/+nf4snvPolf/iefxb/8r/93nDu/CZno3tvEPs2Mm0SbnI7JUUcQztqWfAPSkveeHpa8BZuyuCBa+XSy+x+5/W48/Mz38KUXX0T3wi2SkBe3z+O37/8C3v/2O3HJnjFJSPfYGBquuOwq3HrZUbxy7mxyGo52IixyvqH37pOhZQZqY1qTsSQytc/+vJPCF9Bj8UldwpDCiR2v2szsxLwkSjlGwB5mRDHpSazF80+YwahrDBKogssuvxofe/s1+LE7343DW0mMhSJVwhGmULdddwW+88TzOH3+Ig4d2GtbGGXUujxt2hoA543e1NXbhBiquPW2W/HcEz/AA0++4oaC5fJG+m5vb+Oll3+IBx95Cl/42oP46688hLPbipdePYUoV66lxa6k0gbc8bbL8XffeTIhfbQE4P42hEIStQVpmjF2hhoU5jSgquWskBuJ3Z3CY/8q2ene/sR1J/DiMy/4dczI5nyyS9Vllx/Fay+f9i0SzD3RANCxdfhSDNtnsM0GUT3vz4rSJmPOp8YvQk9f/95w481X4Nv3/wC7QwbwnAl4riXJ3JPPPof7v/wE7rrvNuhirbgWinyMoXEjNCg1GwIoRsz+tGIn52Q1pjd3WBJ0BQm8NmQNU/AUDXdecSn+57/+KnTjbdUmP0DlC7Vz8Ry+9NxLuPeaE/iTHzyJ6EbVrYbgM+94J776zFM40lzJefqSBqWrnatoA/Zu7cXOZu0nVj1VNUrhLCRQAYBMPYqEURGSrfRuhTSL9nDS7EQtEcIwhtVnJ2+oephEmdUIRUzGChPuHbo/dc+duP7YfnAhjx46hFEnbO3dh9/49IdwcU10ZNe7eOEM/tVffBU9kMyAY3sEr1+YMMqAXg+GCbuEeSbLY/7ohF5SsnYa1crP0TsOH9yL1994KYXJHUWTAWjFMyNrQ/buW+HiufMmBlFi74Sfr8OBI0exPvM6tic46mApu5OWZTyIzILVRqiTwyaHLi/l2aSZRqQR4SYmiRuNc4P0LiXxjOVFcPwtx/DqD58FRHDsyAE8fO5ihCisSFUoDh4+hOcfex2qigN7Vji/vXbUY+t27PglOH3yFADg6NGDOHvuNQTqIPkNHiQzBevavU9FfXhzFuwJ/Pkp3tAGMXLfc9fHVHx79elHnsRH77segu+E8osMHr5QNiW+0wRnNsRyKiPaIAvv5TDJHjQ8Zj/OIDMloT4JQABb+w9i3jmPHUghblx4m3uHseHbzz2Df/TuW/Anjz9l7/HY/bq3nMBq/QZeOb8B5Fx6viC6nPl3tHPZwYM4efZcGiMihnoQrXerh6ndoocVRB2OMd26u9aCuXxJZKObjaVLFSXdqWBTm+jzUbGjAHu29mJraDh7cTvkWaH4/77xAPhgQ51n/Eef+QQ+95d/hXvvuQff/+538PirZxMxzVbv0HluQQTD1h7ozkWsFTh0eB/OnNvJbEz3JitwdMSuYk2SrDbtcCOJWIcnnn0Ff/8Dt+Frj72EnQ2F1bNX7GkR62NKvW+rYT0pNOJdpMHy/qBXXHEcL7/8WohjGwccPrAHb7xxzuRAi8xQdCPzkqn9Gr6FEYRxOfHYCggamw0pjA+ZNwv+JIyokrC1NTly6WE8/8Q5tLbC8Uv24rXXt1FJZhbU7d2/B9vn1hj2HsAe2cbFnaXSHbnsMM6cPAOg4aprr8Bjf/W9xdzMEPi4lcVRCFSgHjJWFX76qddwx1034uv3P8WrhGoD2cQ4DSggaNizZy/W63zuTeIV1m14iM4wV2DNhbwCl6lhskBBttGbCgDdrE3QpinqLhhzhzJ3g6rz2ggrbJx5rYVFXsyFzRqnz7yGrf3HsKXd6ho2G4gCn3n7rfij7zyAQ3tWOL297bUe3U5ebtbI05h2zROXXoIXTr+R2Yy53JdszaI2wr0I01+sD+F7yayLnS/Rebbv3R8o1JK8jDCjT/lUMq8FEcDGDABd8YsfvAe//P67sEd8rdTmNO1sY72zg/V6jfV6jaNbipfPXMD+rT04ffYs1usNNus1di5ewHqzwTTX9CmwGkfsTDbXy/aNOHlhjUi/toZ4onyEPGkQKky3NWEqUvHK88/gyw+/jI/efRMWJ1fZVlA9HItwQ7F3FFycAPAsSJT5zxESHTt2CKdOnYHOG/Q+4ROf+DH81E98ANdcutc5oh7GAb2jz5sQeIZBDBszdew9RdW7hIsgH2TstJy4AorXTxSDlM8tQdRbHNi7B+cuXMCBSy/D9MZr2J5mRBs7Rcx7HAU76zXecs1VOPnci5jZatDHtn/vXpy/cBGA4Lq3HsUzz74GtuXj9VSnuF6cJIZmGBmjtf9+4ff/Au/6iU/gxz/7AVx7ywlcc/N1+NBnP4477rwerEiVYgr4decH3o1Hv/VorGUAAkcfNiYfVznaXx912NFlzHy/hAGww1msgyCDT7eoCTGbZU5kGDDrGmdlH04cPoDnz11EtKdDjtE83IRTa8Ule0a8vG2p0NuvuQWnX38BL5zfxh179uHlufTN6Oodqyz8MU8/4m2XHcMXHzpr75uLt+ShMp7VH1Z+itWVpnnZL6F4mTf/ZX9LJDfhsD5QxGRGQlaGbLISUjxUMYV88dRZXDJO2LDvBoU+6jhskwcIZjRcdnCF1y5qPCpBVlsp3wo/Y9PRBntq2ta+g5D1eWzPPvcKtYXl3iXOr48jiJBG4yHOgOAb33oAGWIyy0Qv3aDzGoePHMPRQ/uhXXFw7xbuuvM2lursUkbzfjdffyUOtMtw5fU3AKrYbCb0aY3TFzaZDWMpuypas0OG8dyVIkskmsXvUU93AkDzRr9UnDinoaxzQMoxsZCvxTiOmNY7uO09d+KRBx/LOUjlBUZ/IkPDLXfchMe++2BRVPPK42oLm+0dHL/hepx74VnszKXC0+WudldLhOBIiJFUhCkd67Pn8C//29/G7T/yDtxx33sgOuPFJ57Ho999PhGIj1N8Pe/77Cexd/sVfP+7LyzWCM5fLJPgucBvOroAxRhHyHtH7ewdiMChuCkB2XvGq8jj2ar44+89iF+++/34rfv/Fq9f3AakYVjtwUduuAX3/+BBnIVZ/bMXt3Fw717g4jkMGPDjN9+I3/7CnwMKDNLQ+YDgNgLSjfsQiXTrwX2HMeycxhsXPbUGSY85Z/HKnTfeivnCKXzn+ZcRZdhOOqpXpVpxVYt1yv4Rmu+fGbJ4SnSztrGx0zJ6FAApC9EcnX3+Gw+4R+fZF+Daq67AfPEsXjh1zjmMFYCOPfsPQi+cxjr3qXAwNkadrTvUNE0Y24Brr74Cz730SuyBLUdbGPXbbr0Zezdn8K0nXkKexNQFv+NQqMy/ILmagVAFZMCN178Vt7z1OGRYYZy2Ia2hUXEJ9UMhga3VCo99/3v4wfNGCr76yqu4uO75PkEhX3soUnAYPF/iHpeIkB3ci6Qnh6GuHJXAh8C6YbmB6FnWjJ7nft7z7uvxu7/5Jd4I3c/Y0AAZ/7+FW952Gf7VH78QyNV61+Ta3Xnfu/DAV+7PdQQzEQuzimpmk88xPqsirGm9gwe/8C08+IVvxZyMe+B7LZi44d2348c+8z48962H8Hu/dz+go+0vaMDhM7V9t9/Ie9WiMApj89QpgOh3QFgfcFUAmXMxxDegMXTxmLcNePaNl/D7Dwv+4Y99AmfOn8H2DFx95Ai+/vSjOMfjD9pxflpj/7gCmuB9N70DT770BE6uLR6e1WvaFVH1KAtPqLjz2uvwwNNP5/ry4NvocWqfsXfvQXzkhrdisz6GB59/BbXfAIYx4vuIx90bS3OBGIC3HNiLV86eN6M4rtxoNrPH1VuXVKWUlCcAXHrJJdicP4MzO97gpg2465abcfHk83jh1DlHTRYJ3nzN1Xjs2RdKPUjWXRDZsHHKNM3Y2lrhXTdeje98+5uxDqpq3tkzCOOe/fjYe27G2C/g20+8BBn3pFC04ii8bDw7U80xv/BuYK8M4IEHH8YD330Ul11xFfbNV+PL3/i+b1GuJcM2UcWBY1fg5MlTePaFk4B27N1/EFceGfDSK69nWATg8KEDWF+8gO01iiHLqsaMursjDkNYxy45gnOn3sBm9s5Sioi14QbO7F1ZV6jvtw+5KTbThOveeQfOv/g0zlx0khUcYqr4ZlacuPkGnH7uGWxviFZ8ydAwTWvsO3oZbrnuEP7y/3oxRm2qVrqdKdPEbiBIVJavPJ5Og1AfOu05DlUM4xbe+f47cfcH34kXH34C//af/xucPXMe7E2aMxDUxxfWyEGKniVNatUYw9Uf/tA/lUMHV7YgA2Q0OCXDYI1cm9cPMO3YJNrKhwLbCgEKnLpwFl9++nE8+frreOrkK/j8Iw/h8ddOhhXHMOBtV7wV5869hpPTgF969zvxf3/z61hPJlhXXXYFhs0FPHfuYlRsJgIVNBnx83fegT944AHsTLZon3r33fjsXe/BB266EZuLZ/H8uW3s238A77v+Wpw4egzvu/EGHFkJHnv1ZKSEr33LlfjwDVfhkR+ewjuuux4HBsUb25vIdvzUPffg5993Bx5/8QWc3ijuuukm3HvdVXj81ZPoAO6+6W24720n8Oxrp2zsQei5l3Sj9bE734O2fRqvnNsJY3X7jdfj0i3gged+GPH9fbffhKNHDuGL334I59YTouN2gY0Qo7w+es9d+JkfeTv2HTiEI+OMP/naw27/Fddecy3+8U9/FD9y2/V46LEnIas9uOu2G3H18Utw5+034fJ9goef+WEYCuuVYSXBi54X3rRGpDzioQqyfQC333YTzp98Fc/88LS/xpCMtRmGuq699gT6xbN44dVzEGm45fbbcNs1B/HYU6+EQh8/8Vb841/7SVx1bA8eevR5XHL8OD718XuwfeYNvHHmIo695Tg+9fH3YZi28errZ0ORr7/1ZvzGr34a+9sGjz/9Q1zx1hP4+Mffi9Ovvo6z53dw5TVX4ROfvAfbp0/h9NltH7rgzvffg1/85U/g1hvfgge/8xQAwTU334D333c7/vD/+TzOnGd3KxpQ298mA667+Ubc9d4b8N3vPIOf/dXP4O57bsWjDzyC7bU9U+Tg8cvwqb/3AXz1T/8aTz3zKljFurX/IP7er/8H+MhnfhT3fOhOvPzE0zhz5iIAYN+Ro/iFX/s4vvuNH+DYiatw+9uvwEvPnwxFp7GsIZmZvoYTt9+KX/zPfhYXf/gyPvc7n8Oj33kK2zs7C4XffdZDwjyo/5V/5/+yWVGXzaYJj0fPdmBL1xt7tsXOjn33U6a6tjSlrtfQ9Y4/a1QRB5vWa/O80wRs1nj97Gm8fOYMZvWCL7Z3n2d0VTRVfOhtt+EbP/gezq392PpqCyfPncPxw4dB4xUoyAd994234PFnH8e5jWUp3n/bu3BYz+O/+5N/h//hL/4Kj586B7SGs2dO4Y8eehTfePxR/OaXv4mrDx+0zfYTqp+8/e146DmrEr3xLVfi4KiGZDZrHD98DG87qPjK0y9j/zjgnddeh/defhD7Dh3B2w7vwd0334L3Xn0UF7CFu686FiXgh/essBWsPIDesX/vFi5c3A5yc8+efbjp2B5ccvxKXH5gy1FZwxvziAPTObx0fgLPxhw/cgh7GrKeQ4EPve9OXDKu8c9/7/N4/o1tPPL4U5hYGj6s8FM/9m78zh98Do+8egHXX34MF8+fxR9++UF857sP43/9gy/j6uNHS5jQcf1Vl1qmYJ7Rp7WRayRy/XedN/batEYculKTl3fffAIPPfaMyU4w8Jqnkz0zdebCRRw5sA9srbf/4F5cPL+THcSGLfzkj9+Hz/3ZF7Fv/16s9u7Dr/z9j+L5l17Hx97/Luw9eAi//iufxOM/eB6f+NSPGtzWGW0Y8elPvhd/+mdfxYED+3Dg2KX4hZ/9AF5+/QLuu+dWXHLFlfjFX/gwHn/iZXzs4+8NXzzu3YcP/ejb8C/++9/G1luuwoHBTtlun9/G8488imdfOuWk54StvVs4fHALcMKv9w1Onz6N9Zk3gINH8cBffRF/83dP4N77botxXTx7EXrhDO7/u0cAVXSdIG3Az/wnP42nv/4N/OZ/83/gt/+X38frpy6EEr/7w/fg+UefhKri8muuwfHLD7tFUAzjHlx1zXFEiz1Hrw0Drn7HrfjMZ38E/+Z//B389R9/DRcvbqCBDLIBDmtAjMw0QrPrBD5zxJ6XPvn3GR0Turf/UyiaMnvA498i/jCetjwgRmsWjwksps1/VRZtRfqSJOAqiUT/OnDgCO6+4hj+9uln7O+ucM+9/hquveSyxclQhhZHDh3Fh2+4Gn/+xDOBaO697gT+8KGHoW3Ez7/vXmzJ5Nmbjvdddy2+//yLOH7oIE6eP29j6zOuvfwq3HhkhWdfPwO0hkMH9uHiehNz+8Dtb8eXvvcDrIYV2rjCp2+/Hv/6K9/GmZ0J+/cfwifffg1+50vfxBsXtjEHN6D4Bx97P47t9e5f/siCvauGCzve5Kc1fOA978Q3v/8wPvfgE/jgbddZVNQGXHFkH7731LNRBNVWW/gPP34f9rN2RARtax/uvPZS/Nv7v4uNCg7s3cKrp8+BJcPXXH01rjnQcHZquOXKo3j2tTOAKj5w59vxtYefwKWH9uHkmfPggavLrzqBT997OyL88ozBB3/0blxKQwYsyOrsvSC46e23Yn3yBfz/bL1ps23XdR025trn3PsaPDz0BEECjyTYgKQEiiZFihREmaQ7yYoUJ7GrEqdSqXxL5Sek/wv5A3biqCJXuY8ix5EtdzIlUSJlyaRsij3YgATRPeB1956z18yHOceYc1/wFsH77mn23mut2YzZv3ybTtOMgAAtZT7O/EcvvYZHHn0QDEOe7hfcvXcGeNjk73rm3bA3XsT3XznDejzi5z/zCfzhv/k9fOWb4W/687/w8/i9f/E5/MlXv4+ZqMVswQc+8pP40be+jtfvHHE8HvEXf/E5/Nb/81t4/vuvwsbAL/zyz+E3/+E/xbeefxFrltwbBn7m05/AvZdfxQNPPInT89dx6+AYJ5fw0Y8/g7t3722cpp/9T/4Cnn7Ho/obAF584WV8++vfxR//7r/FOL2CF7//Eh585Frko9iC5/78R3F+dobjLPPuvR//MN5y6Qxf+OI3gDHw1/+7X8Gd2/cwMbHsT/Gx5z6Ir//JtwA4rj54Bfdu3ZMP6P3P/TQ++jPvbZqfYnnFjfe+DX/nf/vbeO3VOyjtWiVg0F98fpMJwvaIhV7i0xyu3JHtwBgesyYyf4IEwc8tA7bfqw+FytOzloQhJdufBFRlr03+p16bJt+DGfCZ9z2Lf/GVf4dzhOPUTk+BZYfX79zE8dKDeOr6tbKdlgXXrl7Hf/Pxj+HvfuHzuH2eJeu24ARHnLnh8pX78aG3PY4n7r8GGPDMO96D+/wN/NFLN7GzgTVDvJcvXcFf/cizODucY93tcXp6Be979EE8cPUKYIanHn8bnrx0xB+88DJO9if45Pvfj9/59/8etw4Tl3Y7PPfsB/Fv/vjf4da9A07HgoNHKfrPfehZvPjCd/DDe2v4N3Kthwmc7MLh+fgjj+IjT9yPz33t+/jha6/j0esPwHZ7/NJzP4M/+NJX8NMffB92afZ9+qMfxre/+XW8eu4Smvv9CdbDOQ7HiXfduIHTeYZn33MDtizYn17Cr3zyJ/HGXPDf/pXP4jf/9e/h5t0D3vPu9+LyvZfxpy+8ht1uHynGY8Hplfvw1z77Ufyjf/EFWbM0J7/1wiv4r/+zv4B3vPURMY0DGZkITXPjHTfwK899EP/gn30RNvZQ38mMbGw6WsHxwxd+hMefeDz8UWY4Hh0nJ5dgtuDytev4y5/+EP7Bb3wOu5NTXLp6Pz7w9vvwuX/7bZzud7j80MN492MLPvfFr2MsJxHRsYFrDz2Cz/zMe/GP/78/wMnJCR58/K14aLmLL331RVw6WfDoO27gyvlr+NJXf4Dd7gTr8QAbOzz69rfjp555HNeffBJ/7T/9JH7tb/2/cDP83F/6FL70r38Xj7/n3Tjdh+J469Pvwo2HF/zRl78DFgqaDXz/m9/DE+96EndffQ2/9ZtfxI2n3453/eQH8KGPvA9/+b/8ZRxe+Aa+85rhybcGOji97378wl95Dq+/egtmC558//tx4+m34aH7L8Ng+Nlf+XN49PoJ7p1F0t4zz74b1x++DgC48sBD+NRnP4h/+Y//gNIbHJkIGD739/4pXnr1LrrvoRyTFCum/hZGt4H8Ffmqjez4Xd8xGCYmHLDlbZ/99H9vV67sNeIuD5i2aiAXJq4QZFDLsM9F3lwO0ZZeS093Chi445m3vQOP7Sd+7d99qRyPbNJrju+8ehP/1cc/gXk84MrpZXz4qXfiP/rAM/iHX/w8vvbSqxR0ACaeevwGPvDYg/j0+96H3/nTr+Dn3vtePHz9IXziycfwNz/3edxbJ26dn+OXfurDePDqVfzlD/0E/tkffgF++SH8xOMP4eefeQ/+6FvfxnPvey8evO8afv7dT+J//+3fx53Dig+/+2k8ednxq7//Zczp+PC7nsbbLgO/+ntfwuqO/eUr+Mwz78RTb3kcb79q+LXf//c5oXHKQTR2p/jUMzeA3Sn+yk9/AP/yPzyPv/5nfxp/5ukn8e0f/ggfft97cP7ai/j1L/wJTu5/BL/4oXfjnW9/G27cZ/i13/4jrJrgNrEej/jIB5/BEw/eh5/9wDvwN/7v38KNp9+L97/1AXzqIz+BP/7jP8bvfeMlPP3YNXzjh6/hfU+/E5999gb+1m/8G5wdJ27fPcOf/+RH8NC1q/iLn/wQPv/7f4g/+d5roOfdcjrczVdfxddfeBW/8OmP42MfuIFrV05x35UrePiB+/Gedz2Fzz730/jAkw/gV//BP8drdw6iGUUqRGiMojjm8Yhnnv0JvPK97+DmnXPcO3f8hU//FG7fPeCXf/E5/PZv/St884ViGzQoAAAgAElEQVSbeOCxR/CLn/kI/v7f/Sf44Su3cP3hR/ELn/0z+Pt/+zfww1duw+cRH/nkR/HQ/ffhs5/+MH797/0T/ODlW3j8HU/iM5/8AP6vX/0N3Lx9hsefeDs+/dz78Wv/x6/j5q1zHNeJT33247h+/Tp+/lMfxN/5W/8P7toVnKy38errB/z0pz6OGw8t+Pt/719inl7Hcx9/GuPSVfziL/0M/s7f/HXcunMI7ZoMd7x3B4+9+xm858aDuPbYW/CJn3kaf/tv/GM89d4beOX55/HPf/MP8dJLt/Af/+efwZ07R/zSf/GX8Ll/+Jt410c/jIceuopP/PxP4nf/1ZfxiU9/CDd+4v145NIBv/O738TPfuZDeM9Hn8WdF76LJz/0QTzwwH34s7/8s/in/+c/wgsvvAGk03ayHH85wZ/7q38W3/sP30LmYitqUz4JJtKFwKgGOOWdCGdrnZ+ESv52Ox7tY//z/3AbjzxyReP1UhhUEhRhMBFCXoRhVTI7BYuyO1HhNyZFWUQgPvWBD+PlF7+FL//o1RAgrCNptRbXL1/DR27cwLXdDj945Uf4o+99D2cttMv7L8sO73/L43jp9uv4wc1beOyBh/GWKyf4yg9+iHOGUd1x36UrePqxR/Ddl36El++cYRkLnnnr43jljdfxwms38ZYHH8Zb7ruMP33hxXBSjYG3XL+O4/k9vHzrLrDs8b63PYHz26/jGy+9qq185xNvxck84qsv3Yx6GM+mvpONdnf4qaffgcfvO8Hnv/ptvHLrLt7+6CP4ySffAvOJL33tG3j+1TvgEKC3PfIwrp8u+Mp3f4j1SNtzSBNcPjnBu9/6MJ7/wUu4efsOdvtLeO+Tj+Pma6/i+y+/DgB46om34ife+VbcuXULn//y13DnPPMDYLhy5Qre/cQj+P4PXsTLr98LDcQQnPqWuM784YcfwtNPvgWP3H8Vw4DX37iFb377+/jeizcL2NqABhcxB6dlRVqimafe+Q7cuB/4V1/8OnyuuPHOp/CBdz2OP/ny1/D8C68CPrE/vYQbb30AX/vG9wAHTq9ew8efvYF//Ttfzmsb7rv/Przrqcfw7W+9gNffuAOD4fTKZbz14av41vMvwh24/6GH8MyNB/EHX/ya2OKBhx/E2x5/AN/46ndwN0P773/2GbzjqUfx4ndfwL/9w69iXaO57k99/Fk8fP0Svvg7f4xXb94pf4xnhGRO7E4u46PPPYtLu4kv/PYfxbNYNo3JPIUbz7wH73vmCfyHL3wZ33n+R7h83zW8491vwXe+8jzeuHUPT733ndjjgG/96ffgDjz5vqcwDvfwra+9gKsPPIAbTz+O7331m7j56h2ZcJoj4gDGgp/9hY/h87/xOUSOHs8zoz1qPpw5Jk6Dg+9NWSAl7CsawnUf7M5d+9j/+j/dxoMPXLHdLok8YW/L6ovvx6zLuC8zFdMeckRGJAVL9uPsse1tCDAh0jqzEQyflv/XIi2ztBM4X4QRmNn+TZnI5KesJZEwov+F1azMiOS9vDYNzoKcfu9I7iJ6c3YTy3b3haRQPwp15nWU+dl6O7q3decBs6dEv55ZCqDsB2oLaiZpPf82dJmdxAFlrm58SaOnqBuMtTgiuBwHoTGD9EvFR9R0yNmLwtMHwX3jeuIz4XtyJVoF8zWl1PYfZrDZBxY1IdY0HtKhqOniDdFqwhp7YnCojz7n+u18vTFYtBw4NmZaRRt28Xkb/ZLJrD3Pxb83vMF6j54Amc/z5hEHs3hpk2cR13Jfw5TwcFhSIFSCHEFBNdWxTcPmxITM9XDAseJg9+4OOSPlyEwzg45Ms5z/MBJqMpvOIntyjJxG7uHE5ODibrMyT2JSGo4SEMrpsKrR4E8XOHzOZeQsU9v23iSM2qdjjsQwIwkLx1Xr20wn6/0vEwFF/Qn3gRPCkshzTbbsYLtdtc7TPtbaZaIB4CSuikTU+5ony329SFD09Yx97mdqFu2xoSO/eAaur7Xm6/NZnF2neObYOK9t7FoUhoLMav7Kbl8IwqiByjxV/g3zCbriyc9wilm1n9ueZdXotFRm220/h8z2bH/H97NvanAdKrEpmb6eBAChea4xR1y4d8U1YLbL/1qIGa0lHWlG92GKer3G++i3/p9rmu1zAEcIbFIVSK5UkobmwIykrz6oiJ+WToLrmaz7KDbp4u2ssCCyduYMZrdO2AlZWF/gUVUZPR9S6uzbvBHWccyZtSEuLcrakWjhj2ixR6IdbOeXxM5BM+rHGdd0oN5bZ/YJPWoxyjBNLVK+E9scaiWcEQlY1o/odOu5ktj9eJ6zQlMap9NW9THZBwMzsjfVQyLXUHUPkVIdGZtWzGzVFUtrN7R+ma5IkfvM14kc8hm6uZfHS4FUcicQn5DH0s7cIWbn4GVvodN4VleYk6X3CqHymYg+eG7slr4eK7V5dKFhqFZ4RFKzXSd7RHr1ytQS9XlHF1Q68/ybGrln6QpttR8JLyDuJSXCxK3seQGHO8dRVH2MBJKeh4gimx7rwIkYEtGgMkj1Oef3Zt5v1Z71bE5dks2YJCz5iRLyQI4rJDTW+yXA4J6h03rekYJ8wrGz3c5gFqXWNBFYHLWamsOE8zM1yPRokiMtmZ+hk1JwKQ9oZWahA7u9oK3Wd6zQYv0EZMWO/ScsPrdnJiVKELlVqDX9BlBCk1cnLzl2kALBampZIg+N1MvS80AqmTlHoUiNwnJ9IPJOsrmvxgSysCufx4iqsjlPQfrUopPFd+uGoH2uGLs9elUr/63xct4mkakqM4Vwh/qA8lek+SSkInWHZfQaIjWz8CkHOQv6b2owIPPDRPiex7ps1ifGcJoonvKPJgwLvkIgjjYygEzE4cW5GSAC6Wtkijh/qsKyyvXjGb2Y3GdEd7SmnMjOzt/MnvTMnWC7fAo4IRs23KHSmtj6AifQzE318JCQYbk6BU+V2dN0YO8JS3QEmo55vzrxFAhdljiakAIcYb7InEsxtvpBNBpDLNxT2y1Re7DbJ1qZOXej4HBETUz+CmlqOLA6NEUdVrUHu3214psrXBuIEhJ8X2nn1NDNdLkYDrZMOMlnLxRhxfD7k2JwA9A2o6AuwryZufFzwvYnWXXKKtUkIAmYFAzsdNTsVgfC/h9LtvjjWMOmX+RvQaVbU5CQKJlxR+czsM1XIUJqJpADKhZTw1pkNl7bV08oSrsVhPLuNR0sNjcF4tLOaClF4J3BIQbk7A7OeA3BAPTsThcuHqIBI/WimN9pU+tskc9O/0quRwKTIzapVUF+a2fuUgK8JwvQxGi2AJb9S9jbFKwPyb1ol4dn34+8r/wETkFzQWhbdKHTDBtUYRfL//OgG+HT9LAQRCC9RMl7z4MJEJECSeYHYD7gtmJ4mX81I4TfpHEU5zlswY4douMhalirATGScLfTBKzQOEsuqqAe3KW5pRRGLmyMbLFPX0cu3EYSPlpvjAajR95fYdl873goQcPkp4GwzVWE1HsgeJpAFS5iVGZDTDKH8n698Q5mmj2pdeW0HJWIxjGQoEZPW15Dj0OrqQVANjkpoUjH7ALLNoHaJ5R23xBACjyf1pisfjRQGpZafVdCqpsnSbhCid1hyx6d9AHV1WXymTXBi9DCHKlQxBDvh5OcFZde9J8CQI48vWENveih87Osl0jUUTaKirV6j04Jfm3VRGdEIi2nEqPmbQ5WzWEBYNZrLiR2MjGNjJ9ORKMp49v7ERW0Vv8SCIl2jKaDFBKfu74RQgDQGEvuE7jO/uELdIJ0fKKuXxmfvJT72Dhg8q7sdQhqtOao25R0U8jM5lAj02jDAXUQarUlmlVhqOuLiaHaBEUb+Jyskk2noO1yYHErgmODHEVlFjrrUEOGNPyHCKeYT8KADsgNlG8H0Q6+ck7K018IIJ19Vl2rBDv7/soUs5w+NuoZs8M5/+a9iGyiScyQGUIUxOHAQgJyltmF5ZBxm9alE4w+H8/PidtIE4VK6oIz5XI9bx8KXL02hlCAWT1/L6MPx7K3tWevSqNmNfkVaCJaf/40Y2ok4wYO6D6C8bx0dxTn+npfUw5QklDqIEYOxEBALtRzQQnws2ZgRy6djzG5bVx4vTelYYiawqOeqSvfMi+4li1WAZgeDtDXQWGR64l+FrKVUoKxVRz6DSk81jXgPftGUAjMmVA+IbWEiG3NhCxOcqyhrdchxhfzsTHCkqgkpSaIVPiTvSYkeYdtoymwejauh1qCs0IccfGlHLYdViNNDffZnKquZ9GhMBQISw1HZojDNQBYlpoQvx7hY9kIuUJoBjlFqVUbjcO9ESSZqJxU0TR4KdOPhCyn54o+AEfPf1FgpNDw9A31KeJhBsza31yjq4KVxFn9NIE1akaMGrVpSzqyx1JjJAU2CalRCNa4HSkwm4avtnNBR3TYu9aQnCJTaq19QGlaIB253HrjtfOPjQJpeKgJWQMTqHLfo3UbFCb11lci9+LNJezYrK/OiOwdodcQEjOXR1TnuSJvz85bd7OokFtFt0ohuLvvAFhvwuHCNHxGL423sf298hgIfWjSOLamQNPg0dMSW7uXuRBCAwnhAWCXWjQjMaCPhD6TkfkGFCJd49sS30tHZDR4aaYKUQURyAwmsiQwHWBlsiBgakpcTnDPqefOiA0ATvWmc9VT60fjHA+fBxmYFaAL7xdCzTRlPqaEE8159s2sxkX0+XShw4I2Ct+E+PpMIwZpSyII2uO0p7vS6NDd676eZgnnj4oRKTjiehWUMKGUnnQGdzgVytoc5jlSkQikGvN6e2aeT/gdTI1sh9AX1zhkbjRHfM9tsaZVUe0C3Y8bxq5uYqHd4xF609waSRChSR4xFcrAJudBCVcxIKiKvyKaUUJg6PUScVV+QYKlL0e+Ka2H5w1w5GHRw9R78TMTWQCS1m5k2FzIIQYLy2GZjCIG4efAZ0/CX9cSFBIoSehokY8Lv9kkVwLtuFZ4VWHWoVvassumwHuwkWtSaoY617o/EAymXIORWnbCZhNu1rpLjSrF1+zT2Xoxal+SpKxNyxbkzGObEz7P64hENeyz2BAcEYAQU5WTwxARIt73Qv4CL4HZmr1upsHTIUsEk8KJEZ+5ah+i5UEgQuM8C+uMHVpNQoVjE7wlRPkEyLzptFPyk0w8RzFfan9eQ1oXKXB3IfRZkbzJI4jeGRUhgCI22os0NV0blYqJ6QLdfLVkK++av2thu/BfY7G8h/vhAiOmoGhzTMD3U0ilOKsz3yDdMmsufn872a2hJJ4Fui+ijI66LhkrQEP5MQYA+A4G2MlJtInri7YB7KMbVEBwSvIkhtbVSH4E3lhMlJK/zzmlJp0p8ZUpml2a8jN+ziFE6Zzk5ziDQw1BqNGaQ1PamYjIAQnCtP84GmAmdG/mjWxbh5rdKtmGDNB8ABJMXXOOnUb4FVNCoEyCzVM70A6fazWvUYd1wugkBt/Cxv7bZ/pc6JFnGNZrbwFLJqrkNCNRyf8w5cAMOg5hHD4X7lcTUrYlboY3RezKxKTACDoS2oQD6wFg1mRGCeQUlPORkJ5drnkmHQHEd50Nb5tfIZhuFo2QUXRw+eyAGLqnUG+TlrrTHoVkeG0n47q+IyFFAZAKi0K0fCL8LMPrzQGqbQ9hXSZGExBqFlT3D2Ty5pwPfpc9OK1dh991n9hh2bma2XBNag6LDSF37zI4CxWJMHoLPmoa8+a85GdzwhiRAE0UMk+LjPjhUJoxCYbdpUO7DPlRbBQDs+19CJk1O1k1+8wGsMtp7kx5VjQAqaxS07Qs0UAfVUPTMHUqubVQR7ZhUzfsmICUwmENjUUmdjTIHYSP9VDduRR1QWhOoSDmRORhT6YGryIEcBYrKn+hOx3lH2K/EQJUGxEFS5PFEJpdZy5Thr+DoMuJB+1phCBzD8QMA8hW+MVgo/loijlkPswKD3JoUk33Sp9HCpRBYUjmNoMZw9/NpGauRWPCytBsqIL7QD4Bl9K0dYsilIOR+1MCgs7QTSZp7kMNHertARmeDrQ3L456xNbE4L6H6ZK+F2uzQZzoZRbtNgTCM6a5YrmvOzMEU5Jp1q6BgJ5x58ckYI7ec48MyO7UXPPf46SEC02UhHbSaFYLI9rwbMgb2q9B7ITt6tjEDWkNVnhN2fq0oeVrGbpOtLKbkKPv/CzWIgRlhUoopLJlnqAqKSbzIyh8DKbGs9VwNp1aSr5BCtRFr8scW1JDNdRV6b5IQnKw47ZmpC67ECZM+kpC2mZNJgMeV0UosDb/DQVFEk0I5RyFS4KnkON+ZvEVRjmJey1M7PnadBzNkEQAQj9vJtgyRwCw5kE+Ff6y9BGt+ry3PROaS4FCRDLX85b41BB1MummX6lDz5h/AIhcGDIhNOS4mDhvLB+FZtGksGOh4EWnYg+9giMnvYSacE7O/2DbPQcRV7lIecXZBEsPi4KfdtJWDVTmFQwDO19DQPhKR5BHXkIygC+ofIbUXji0pJ/jIW4yrHwMSchOry9zGLKYy5Yd/N5dlOPL5EvgrA7QkckcDTJ2Ov+YoWkURoT2DL0BcpwWGjkPQUIScgMOZ3X47O5EwYQd/CwqTgFkzkRK6Rw6ZEvXYIDSvEkqM2edSAtb2dyI+6izdjKYJ0N6wnJD7m/uCzt/q6APgM8j5qs3YZeuYpzuYWNgnp1nk+U1CbZpdV81sjK+n5B/zhLcDTlEqvqMnqF+LKackcXo6wHuA2MXuQfr2V0sJ5fE4DZ2WM9uw8Yeck76rDkmzO4kGuumggNzPWLs9oDXmdNxKOSQqCHoJegv/E8tB8YN0w9CDOz8xUIuhwedKMmMTutk3Jl9P/0Y9JOCgVxJ86rGJdIcPJbQc090WULGaY6lQ9aoWBPVldCaTWHkcxugoMDGrEHRZRDnVmckeg6EQROlBPXKIUcYmJg2zCz6buYhY4l/Wy8k2+2jfmQXlad2chIMoJyH0PYqROpwlZoXUAcrPx6qGKyvBaimOXxjyWfZn5RJk4leElQNVWCuZcoksVneq1K38+BHPjNTw0cUSFkznez0Sn4/cjqw7CuPgyGysWy+U176eI9zT5R/oRyCEaMTGbZlmDVNDFtyn6nR0pfi62Gj/eCO4wvfBy5dht++iXm+Yt69hfX2XRUB2rKt/4m+qhyiHIhIHbHMct9P2rPscXzjJuhQ1es5GWye3cFcXfu+3rmTlmPUdMz1iMOtNwADDrdvosb5JSOMOnM5WDkDxAbOb7+OmEPC9OPm2PQVisgJHcV3x9jLLKIwicYxjb4tZ9AifBdjOQWLqvjZPjg5rsVakv5fM+HmUYJIZ53vzab9aaqYfu/KbJPKSaElQ7HMuUqbLzTIMnkWiZHFGF7lX8Ywrta0YKBGKg7bZQp4vD82nnJIkIcW2adGJaF7ONBAP4LsviauFuY10AzIZCVP88SsGtGSAfib+Ra9dZ9ngdbZWRt43H/y3ukcdaC8/7yWPP5WwuaCXb1Jo/Yk2OxFSVOkNj43yRqREMLJAWvSnqrVYF4FiUuCNPZEQiOoINZ+OCtHKV8HtVdcY966CbtyHcvlS9g9/AjMJ/zePYwrV2uN+ZtMwhzceE7ec1Ylr3syYAldIMKABdUJ3RfM8wPGriZ8IR2gSjhq+S/hIDWA+SC2JWJGa+Z6nswWDu2LZ66xh7B6P9cYUQA0gdD9LbxGMTiAnGKWiIZ+DCo0cdxF+gP6QGJFp3I9QwI6EYaXecFqWq2bomAemj/D9KuHSfmznafSnPT6fUGgeX8/7jf0DI6qUm2oKO7rw4/T/HAIITBa9mHatcqd4M8yakoZswiBanhDaMuD9EQSTN5B5iNweA8de/Q9dFuXQoRMJkm2NWv0Wdm8qAM/z8bCayaBHQ+JcGINznWIQUJbR5Zlg5hKJV/FELSNlc/gFVYFkNBcJ5l7kRPLZZ/mXvP+84jDd7+bvGg1WkD+nUqOoqNzff0Wdg/cnwdrGJdPMc+P6T/NIdbrIX1CBxx+9GKik7iu37tTPigKSAk8ANKUVBR0qGbyVJqcku/roYQn7eT1DDIj+cNiM6CEjE8c7twC/VJmBj/cw9ifSNOX1y1FXjrPvTFb/K6paDX1K30kRH/0QTT/VzkLK7KzMSl0L0AOTgnxo56D7FeDntqZG+rMdT0KESaZWX6uIj89Ndv0POmoVPFemlNtypj7mhWlrjUU7c0m8PhjYGNfmku7mrJtIRxsbJGCiJTXdtnMOvjRNA33iXkYjmRqlHBocLg0bfobGHHABENXqg8JyoQGHPGl42Ez+FjOwhxOxPoX+Q6YM+HNEUdtQG2fTXeCBkpr2C4F6hL+FOtCsOflx6ZCNQkeRKO1U/iRSQH42T1gOcHu4fsxb93FODWsr9/C8vBDmAnhsTrG5Uuyb/14Dmc6s6JBsUfrGzdhJ5cxTvaYZ2eYt29h98BDGFeuAIczHO+cYblyCWc/eAHLfddx8uBDWG+/DseC3dUrWO/chp+dYbnvOsyPsN0JDjdfw/7+B2JtcNAHs965pUjGPJwBtsfh9VdhZhj7S7B5jnF6JcKjI3pirIczmM+syp9h9tjE7nJ0Yj/cuYXl9Arm2T3Y7hTnd29hf+m+YI/1GEigJEcydoVWAYZR82zNy/fWnIloAgew7dwOCzapSEirRwGPrqGsrGyt56iUA0VyqNh0ix02eS9JOxJkjVYn/RvS+MQIXUDRuWqFQNUng2tnEljerrhJ/M7isryWMd0OfihnFyTlG2bhvydiqjjDkiwPz0gAs+xicc2xtx6zWQ7DhQ7lWcCTYVeACVYURiwhZ7OVdQ3fQYva2Mlpfi6YbzNVTIRCpgVwOChyIPQnRGN6ZumGJDCM8mYjW95B0RvEXig5KR2ciUx6V6kSEj2SY/Dze5jrASNDiseXb2OcGLAa1ldehu1P4euK5b6rAeWXEALjyrU8tgw7ziPm7VuwS5cwb97EeOh+nD//PE6evAE/v415ZvCzWxj33Q/sTrBcvYb9gw9g3nkD8+jw8zeAy6c4e+F7OH38CRzfeB1jOOa9exi7gfVwxBhBVMfXXgZswbh8FSf33w8bexzfeAXjyoPws9cxV8N6dg+GFbtr1zDv3cI4uQz3Fec3X8I4uYL1zus4uf8hrGf3sCwOtxP4+S0sp9cAONb1GLQ+V9jlYNSxnKDnYQi2O/MkGCYkLRzKPClJEIcvhifblQA3r+iMeleoTL2+36NJvXiNz8R7VTLVhLdnrGgEABsYjizgRPog4skGdmAp/+Z6DSGJdrU/FbXZppIXyuhCx7zStuK1CSAKyTy6T4XPwOj0GyMcl4MdjS78N7aLu2j7RyelWUxIqH84L+RCZgWg9O80E/wQTrxonDLl0PSMzPhMb34ymwDAUjYwO1nZPv87uQQ7OQ1HJ00bmTmLnKt0WEbYMR15ac/2KAazPMvWAJRZaCnh00sf5e6tMVCH4yys2+/gd+9hff02/N4dLA8/BD+s8PUc884djAceCERxZLMZh5/d1QAozsj08zNgfwW7y6ewS1cDHTz0GJYrV+DnR4yrV0LgrBYO64xsrXfvYX/9ehDQ8RzL/Q9j7Aaw7LDevY3d9YcBGEY6tP14jnH1OnaX9oEaRoQh5+qw4Tjevo15fg/L5ctgMeF6OMdysgfmEethxf7SKZbL98e1djusxzWTgGOe61gG1rN7OL16PejB2WCIJkMypQ0A4RS1sdfvsZxgLPsI/5qJNoj6+t909lUXK0briAy61q+/I6kMIfBRxV1VOAcwB0MEnybslHnEUOraXmd0wjW/Q8IMDLmy8G1gYBdOSVv073DO1rDoIaenoYYNlR/NNr9Rgid31zRDgAzBjzESMRgtQUMfeQn2YZCmzE0UGmmQGwh0kQVi5TwkspgNAaTpIIZqLfzSScp/M4qhStL0dcjZyOjI4TyF1YwEHz6THKpWSCQrXnkvEoEkuKIBpUkkMICWcBahLTowPQUd/M3IwpY9cPYGmHthuwFfHYYD7NI1mE3Y6WXY7lQEPq5chZ9nB7P0s8zbd7F/7FHMO7cxLl3CevcMuweuwdcj5uGIsRsYV67B790C5gFYTuvBfYXtTjDvnWF//UGst29juXIFGHvsLp8GIS0UxidY9nsc751hd+lUeghwPd/pgw9jd3IpLj6PgYjgWM/uYHf1Oo53bmF35T6shwPGLpCXzQPG7lIKbMdy6Vo4RMcuhACdrcse1hSVEf6nz8Uxw1nI6NHFfAoxQ+p4OoAVNWhmStjRYiNvpodY6oJAoANTfgOkkONnZfpw8E/q8y7EkpGH7VH5EwNDAkAHB/koMjTLie2Fmiz/V+abpwipfJHuSG70DCAzYYLpKwMwAfjhoI8rsYf+iXUmIov6i5g9wo8Pvad0WDnwPJhzv29Ncy39Ghl7twEshPwJ3RmWY9etZb/tg6Fu40jGT83jDtudqA9FrLyFLmFbJ671AqYOJXOP1sxmnOcSSrweoaiKjVB2o+plDGB3aJo2gMX6xgK/d479O9+G+eqPcHzhBSwPPoJ55zaWRx6C370Lu3KfzA33Cewvwc9fwOGFW8BYsH/kEficGDvDelixXFtSmGbC1jHyJQ4vvgA7vQpMx3rrNYxLJ4BPnP/oR9g//CiOL/8Q894ZxskpxjKy/mYNwmabQTY9YoQMBjTnoQ3D2asvY3/tOvx4wHoI5+Lh9i1gPeLk2sM43HwJy27BMQXBejjH/tIVrPdewb31gP3JDsvJKfx4Dxo+7SFwNt3WjFmU1P5lEvMcpLxSkVXRFZoTk/C7OS68HIjqtn7hM5vSdfSMTrJb+URCIACcdq7i8B4UaKHhEk5cLPQc8l+kMCznaCi97n/hs9BXobT7Fs2p10d7PRCPfex/+R9v45GHr0Q15IWIRHbBtmWnGglBaNVM0IFUm6KKTUBl2epT0Os12FaOB0pNz4Kx5nSMRjLRaTk+/uaiJd4bnpmejoKQ3YHZNhB0jBIJcI1AmhzOxHaD2X8AACAASURBVDxsOmQDQCs1jiStigRZJ9ZurhEx9V6hfLZW/bsxVfowp5a8tfEr0WnW1ylKbsRCoX3B+SpGT4Y8vPIK9g8+WOcBbKNiG6XrF/w/Q3tFNCYl1FrroTHJpr8HGlJQZAUifmUpdjtdfoELa+X+EvE6Wljcaw/zfZOD3/PS2zOv66aGptOaQmTTkCfNESaY9aiGPk9HbA+r5n25txJ2RDN9PU3AtTVqHzafM6gIzUtQWE5NZ6u+uIRrrQ7Hanfv7DDyQC8mDLHsWTkS7XAszYG1PTwg4rae3zCyWzaFTb8XoyTuleBFvweZ/HDIBy7/QaVvN9sqtZuB6eSBIvxY9RrhDWetxlCWKk0ZCgpbFqVMS4iwKjHzEKrBTXvWNFn0LOz/gU6U9HW0zuSK0jSv+BjR83Lk0OLW6s74HWr1pApnj45WpFZ7wyInrgGlvRjZUFQLOmekfyDOtGerlned+1QjEUbK0WQcA9Qhip/pAh2AtWaygewmMCs/Qy0FzCQoSlN67RsgQVUVwsWkNFUMvFYpnDd3/c4z78VnJbnqzPU+EAV6U8K0OmMx7Bv/HpZJVC1nxQDMmdm87FWR0CAyOiv1PB48wps1ftALLVBAp6Bg+nadOYV4mVuKLNGxirQKInxqOzgy7bdsuE19iE+47DdwBxr01HOGk3SdQR8Lsw0T0u+SiMcS3ft4fUPT+Ll5SxJRY+SSrk1srh1m1iMaGQlhX8OiVR1g8YyOfI7UWkZpnvCr15uILmK9ZVrlj3uNfRzQPWwG8wYqa53IkXpkjAgjLnuN4wsBWOnySl4bjDzlFvD5RGJBBDYy+86yIteY+Ul/S8FhFdsRkckj7/DjGWx/qWko2xI9t9qhJDwlGJmBWZY2dmDTnOiIzTNPBOrIuSFl5kYxVTDGxXkWQiBcc9Oilv1Dgofo7MwdSrM4kEprYOSMSUDatkdLgjSacBExJNz3FHJAOhEzddzYhwLtO0QZYabNNCUj1Jprx4zmxq3Jb9FM7lO7bPjRlkB1Ie4zba6crOIxBybaOoTQbLPmeI/GSJ154CgbVq3wXMRpLYtSzMHcCToj0xYXQdNpCSCmr7MYCiUIiFaGBTohY0sIJAEwuas3yYmHCX8H0Ysa7PCz3JnSmtLsvZRegqnMmWB09u9AaTrmUyTDbByUC5O1Wvv441ES3GU35zOYZUp5OlB7415B6u4cbUSzy5kdGfmQVqfZA4Dt87edvmz7n3tbT+4dnbppNi1Xr+bzNHOH628NcTjqwHOttOslYIxZnZlktezLvNswVNurTK3uuQNjZMq9FT1YCgKZOM3OL21etMOkMuWjJJPY2GFDY7mPmwS7THSSXyD9Cuq4zX2PhYBmAZXcUOUtgwi2fS5Qy/fIS6CRily0bE9du9i6X1MKtH2qmvISnqZQbfvF9639G4gitB3m6tGNaQ3tnxqVZdt1sMi/wyFTGplmhdcDKkHLa939DNeotpQDtdvZvBYFjPP9InR1yeLFaTLJNmz/zbaRhOnHhLmMxhj7HkD5EwxDykQhkYl5yz+y0SJKgWeCW/OFOB2pbQBO12MdKbEFPfc/16gRc17XZyMen2tqmdKUNf0r0RqTkailVfiXvQzMYKdXau8ZRmzg0nlm+ouQvZmqJA9+xFcAO1Rth5cgT6flBrJ0H4Tleto+02ygDiRRl5MzBZaQTcvDQGdWw8yQdlX20rytrNRafE33KhIk8hFOET1RiDnp5oJvpad1e+bXdD9gCRLEHqfZ0p2QjGnIISmkgh+7P0ZaAKtw05fBzdarJbiGDeykbdWaDeXc9CIMSlk/NptHvTqbApq+rXGQU3OpYUTcKzKCA8ys04Y2IqaW2hxczzJV7gM1MgAsYIJWlKznoXSnKp9JayjbcfPjE9HOf5XQCNTk0sTb3ymA3NPO7yHSkRGQpYVvKYDIoCQSCDZX0VJPOmPWJjVeOZwp7LuW18rYzYzCJm4U2s+LsLSW7DZuQEYgKorA/VGuATqx03wq35ae11r4zpPgLRyDnj02VJHqnrzTfm8chYjrs1cEJlT6j8aQisyt6Ijhx/3EfThEKE2IFE76gH4q/TqExIIqbJs6441fhOuCv+ma5YBsQoXREAc2PUbBv4FJf9jm2aDP0DHcU73l19ggibofhc3ExA5zhtpYyLR8KI/O2XPSsVsMmu3cRdljpHc/NRAPvjHiBhGYxbXmYePw0ntAaVIg7a8kHJoxux1wOI+FHr0qQZumBRAh3dbKXYhnPVZiliItufk5vtBbe0DPDFE1L4EpAQ0b9BXEE+Xux1qbIikzcicoWDZh2wUlbCxCnQYoHDbDL+Go67kXGqkU50RD1OhWJkeEXWnihNDtNi/9DCKcfK8yFPPvDLWXpkttP9tUNvpeGlzejljwlElEEAa4HGq6lyIlFqZuEHdmJVpfdyK41kBGZ04kiSre6g5N1ZwomoG6L5cNy0ty3Xojn3fNnhHp8ETtg6MXhjFsW/6UWn9ck6+HWEwGp/DbICOvJ5B5ddHM4V5IrDaBgbq+BEWtSZ9zYAczJ0qwnF2KBZJ3zA2Iq9JBlIwijz6ZuBUK9TkcqiUZ9Z7sfZTWZUSCzq5EBUZzAWgDjg9xyWVX+RozGYr3Vau8TEFnnwShgLJTNW80hx1jzsj0TIawJUrNsd+H4y09xmQMmS1M/jGD7U/zMzMFatr7FBQg4QHKCxg7zWcBEELYc29HRnrmERh7EU8xXkZUEAwYKIDm3Rpl52S6fmagcLWU80tBbbNwxGZUw3rxHs2Wpa0dBpmv6eMyEqynxkd7XhJxnon7WjU82tsl6WGtvydRwxbaF9IiW2z9GGIiYwZkCSM6iaXVU/iNsZPI6YhK0Zxm9oyxl4yNLl4ObKIsjWbkb0oTUr0pMj+ohYrdZ0VQACGZuDfN6Ivh11YKr/9mrtsBrzRyawJjWHUkL5/LwA7Hg0UFqUUmoCHCdZyYnnZ/26EIZ2aPh82hHbMN3tIcphQEDr0eUYJmAtDROOlNDm3NUmjnJPV+TW4ZIzkZUagekS4TJj6/DRlVKXmms88ZXdpbjoKv2f6On7cBP5xvw6fJJCzdl7nga9TbJKFHGJUVroRqXoIi56SatHVpdflAqCltQBPUWaTG9PvsUO7yj+T3qaXnCnDamQSBwS3DeZbJTl5ICBZtDCOM25oqw5VbsnGoumucREQGIN+BhKnMhjgHZScylEgT5MeduVAak9+GBFG1FGxnzu/J1q+QKTMkkWYue4f26M+cHFMIlLlI30XT8e6IBr1EFhEFYniSJhQjU9U2r+hSbNZ8YxRyKgCT/4Z3DjpWGnxDEXFH7sNIcZG+EdBxCnjbLwqc2WtK4NhhLOHgtKVClnPW7BDZjZDnv3Iw8qEG8+vbgukT4KLm3FacjqUIMpO/YBGcifVX0pItAzVQeKiRrbFlXgoi730k1xXVYKUkeOzZAAa1STKfUtajLLfsXdT7TYgQNW0qcBVfN6EsG0uNQRRCW0rLar9y7dLoC5gXwveDuR0clyA4LLOEAuFYhJYCUQIow9DKW5AZmKMGqRZTGAghyMZOW3YMOAfyisbTTGNvzJmZf2RPOZ3YR5Np4Sga6agvRzxEl7MUDGqfh7jXXAMtAmAjGPd6KIHxFEJl3rTWjE6/TS5EQqDse0ZHYAx3trwgmWqjvue19mLUECCpYZqJQ+E79J54iOFuAxj1kRJtZqfmnhpA3wTXqrQD1LqS0THfVJreUIbOPChpVx2kE0FY++5I4oSByVs6iGUR4qC9H1mgaedTsOQDFORFtbZLaL0ZK2CIDaLQWMNcGfvTCsW618Aelp4bEQJS6Hk5292zRfxMh3L6Q8ic9HMQxi27NDkdsIToZunR7hEGYDPc2JO5bEgwxlAhmkUtlDetrkOTLLNbja+BAjeRhQYQQSHXQjlH2d3xmOXnkDBwpvP3Zy7tS1LyRDzlA4g337zuELQ1xrC9z/1gjgNNlaQlmV9kJgoIYXjAsrLU59YnQsRiuhaTqmaCqPTD5H+ax+GRMxQfKQcez61r7EKI0N9CHWSQvkZj5IX7S3NHbk8wTCn9oLstyHkUKKETe1hl5HVdoUJlsvJWFJAhcKrNQ3yWdyyfBH8606dAdCS95KwSd+ywmNVEsPy8nJxoRVb5gBbCxVdCGd6DmgE1mYxEzkpWEcasEObMA1EKOCFoQwF5EEQfMISPRWXxWa+QNp4kdRIfTSNTuz2kJi97zgzVdFdh49wTpbsDtCfLydVMnUGE0nwJlkTO/QShbw0MlnABULNRGuMk9GaaspkB6Xzug3hCKKLmjVDwpb1vKJ+TsmGJZIg0vOVodDMg0UiloVPjFoFXz84SHtCjtCxJb0hP5lKD1fQ5qWlx0ghzHAwp/PJa8O1ekuFHmCVBEy5UUAVcGeFI1KUCNdCPUOvxdl3QdKBk/jERCEshWyhn+70qemOtRiHzHqkxUCgYkM2FlT6O3NfNnXv5AzbCS1msEDHWd35cAVkKSIqXHbJ0F2sLBbI1njIpJ2AtyCMAkrbpsqSg89Lah2P0mWA3LRIEu3x7NuJd8vCPEW0I3qWZs3WA+hoDhUB7rtn9FQ3xcsLmptrupJK86D0nY6/FtOrVyE5QdHwdzsAMQTQzB8Oh4Ud5DJ6T03rqszNESphPoQaUsKEmQzp26Zz11rtTZkY+QzKHIgL8XCuqczmHK4xaU+777NFkXHUEmzUyst07HilRTK5JHcPWA8ZyCnoFlAOQz6vOUJJBawMXo5meAM0D+BFm+6bZExY7EM2Mky7TDPPJ/BGmpl9gIvlcGrLo/0qzbU76HoqptFcKXeaZqw4mlRMyg9YJ44nZJGJ1FjQ1SjAE3VYEI++BRnsb4eyb6wVqys9ZJZVVp63mOEY9L4hEAGXO9qd2TOzg080seikcS5Lbfh9/u8NO9sGEx0xqSmeawYD9qA7crd+lnZ7UPguFNRuNEJoCd43DURGaJWo4HKLZDrVki9PXKeYNRtj5trvgnVff0NHMlnx9yVbqh/NEQNHGztcp7WuetvHYVU7HpX22B5wVxQEa3K68EDdOWwNkqtAXpDaEhVCk9Vv37RoOTTt1hABf12gijBHjD6cDI52cOU5RgmfOGt0AJNo61nmMvRDjWKIJUXQi36UvicJpr8zN6udhGFnqTq2qtOWBoiu9h2TI0Qg6fR7zUHvRSrGJVKzD6BHnVy0WvdClMT8iGzElU1n6fDxNRUV/GGaGgRPYFD1ywJZTKG+khVSr83ZFItQxS/kKhV7m7NXdcfZDA4fo57gQVu2M6yuqsS8FdiGlLghi3xbda7Bk3tkgiMO6oLEIjokB9rmIay22i1a+qii1AeS8TVVvpvNRC0tzwMkYMxvVEFHMGcKFnatYbNaiBNpl9/CJNE266Tg9V2BJRw19KvnVOqwJZTNS49PkoTOUqdXHQxJv88qzdd8uiTLzL9TKj+MBGM2Ys+pcaBotBswjbHeKfrqeFbsxk6XyOEJrhykTzsCY/KZOY3RKttEJuq4XzNzMk51sJ29CO4GqMwJ1PMdYMqyHNMdm7mNHIUCsNZGKGRFIaEppNDqrM4kqhMsKOvc2cL/5rpzPyoQyB3rqOdvQyc7fwPuGctxDicRGQ+apj0QjNF+JKJOeMOFuOfmx51ukc9IgxCX/Ds2fGfdS/ceckYbenrFyM9Jsk7nmgbVaxmYl2oH4qPaESoImnNAFa0+wQUfy2RB1pOk6WB8Erj3vfSG3oqIt8ffMPhgUXA7Hzoyj7tBgoNfh9WpRA1gRGsOKU4rtW8wfCEJyVFPfuebMib18EBFKjAeCQ81tqKUKoiXBZMu90sBFNDVPxKHaFfpAuLZjNqhlDJ/DhGgTr2sL7aajiuiCxDIQzwBUyHahXU44itQwSM2fMyqWPdyYAzI0hjFa8rOV4Iw+HYli+iAhMY5K7y2Pygsp6NxGaT+ZMelYU9l87o3OfNZ9FHLldeIsGJUAkM/chADNgGRcz/sOhsBpaqCcycahRM0RKqzuEdUYzIDtfgH5H7aIjFqaioQ1PNUHY9beoMzMPPR6jWaGMX+hhAprUWhOVSesOvcadtQEidAj8ho965g0RnPA5UjdzG2VmVJMvvlN3xKYPk8zqJtjNA+tfReoZj7ljuUogahshe0c7pYj7uxkydwA+gzy4SZ7WhzAnCYymbIcs6FLCA5khuVBhNcdhzDWVeQmsoemYH0zEzyXtCY868ILqaW5bitGUlq3ByEoldsza5Qhz45CNqHPXeQgSEuwSjM/kxCcUhzOkQf5HhlOzHSEGHY9BztNxeMdK3pCBXk8FIFymI2ckChBYiPpcIJT5WLADrIGJpmLTGQjGCN7oW4aA/VQbAoyRj0s6UDoMDtKScAxoqD8ldJ2Ev5gP5IRIdCZc13nhLdpZqUIZmx3RiF05mRKVmKSCVpPzhAOoc0j8NLHDSz6DuRHYUiZEY0miESEKYhNd0zBgVAMQn9MxirNT9Q1bA8K124K8KzjdynEvsbKhTD1niBCUOEiji1PhCcXJiufa2AHv5AlC316oAQH9L7DfeD8oA3zTas7lEbJaeXsyUkBQoRAWxGE8mbA+VlJt2HZrLd9n/CX1yIh0lzgItxzEE853gI9UADkgrofQNI+D49t91DSFuuaZkVcn8wJAJxzQgYyRU5IlOV8peS3JlSqhNw0xEj2tpBVDgpmBSvNCaKy1PqWQlDTx5yaK/c/nVgaP5nMJI1qOayH685xAMmFiRTKAx8PaWLmisxQE1sih4SvyhhFTWwD0WefCZKRCBKhnIxhNrF9v5hzbgUXkVvvS7lpjeczmXLyECPzkvybdnohoAmOMkBjx/AzeCFAXZ+ILeiqdLDp2jxzs4Fhi0wJaWxGFxLuV3r22u7THKetO9bWMUm3bjcl4r/BSlJOssvvTo0o4P2acNNVM0xq5YOjeRQ46eQkvOv0E9hIZsxFrgwb5SYZMrMRMSOVk8xoLhDeswfFTOGzS+FgozR2rwvRxqIiDNR0EgQjEaGVXwHYVKHGWACmqKcgY8r2Lkvbea3Wls96aBe0VUMay0cgs4DoByh7f00/QRVUwWdoAAqD42GTyi0hSwHrIQiV+sscFKMAyzPISV3ViIbIJQUS4Sw7owOh/VP42jipFHkDqn9CPXdbRN4rZ4Tk8xehpQnSmUthTIZnDfBjaDmVd3eNVnvcBTzRIo9ZPSmVrGYIn0lL4GNkKElyjHKQBjpjazy0iFNHu+1Mwm7DpoTc+F4JJoPJx16mgCeMP6bwoeApYRAHG/cvf0OLYMjByXtD6CNebT43MTeb4QDVE8TbdV3335oivjnTLqwmYh79kCOPORLUlAttO8BGMBPrJ0i4asnvQUR+fq6zDsSU2gsuGx3w7ENBSF+mSSCX9rs3+tVBNGJEarPWF0IagR/13AIKsrV32IY0uIhD2gyhGXOKWqTAD/07djEhNJsAo7Q6n5cRCcJ6CqvK6DSog7qa6DRh1wiwNAjquhvtRWHVwtyZcKboBT9L5uD38jnEZVQcjA4oIrArgp3HjGIV+epsuEZpeubrzHq6RKZxZoueq5/fxk9Bop7hhBZcN7R1c4tir7x3yVaYuFKnheLISE3ogMIJaIIw1jaFhILN4vVkuebEJ6qSshHKyP4eGwHPc+Re1jri1uuFz+Q9sry8dihzI5z9NiChUiZGoZT6IfpLX03+/8DA9IkRk9NDA5nMhNRKqZVl/7AFPxnbPTShR7jSTk4gD28yWdBdMb0fDhd6b6KcbpS2wMasMM1FzUNtCUUmQZH32OUEr6UKpLQdSqdOQcW1MxycOD80zNo0N+RziD22zfNrtEASe5VoJ8FlJCXGEDaikZA3/VPX4doyzOtz3b6nPUgn6aj5nVovBV8jhhrJeIy9YR4MiJpo/zapr9BqNbKJc4h2+9oHa8Kd0QjPvVN5t+kepBWxEJUQUjl1xhE0LocllUNMeQ/GpBCqJdce0I/AaEZnOjoTZfI04bJlqWSgEShVolph3aSBRKcznd79FC7+lKCIhLih5j+sYKVp1D+XTC3ncbF2/4vXCUHKNPCtmVGoovbJwWwZmWVOsZYE6aVxCNX3e8jxk6FQs/Yw6USCo6Zy+1QmJqMKAMAmvT6nmu+iL5AhOYeGKId2LsEloSFNmM/PXp+bbNFEAbt9dcmSCcB1owkQFArIAciC2JlYtMlZ4Nb2tnlZDyHEYlYIJP0vFygFQlgZjg2hgtLMCmHOErwUCmQiCno16kmt3dvlGz/PPa9YvwSEjTRZ4jzi7JuTkntEIpMQnYo+aE3cn3TmTfkIeIaI+86o6XGGNvkdETJ+zPMj1mhUJMUAln6ayiAlfaEJEibh5Vqa0IUcpelbgLUnaVpeyj8FrJXmlh/jAtLg+imciES8RWNYEGYSGDQZ6jeITjoSSCElf4X1z1dUxVECkQljowsldH9J8fmORB8jA7FpaIPJDj8AY+G2z6SjkQTnLvu3+iim9KcT9PQkNfgoiL2uwMxJU2bAbNqah9rLoeVY9fqcRGqiISIFEhWJdnpGbQwwzzZ5bVoa8xvMqsemhz3IMJmGJg02tcn8k2b+OFPbmc68O4lU8ZwaP5ApxN0xOz0jE7V2DSrqTlISp6eG4b0YClzpDU9NRUFLYZMFbbVuVKhapgMgmzp9Do6e52FKvFMOQTPbFGoFYu1zBbBk31NvAqUYSg1uSJituK4yIovJukCIx6xBPp0xGLqVE5I9QDObtUdqlAjl3pjF00Ga/i73vHU5ZiPBiunisWfDdjCMjNpbMV5XLl5rq/VUUlkwefqFHKiox5TpUo5SomXufQmheI5jVBOj9jRuQ/TYUBcq7Xsoe9WIYCy6e+9aqNIQjrolw3DLEsjAgEqvNh1ohVhHO+Sm9ekr6KHEiRIomZHox7Wa2+ZGSwMdj/Cx6EDhQ0lIscCMTtCrvGnvb4ieCkzEyvsuIz7OBKtcS0HchHeTLIh6fq4bSF/GonmrPtfIQTgcEPNjGSGgNvISZipLzwzYjHrAWJWZ0RqrCkkAWQcTDlMsO2lBW7L3h2fFIwfmjGxBR1RlS2R7ikhyiRQe7PSk9ZKok3hlQjCtOdYThWZ55kwlJ4/Jkd1seK35qNsoNMywMJJWqOmdz1NVw5ZrQtro5qErC+HEmswMbtGvoZAPo16k6zpix8XX6H/h+ayZERnmg3usYzJaxWs0gehKfS+hE79bgRtlrzQ9MP0A1tY4FuVhjNZoR6ZD88GUw70iUUzvKuFQ6KnWTuErYeIDmR3LQcD0WzggOL9peMIHcbQsPqTWaNBFHvEGSflds7Dzu8NnX7F6ZSGmpoemj7VrIJ8Vlr1DyfBrmTB0TvZSdf6s7fNw+QbCNqczzkrwNDvYaVJYEDcrS0XUkx2qrQQPQ4GEukRdWeuiZjejCBEO2P4ETEdW4hZzEtKuVzLYrHwSOQnl5OrIbd1A0AppI5kKGR3qULTgN6NQFS7kR0ozetKI9TNndm5+QY1m6ERNnwx7g1o2nUliTQRXTmblFjTE0sOZG87n8xJ1oO7L/SKjCUWDgsI3e2G5D2h3EGynacM9kLmQaDNNpyCPUe/r8wBDzry1u6cfAyDTa3I6mhMT7Vza2uPVLZLoztXKXm0IpO9bmEIW/dKzD4QfsyVaQl2iCxaLVSagQ5mFzDnIz0dGo+dEdjJrfl+JUklkY0gAmGpOvL7HRY2RCV5epokcnIs02+a7zbbX33LmtWdwj+t2fwsjAb1LFR1VtMu5pfINMMuv1sbs12rc0w6RWh4oHwFyHVwbO0Rl0lRnJpDYuD/6vsVjIX8z10EmRwoIrqO3/hM6YDo2MwuJBJg0VGgnMltz7Rm+JXEqlyS+VOekfUuFAPoPKJSCeTkb1pRS3Rx9GyifQsnamYsJm9NV5xbrrVLyFAxW6d2wTE6yOLcuEyFo3kLgyTNbkyjuJbZNARAkX+eP9tkK008JlHhCojQ6Usebvi/kQMFH4QHuXXZh1+9M2cq1Mnu1EukcFT6NQjLQlgtCoQaZwPlaTDdnwOpeydcTtAQRLe16rsPabAlADXHYAzM/45rhkZ8hosjCJ6bqWk/93TBhu1/6GwoFefw9uyec+0EBM8KUsKjjiFBiS8ltROXmYirZiszHGCiBu0QxF2tL+FkHLjSjbbkbhI/7kzhg1rMoa7IAYuw3kURb60gN0czKYJBV5FMRjUQ5gf3LoZvmBox5H0XwJmbLdbJmxLyuTRpCnqez+W1562OfKdiIyBaMXU3Nim1ntIxChSxAwWJbJvU414p+9EgChADj38dicgdUdMVnF505oOzG3HenImCSGgVGzBjle3HmgQfIgkQMyjsBoo7DLIcgFzPrxI3rSpJ1milkHDI3n5dCjHtWqJx0Fg5WVmnnuowomd8yDDcPPJsl3W6WpeIkIKv0aiID2s0XGuWImJah7Ma4doVJHYgqxyUiFH5+niZHagUJENNvZi5uICyFSWO4eKbZtFBpS2rFchxm0ZXS2kcmmgXRDB7+PJR2pzDk57MUXU1vdycQI6fpczFKAoSj1FmlS6RDQSEhSLt+6v5IbzvaEcoeZou97uhNc8WP5yinIZGTxXeSsVxOOq8zMwC2q3BqbHD7d4P4eW82XymFks86j4Clb2dt83NtQe9wTrNAAov+IySKEONbO+OJ3rWKDKbz17/J/MkQqG7tqgfx0q5xuSl6if0+Vtl+Q346czkdeT4ThqzzUXp3RC/cIixaWKpMCCXV9T1Gz9iEBG+JzqnPTLbyc25LCalCGz3d23Xd1C68SxxfRqh2GMPLGQlgHwNqqycEEk62i410vfS2aDOjII6a9EXUkujD8rtwRAo360iA1Lxt4JChDrincq+zXqeJwxg3UYv21yvRiZCd2pCMOhpTZrmztMTIsubunJX5YJkGH9moG7jNUKeYs6Cwoif7vUKh7t3kSabNBru9kMxZSZpClDa8HqVSSgAAHwdJREFUqzzZlWCIFlJkebxtMnWLoRRe7fkvGydgIpeOxKidfEKjEzcMyvM3qEENy/y7/4tnpmO7AOOtoYx8XQzlKITUf3p4tdNC3tNApFsCth5gyWctQbNpXmQDSE1cIyzr+8WATainsIkScE86HACL6lo/ieoen5du16p+GgD1/vZOpPGMwki5TERz3hIMZjs6K9tup6DQdvLVeGFgTho6+WaDdMtSIVWrg6ETNKIogNrjcYHZ/o15G0DCXU1a74jAi+hURFT32vgiSMysUZHfg/4IK0aQc5MMgCpfpwOxb7XQVCAOawJUDq/0TchH4RVSVSHWRuPyeRJtsdiuddPyzK0QM6QJUPtTQqYyHVE+iMwvCf8BzRHK2innKJ8nzJPujGuEaLnWxmzlUxi5Lzl7dZNda1CZeIe99LNoTXVZQf0uCDbIyiEfAs8EVRMB+opSq8fvHgHJx1L7AmyYcENjSEbDELn2ztvl/MzIge2amfFmRyoyWWp0hMi9BwDWqfCgtC/bMwdadIP7k+tnLkXbUq3xTY5Kd2wdtHV9aF0N4/T7oByhMQqgIxAS3W6XaIF2eR7ibqkLr81koRAByttPDUni4wR1og75H1AJXZPSNUuhqenTQWaDuRCjrpWmgA7fMyzHBiAczMzPA2XWzFndyKnpVF1JR1O+njkK1X0KoaXaLJGgMWoMNOLNz6cfQxqI5ko6DCffI8xdo6ai1sYK4GoBuGmtRuE4lo1fROsmQ036dSACiUelACdNtCbKSKE1mmAUYzPcmo5QMWhzXspvEQQ8VRwXTDkprB1lYiXjsi1g1ZBgY3LQP0E9OLLfRCEH0mVqVtFOCIpND1Z+Ph2kTJLa2vE1JEkoWHzeC8IgPwa/O2ejK1i9l8hF4yJQpuZofULCzzAvrB2wZpZ0ARZ7RsHWRUx+fhM9SYGhUYmgsrCd1FBcNSIjzAJk9SlmDjxORjQPQhwMG6IIikyZuRolLT2jLtYOKt8bi0YDeGoiwVXB7WKY3uAlkFMxNxwxmBg7aBJaRmNwPFYjYZoHGb2pXAtGPVyvOw+Vo/e438cVvlCbJ7FQYPZBN3QAI/1CZFYgnLgNaZgtxRAzIjEFEfO6c1aau7uY3MaSSCeFxGAy1SwU0aeg8bq+hikESNjGHsxiICHFUSYqEQOF/kyhQVjvQOVrUHMlQdqIIcDK1Mwz1xnkmbMhL4bOn4ixmCX3xTpdVQ6HCt9oAohWcp0MQ/r2d/zbNRKSe9IjVtTAE8DG70P/iUv0iAYiN8NqjxhaRV2vK38T3VMgowm26GlF+5Nra7gC2xA4H48Zoqjz4l54CVh+L6Mh2gUoizI7X6lNvrz++eGeDj6odS2coycnG7hfpdgpFCzSv+XBbYwSz5FZf82ZqcMyQOV9FBQkWmkvlMZYdk3jDNWLBGJIuS3/AuQY1KZSCEgbp8akPbskc65t6E/6AGgbq3ELY/orHaN5IG2WiFMIaO2lReuQe5gRJZyG1/4wSuXRF9OWvZyt0RvC6szjxRCEG2JvAhgpPHUOGTY0yKnM4i7j2ibj/3yW0pZ636GOYWX6mBDgm5rRbnwTZKgeGbL0z7i+K6d2XWSzB5vmNYIG5QhkJEPmyhhhhrAPKeJe0RavkGXw78gtXGtfvMKRm2pW/WxWrGfmO31HrP0jkg6D2UMQLJv7bE2P+JkbJ+eb7ydBnH/VrFOkFJ9epgYJhOiCnZU39nRqybHLFOjKR6hS5oJq3srJ44m7KbJGtStQCEWL9ZR4+azO/AMDkNGM3V6vcSiQIicDKB+Hyea23tOg143QlxAPEERI5yygZyYyUkZpc8S96dzXi7NNaw9qBMHcalBqwJbIFfkbx811YnupzTvzIUPCSWrMONUQ5lq7yKmHDTMMblo6k5KmUJDi8nOF2wLTFwwQ8eppNkzvGq8IQMKlIRB9NFEEUQcyUpah7rp/Qmgy+eYsKiOUl+yTxT33LpS0x3vmFzS1Q74Mvd7jDHG/AhgF/bemQ3xPbQjTz9BNC3bsyhzOhgLil6HOyi9k3Fa0I5BJ3KfSHuId5nDwuvFczXArpQ7DTnYnlenpvnWHdp1td1oBiM8wxNbyJQSH2IV7bT4LWAkDR6EKZczlNdZZfoalwfLOfTww/ptIhpERls8DVVg2RvlZqOWYrKW/l5o5wWebE9jtYdkm0I+HgnAypZgDkg69We3stDe7NhoPCGE0tolPQkn9XOiM1RkAjPEXGgEM7JbNArgFwFroxyPCw/wJCl0Oji54Du13i/KDGaKBnEeti2hnqT4bPbZ/sVqS6eJx5TzXDIGyo1Rcmtrd22/a2Tx/amzU2tLMEeO1BDMpuNEcfVxD+qjkH7AdIg+j5ZoU+Kj9aY7MSjDj+7kWB5jDEWbGhAYOVTOMFBoWafs67P6vi4lpM3+3DGIE0qlCuDfzjxLudMYlKJBsXGIrnmUHwCLZKu1SdvROc4GQtsJErXBGCGNq88RkKKL34zlY97CB2ccZDNTmeVSX8EIcJTDLsdgPCI68Rn5ut4RJxOzOFl5ltqlyE0bbSPkrmqSnecBwMHNSFIP3+jyTm2AhMxOa614JdZ0MlA5MwApJpdZPkFyOW167CaBAUUwiGxIuvpYQAgBVvxJRUPCkcNLwJiEVCpJsz3dRUOu1Blc3qf7etH0pg9jbtUzTNAeR2Z4bc1TPkpo9hUMgzA6vaR7EPldRFye/t/wNlmi3sPAma1EzSIg04sydGKX7OciYiuYQcUX+g9CUzjzWRAGve6eCq6I21BnoOeThgHJEJFQHWD9KQcFrxx0XeKLQiiYRqfD8Gk11VLc5DffyWcALxgKVms1xeccVdnIaGYk+w/nZYDtTkp2OTWonVmlaa6ixDJWq27FnhFoI3HVW6NMzPq/wY96QPot0+FW7PgoY/s4ITqv6K/OCsLIhgGwt6MzPJzOLSOIaZkvMBT2eozv9IrNzTedi1qyw0pMMzD4ZvYRd/olEa2Q0OICl0A9BoJv8UKpxMJRDGADoS8g8EPN2P8YIG5KoNvIJm+cRY3cCXznYJrU9aWTW3nTnXqAGnoe3c4kuVWh0puvxuYVqVrhSqikUeK3m6G5krjM0A5vllgmbwoDrRjHG5JQzFp+h04cOXciOkbre0UoZxpkApypSmtgpGKaU7Wx7ScamQKs9i/6rszKis9FNRTi49nzXluwgzmzTqlit3AwKPW9ChThvRfTorEQtitxS8wxrGqDGr3RGjgXY56ExJVzwOA4voO4aJexyAuYGEwbTSThy3OCCFkpFer7Xmla2C6FTMAo1AAmMukxp5E24lk7MgRzBmJsqDR/SVfvMCItNGJPDYDVqMQmamkEdknd7ITAlfiURhNAcihjpR4jGeMISrGpMLNPI29lY7Wt3ghIwEjXMaIBrWbXqFglf2+ThrPFJc8TYFZ2RhowuyATtk7+SWJmZaGMnbaUlWusFkiZGMBPvyU3NMxcCo0IYoZBAc8Pb9fIajA54anT5i6pGI/wKFCLcNxFcRqKsnpNsQWYR+irfkBKnGFlBaPAyjehbaTuuz/K88nspQEaew/AoJyjhhY1Q8FyfBF6iL/YIZVcw9vX09v8URkQ4DJ3H4KbKq+BneUdHDAbYydY/OYkNOx7l2KyszXzMmZvNw6IDdDhslyBlWaCy7m73y2mXW26IgT70j1CzUlC0nAh9HqjZHzKBsIXcQDJji8mTEeJ0RCvRIi4FoMroUwtQK9JrvlbICulX8XxmmVbJ7FF2Hr1ANAiGhMwaETEmE6ea4KIQlE3eGFmQPO1hG4qoMEqiGSjTYAvPq8KSfF7bxSAon0dBXcHzgg+g41Y+DW5g+ndoQoRsCy1uGRkhgDbufZ90Tu07dmWq9R8q9p5YJx20oOAzk6cgIUiGJkqKhQKVYLeTKcR1bmh981qLcsifciGFXoKU52LtWQ3Q0KL+fF57k9dxVZUC5Rz1zXPQuVtMH4giPtlNGNNr5AVmS1ST4EIQrtOqMy7TxrHz8/N4WDoivZ7PhiUyZuq3pWNopBMyEYSl7dbDVF2ocNOX+F4MUD5sk7pYMyDBwcOybBI7ipimq38E55IEc/TQJgA/1jORmdugIj/GWAA/nNfa5ahk1CGdQN20IkQkGmE0iI5Ir8OV9lb+xEQNWkoCmai9aPa0umoxzOrttWWv6zgAa4Qf+7WTD4VTp2RerOep+Sts/CYo35oBK1Sq9PTm31AqPqCCtWQIJBJl2DzqQlbB9vC1pEAWc5WScWnj1Jzq0cFEpv47FZxW49qyABTxPDRpfc3+EADK2RoMWjqtobuGBii0e5XpxToOgEKCZ06TMiMcbNqjMnnXukQbiYRqwNOSaySDE4EgTaPKJ+koIp6PtU80UUr/1r8YcYnXBmgWGQzmA2bw80Me9lrSlt78tgm2ZDUpbelj5k9QKzNPQaYBPeajGGFZSrDIfiRCoM2IEhpAOTz5ulnMUQW2BWXLrkykZcnGwHlN3o/FQ61lXVwnG9qua+WFAOit2bQ31CTHY/k/2sQx1pmIWXhvs0ILPYeCgsy4vmX7zLKnECZdflcmAUPMCI1nm94cLFBrROFIZkntRSGn825nrtqNJNHcN1XK8nWfmYNAzTvE2LLRiX429+CZW30W1oQQBfNA9NrEhhYqwzJyelSWnteq6EtjWjkTp/ZR7eyc+phnX2sMobXW+V8YS1BRn22fy762apvXaAs0T1Dr1+tQNWqhAN98V+XyYp2lXYNH7phI2le3L6D6fmzFBO/lQBaSwXa234Ppopt+FWT0tJery1JSG4ZGHRbjY3PAMkH4w+a4yZRw5DyRjGdrtXx2KwYafRMR2oiXpkYTBOdnvP5jhikLy5jpuPHAk+iIsIba54nxHUG0cw3bUuZV2ZHUuoKqHcJ7RU/i+kUUemagCc22tyoki/Vb31tbUp5Yy+colKPJaik8/XiA+pIQuiuZi2giCTi1oaV5V5WRdeZCLVy31pPa0ylokCYK7fHu6YeQmAHA2OV6y/3m/J6cvwAL/kqxFT3EVo48Pzo9K81c29dteEVHks6zQrQIMwVPN63Zcr8xmrVzZdt+CbJ6o1bfnPNl8uUz8SMbPDAaPTQnvfBVrhuWZs+aS57azUoIi3URZ+rM9W9g54dDMqwBntqQGYswwAqSMzvOYDE4eSbTm1XWJnt4skluTwUeVhmLXbgI+mYUJMcLUOA4E4aUut1qPbLqU/ewtsmO2GWfUK9P+RZSuorQ6giU9+FegojCi+X0zvLxOnU/nieqCAduz0DspcsUuKFpSojEPmb27KTfpEHZ1p9S2rULdkJtIHNFgkjZ+l5OK2Zb2siICgkqGX4G87AGJ64BmTY2kZ/Lsv+ZfpqxqxCoWRCl9byLWrsYzz1S4Ft1LXzCW1RBSUspZFU/08VMtwJyL3pvB0FwVUo3YQLEHgs9cB/5fgjsQihFZ85ycK6PwrmdeTG466+a4ZH7RAWDFFp8Apml/FzRqVk68b1nWnrJryawVNJuBs/MUiOKsqQno1lXCWIj6XjAfGfLYoq/mwGrw9fzSmTqRVVEHjI5oJmfxnDoegwY3EOO7srj0KF038TmkMkAJLqUdnNWVOD8TFtDjbVxvhFJMIeDk8OJeHiadLCSaHNNtnjNYbVgBhuogq+xxEgD90gaG7v0eyRBzaP2zWWW0bE2Gtoi0c2khVUIqgQFanDSeiwGhdfAIjk/0+mVTlTjPlIYCbkFbO1l9T4PYONgjUBwhxvPfM3Q+oR6YfAaviJS2+nbSiHLAUluSdwUtBcOXYCsUA3f4DVnzieJVdAZTMZtjBcHhW1fk3KcxuspmNIkCL3k6aQNFyPRhzNfw0c5gq1nRDIZKs32PAemXEvLk46pBLvfRyxdqGH6saGBFWygy1yREmYdRQDduWqozFmGWnuUaCKvm2aWpXIpYTMxU+hOX23HugTLuaZxBo3AeLA5ZChCqUPwXc1+x0jfRyMI3nXsYDaLCIgCepMUJYChogHJ9NW4xqulfwcPoxGgt+sqJDdLG4hqrJ7PlghZMuy1Zggv2wnasldlqnIv+oTzFHARXcnNlj1tyZxViEUtqurMTcSIhEY048Vk5jn8Kf0VMgWS0MloM3MLrPbRuE9MIGtaMkBT+oW8CJCDlXzNJsQUIgyV2og8kxQEG0Q9liRs1L5zze2spHXzWWnGFIPMZo97HT3vB0TiXL8WhbR39pNOb89L83AW+sksXBX0ibfydWn7QCAj16kzR+SYKFRKREq/h4T2VrhxZXzGuhay7qTEgjYBtW4ye2GKFmVpSE7Pbh4CsOBc3r1S+Ht9idnwHTzdLdNTYEQYVJrWlnRistBpKelIsyNrSjQZ/SIh80eJMb7NM6CJQgJfm8QmAzBV+9gyHpcl0mIVIm0QMR200iRESV3bcjOp2dU8JK7pCL9GOAMrFLvp0ZBwX4V3RA9rromOpIbQgJHhdiK3vkcuBjYyUYPpFU7jo6/Vqp92tmo0AIXrZppieXZG7cloiPZkpk8mojaBOC+Yp10rUsChZ3H05ZT+EwOZNy3sbR9qDyiM4DWTVNpagj8zjZ2sloLRKk/Gc1/of+ldo0AI3mz/uKUjW78Xk6WvJG7r2o9yVvb98HYvXthSc1/gCa25/0HFXU7Ijf9D/rAiKSWFwS+sMa5AQVIh8kIjQRiFXEqI83eEc0f3O0TL/9oA1VaYRdhTvoz8OWYEgMOF3dUBShreHX44D5jOORtzVn6FCBAiHtufqGoVZqSLuje7SDliDisJb10r9yOb1EAzS5OZJFCo4fmsyUkjY9zrMYTnsHKGJiHDLBOtIhFKyUJJbZ4a0tc1zJXjQdEW1S4AImA5R8eA7dpUNyPh8KCnUEoJHqSJ0NK4M+eghgCj3QfSpICJaRVr7yiME87ambM9XF2DjkNGE7L583pADWDm51PIdDoiZB77Fj3jWZfoUb/KXOOb0635PiMYyRFObcp7ldnJfytCo9L4kQInby/mZ7JfZqJKdxsY5YjfR5kP1X3bcy97BCS+q3th81bcs1fu6v28H6aeTZXTea8tUkm9lkjPBbkcEhC69fb54lOx3h0sIgjlswiGcqAgPxmRTh1mGfYoxdgX7Nqxl0QgAgOAbP2vqsezM5XCF2MgiOoYsNz2J8XE3cljpkO0ZSkBYQalhKe2j9GEeeB9shlm+TK6VuOQoRYZKMnOSAb9AlYZnrwpe5ZmOT7Y6p/MN9fwQTgiqUtHGcLLYdqjzTR5wco8D7A0PBiReSiRR5YMTBf6zMQqmgDpYyqfRaGVTYRF4TW0vAuiEGRRoEfPBiETzucAhrqIZTbo8SxQAplT2pT2/sBYTiQAerWq5KZDQkNZFUSpiSAiapOMkM5XKoyOoLRMp0OWTEnbg79aTQkMhl2j16RNyxAmDEyAY+KcBMdGmxP5pLkkP0ib1NfMihIu9Fek78JMDs6RZq9JmJTwIEKIZCzSNd3EXUC0fWnNcswsJ5LNFjZbFviBOQMpEHr2YBaaMcGqul91EyLXR9NAxJEQm448MmlPwkqtKM3S7XoKg+mV00Fbm41TFA0BlJDF+SZOKY306uf96czNdGlXjkVC2JGDlnKNVVQney6YgNosG9GIF7h2jlPICEJSev1NxACkoLDSzKNGJaiAjJpxYS8N6HmhaAa2posEQAoXA4ClDU62ui+1KmsnMkrDOqDajzZOAABsV9qaxMBzbHsm8yrpzDaf5TMkEsl9VWTEZ9jyxjOd2r8wPbrTOwW9TzEG719p4mUHqNmPNHdFtirpaWj/6/tN0PJ6QiYDphqPUBzKD9F9y0HsYI8MIgU2q2koqu1v1YqEwtkmZNFEoWCwhk7yek1QxN1XigmwR8YO7ubU8D0sROYhXOz+ACZhkXmbDbkZidcrOoVOfox/gZtLQTFDKvvxGBELwmull1uaWfu8douqNE8+BrYl8kwLdwsTg6nZyuz0uCahuAjN1GuiCIlHQT9Gpg/3mhimcq/HcNVkJqqqQklTzbwIB2CD6k6GKoHN8Kz5rD0BwK5QSD8LwDCaAUuW1jPUyVD4hqGymvGieWS539SggtKo9yUoKBAMNIUqyclaViZhQusxQQHHcLYGWRd9DUJ25s38/2Vd7ZIcNwhsNHNvlsd2nsquVG53JfKD7oa5uOpsX+2sRh8INdCgpKmJFqfnO5txqhPXJ7XanusPLSwZk1IYkm+iAJk3j/a40XR4VGuDCetIBR2QPhxaKQWCzsdOd1dau7JuO+wKburqzxklC817AVmveXCMkHu9YrSkwc8EN/l2Iq46Wir5i1BX8PpaVZ5OFwfJMXIGvyCzCUDazHrR/UX+xmpb9BqaV3wLdzma/KVNczUrzQpm1qKQ3wHoEn7TFv4IUSRc3YrvyUzgvvu2NSk+CphuMO96k8f9Fetx6BIKD8dAoplyT2pD9Mkec0zsqwvluk09pLGKDSnleBxa9s1xTPKbwuR9oXUDqj9StNosAOefXAlnTarPi3sr23yxkuDGvMZ35TiN1ahakZgxrnk5kFigj7FH4JGHoefYtvvBGW5F0WaK5ROAWJ5WQHLE8z1VCJefCy2rtXb+aER8NQvoygRKMTrHc15ybdI2W0xEk3ntJ2QWaQMTYUR/5pqcY1b1/RlmBXT58ZjXWnT0zep6Vn3u/mfurKsArlndCC70GggLWeannIkhkg2aHOWNGWhi1UgMkqkiKrYzKE8L5DnAGUVQ9wGCEQ2zLTfyvCy4LhCyP8iVRg1t+6/eUN48HJtp4FJASeU/Qq08kZKC6UxcC2pQphqFBED4nw/4X4hkCJoKB6GUbMbx6SaTxyxPoEKUPjrTQuKwYawuVzhMBKGL/q6EW7CVf5bi7M0wTStl2PQqWZBztIsLlzmyew5GaJZf5DzQH1GNos+2WrdDeYnrZjnFxDlvNKeCUPlQPtS+zLCoEHUDgRwogJp9bGqd6AoVPUr5RfdRSxXKviXKqH2itUaPRShkoChzN9Ab35txoFY9f5LmX/TWqWaJiCHFqTG04tb7PRQpn8BY9+PZn9EsfWPeRZIRsXTtHlg124U59i40PCtf74oeFAzmRtT3Rdt2dWmeePfdkQ3V65wIQHkUqqylP7dITJNUBCMPD0vwVTYxlZjCv3ZyCjkot8LjkmnCzSTbPdN+ggiMEn5DAKhwPEeC6dfNnx7TI0dE80n0AWWt6oQUAljdt1AbLV5wpazxDmeULpXsH1cX0D8SrGileWuHolDa3f0c/grH34XAzFRt/4vvX4leZ1d9H2gjiGIwllzl9cSb0YY0oUmAWWbXDP2KF8G5rd/577o5r4Mrk9mmjyI4epcU23DqsmEjkcfVhRpTXJhU92ZC6/cYz01UjfGcFGz6O15zi/wcd3EjtKn7vTJbiGBi+R4R1bmoGRXSGbKVrSR0KC3wRrJ8vVqQP0UQCd5AlonO4xjVnR0NyWz/hajYiL6TdFawUkr3WsiXHFs8wXfzCGzmsCJ3rtV8CoXP7q9Wt6dNJCsBIwogX//WBnh/O+Rayjis3Ip4dNsRlwDibOT7G74CYJin8kXoRPcmp7O2is3wVJu5C4TxvrYu6bA0wh3+ABX3TfSFQ0tl/yTMXuLhIxqLPgrsmNWYKJ+GfUT01JMGn9PUOFlAZWYep05JIc/7yRad/Rphy/LHLNrkPUedTyKuznCgeoOSPyGEJtTn78LPB7IYn3EBZkICkJNQJRjI25h+mgp5vwcqkxMzqGSU5XoIupo8pdvzasNez7VQEZostufxVRd9ABUA7JvimupNZRkDwbjpaToEiqg1mLSP2hcbk0pe83GhIiQyZfQT6DT2evtdadoDkkmrK5tUNjHfG9ODPCjZjX6Sqev7KfjDvvXdnzPkySHEz76sq5yRsy3RjtWuErrOAd4vKgy268pdfN5hUgoxFZ19E3JaJYCLtr3MLxBdTeFcFGT1xe0nD9arzTbDXcA+EIeh+R1yMVy81/N0PMbUKSLImjoN+tTPOT8JOzb1apsqMluQZQ6dT/seMitZEMtKXexKn0TauHH9f80tsJK/VgAzpdvMWUJrXQA9QbHNVWtrEcvYZ1fUIpsxeq7bRFBTRGpEGCZXZRKJEBXZfJB50BsJ4+9nerraPeMpfT7Ysw/E0lGe2X7/f743vKY/L0tus0btMK8H0luzL/pdhZyuRszzXT2neX9+//n1dX/9VTUiPoHrSn4Ygci2h7cU7KPDs1oWZwrYOxArrQjWAt6fogDIHMhDxXblI1nrWrXGuvc05dFH2QMRWUJd9xbEWpn7BB2zWWX95BiCBbA21TFKcJ/zIPfWlhpjS40xcp8EFPJMIKJC24d3rLA+gO1mTTMdsC5y63Bh+1FaSOvdTt5yW5zxEuhEZlDB6biIjJU2Hx1lkSl1VVRpDSerTo5zgP0JrMW2CurlK93GU7CjLKLc3B5rtLUFE1FLFTj7U9OA4T8qZ1I6hOvwdyGSHEosstY8EclQOd0+q5V8Zp5MVpqqPp08DaqpANpfUGt+znbfPAauQ5ykkHHTZElubQv5ZaZ8WUbhnJGfzlD5oKSgD9gOoIhG97H0JJ2aCSBobophp5Fz2doJC0j5KXEMj4RuhkEjanZ1TOXG259PJSXH6vf+5+//AGJrNlbHdTTqAAAAAElFTkSuQmCC"}
,{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)", "background-pattern":"" , "items": [{"x": -626,"y": 96,"w": 2749,"h": 510,"type":"text","text": "","text-data": "TGljaHQ=","font": "sacramento","color": "rgb(202, 222, 236)","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -656,"y": 602,"w": 2803,"h": 770, "type": "color", "background_color": "linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)", "border-radius": 0 }
,{"x": -611,"y": 599,"w": 2740,"h": 776,"type":"image", "image":"png", "image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydB5gU1ba2u3vyDDNkhsyQw5AzKGIAEx5zzjnrMR6z6DEnzDliwCOioqKAIkZQJOecc85M6nDX13Rxm3YSzAAT3nr+9VdP1a5de7/V3kPvr9b6XC42CEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCAAAQhAAAIQgAAEIAABCEDgEBOIOsT35/YQgAAEIAABCEAAAhCAAAQgAAEIHEACiUlJFVwut8vv9/kO4G3oGgIQgAAEIAABCEAAAhCAAAQgAAEIQAACEIAABCBQOgj0O+Pciz4e9svfpWO0LlfV6qk1f5m+dGPPI/scX1rGnNs4Xx445LtPh/8+qTTPgbFDAAIQgAAEIFA+CHjKxzSZJQQgAAEIQAACEIAABCAAAQgcagJHHdvvlJp16tY/1OMo7P3bderao2KlylV8Pp+3sNeUxHZtOnTulpOdnVUSx8aYIAABCEAAAhCAQDgBBAu+DxCAAAQgAAEIQAACEIAABCBwUAi079rj8MXz584+KDcrhps0T2/TXt0snDt7ZjF0d0i6qJ5aq3bFylWqzpgysdRkthwSUNwUAhCAAAQgAIESQQDBokQ8BgYBAQhAAAIQgAAEIAABCECgbBOoU69Bw6rVaqTOmTFtcmmZafP0tu23bd2yecO6NatLy5gjx9msVet2OjZr+uSJpXUOjBsCEIAABCAAgfJDAMGi/DxrZgoBCEAAAhCAAAQgAAEIQOCQEWjdoUu34ML5tEkTDtkg9vHGzVu1bb9gzszp+3hZiWreonW7DhrQzCmTxpeogTEYCEAAAhCAAAQgkAsBBAu+FhCAAAQgAAEIQAACEIAABCBwwAmkt+vQObhwPrV0LJxXqlK1mvw25pdywaJl63Ydd+7YsX3povlzD/hD5gYQgAAEIAABCECgiAQQLIoIkMshAAEIQAACEIAABCAAAQhAoGACrdp26KzySsuXLFpQcOtD36JVm/adNIp5s2ZMPfSj2f8RtGjTvuPcmVMn+23b/164EgIQgAAEIAABCBwcAggWB4czd4EABCAAAQhAAAIQgAAEIFBuCbhtkx+EsisCtpUGEC3bdggKFnNmTC01nhuRXCtWqlxF3iEzp00uNWW4SsN3gzFCAAIQgAAEIHDgCCBYHDi29AwBCEAAAhCAAAQgAAEIQAACRqBO/bRGFZJTKs6YPH5caQGS3q5jF5/X610wZ1ap9bBQdoV4419RWr51jBMCEIAABCAAgWgQQAACEIAABCAAAQhAAAIQOFAEHv046PPrttDLUjEW+g2iv70WORY+i8D9F3Y5UEMol/2q/NLaVSuXb9ywbm1+ANIaN21eL61Rk99/GvndgQTlGD/PmDLx7wN5n+Lsu6WVhJJ/RXZ2VlZx9nsw+5LoovvNnDoRw+2DCZ57QQACEIAABCCw3wTIsNhvdFwIAQhAAAIQgAAEIAABCBSCgMQJCRUVLGpbNLVoblHHomLonMeEDbVjKwYCCYmJSQO/HjX22zHTFp572TU35dVlo6YtWn32w9ipL33w+bDGzVqmF8Ot8+yiXaduPXXSrBRKRWmiylWrVa9Zu2690mIQnhd4+XBs3bxp44qlixceyOdL3xCAAAQgAAEIQKC4CCBYFBdJ+oEABCAAAQhAAAIQgAAE9iIQEiH0myPZopGFPAF6W/Sx6GrRwCLBIs4iFnzFQyBj166dt15x3qk7tm/detd/n3np+jvvfyS3npMrVqwUExMbu2P7tq0b1q1ZXTx3z72X9l26H7ZuzaqVG9evXXMg71Ncfbds3W53KSXz3CiuPg9FP+ntOnXBv+JQkOeeEIAABCAAAQjsLwEEi/0lx3UQgAAEIAABCEAAAhCAQJ4EQqWg9HtDQkR1C73BL5FCb9p3t1CpGmVaVLVI1d6uiQ1dB9kiEvhj9A/fn3F01/Qp4/8ac8WNd9zbrvPuDIfwbeqEcWNP7tW+6Ynd09O2btm8qYi3zPPy+ISExBat23aYM2NaqTGvbt66XQdNaMbkCaXGcyPyAVSpVr1GzTp161MO6kB9s+kXAhCAAAQgAIEDQQDB4kBQpU8IQAACEIAABCAAAQiUYwJhvhXyq1ApqLoWbSy0CCzhQtkWbUPR0PZNLJRtkWKh8lFsxUDAEie23HPj5ed5vTk5F1xx/S25dalSQWpXDLfLs4s2Hbp0i46OiZk3e/rUA3mf4uy7RXrbDrt27tyxcN7smcXZ78Hsa49/RSnyDTmYfLgXBCAAAQhAAAIlkwCCRcl8LowKAhCAAAQgAAEIQAACpZ2AfmvEW9S3kEjRyqKmhUSJqoFAQNkVyrjoETpXL3Se0lDF+OTXrFqx/OcR3351RJ/jT3LbFt51m45duktIyOt2SRWS9ayKvLXv0uNwdbJgzuwZRe6smDoQi6joaAlquW4yCZ81bdIEv22FvaX6i7N0ksK2L2o73c8TFRWVVz9tOnTupnMzJhfd6Dy/70lR58H1EIAABCAAAQhAIJwAggXfBwhAAAIQgAAEIAABCECg2AiEsiu0ECzfiloWEiZktC2xopIrEFDGRYqtF1e3zy3ss8pDKeNCJtzNLFQaCgPusCfSpecRR93R/8nn83pIx59y5nmPvfTOx3mdn2Kln7SQXqlK1WpOm5Zt2nX88Ouf/jz7kiuvz+26+g0bNx09ddG6w47qe4LOa2H84mtuvkPXvPflyN979z3x5Nyu69n7mOOeffOjIZ+NHDPl9UFf/6CFf/lXqO2COTOnF9sXLdRRbFx8/FX/vuuBr36ZOGfMnNXbB5uJ+M13P/REwybNW+Z2r4qVKld58OmX3/5j9qptY+eu3nHlTXfeF9kuMSmpQr20Rk1mhDITWrXt0Pnp1wcOfnvwdz//66zzL8lrDg889dJbauOcl5G5rhOL/s+88k5uApDGI48RcXXGLl+R/Dg1a9Wm3ZuffjPq7wXrM/+0OZx76dU35tZe/hWrVyxfunHDurXOeQlX/Z999d0b/vPAo8kpFSvldx8988tuuO3uHybMXTlu4frMAe8M+iq3sZ1zydU3XHb9rXeF99W0Zeu2T7zy3qDbH3xigEzgi/u50x8EIAABCEAAAmWXAIJF2X22zAwCEIAABCAAAQhAAAKHgoDEBmVW1LBQqSeJEfKokLF2ooUECy1g6s1++VeoVFTtUMjoWCWikvCy+P9Hd+Sx/U654Mrrb2nQqIkEnX9s/zrz/ItPOPWs8/PKGHBKPoUvmK9bs2aVOqrXoFHj3Pps2iK9TWxsXJxlwgTkQfH6J0N/uPX+R5+pbL4IVi2p81kXXXFt+HW6t4SAVz/+akT11Fq1F8ydPUMliV5473/ftOvUtYeMwBcvnDenOL+QlatWq/7xt6PHXfXvO++fNG7Mby8+/uBdGzesX6tFdi3qR96rRs3adT769udxx59y1nnDvhj04Vzz1Ljujvv+W6tuPZUj27PpWmVgSLDo0+/UMwd+PWpsj97HHKuMhf8OeOODXscc1y+3eUjYcI5L0Bk0/LeJEgiSklNSTjnnossbNd1bRBGfL3+eMPuqm/9zv8QBr9fn1dhvvOvBx/Li1PPIPsd/ZHOu37BJ00/ee/3FVcuXLfn3vY88ZdpD5chr1P/0yeODHhx6Po++8NaHL74/+NtTzr7wMgk1z739yZd53UcZFQPs/E139X988t9//vHjd199ftRxJ5167MmnnxN+jdrdct8jT19+4+33OMdbt+/U9YOvfhwjIe3Cq264VeeL87nTFwQgAAEIQAACZZsAgkXZfr7MDgIQgAAEIAABCEAAAgeNQEhkkBAhQUJv8yvDIsciyyLZMioSXFaJxz5L1HDbZ71JLjEjzUIlozpZyIxbC/MSPdiMwJyZU4Nm1c3T27aPBKIMg47dDjtCC+zVqqcqi+UfW4UKKcHSTrt27tjunPTmZGfr88L5c2bldo36zLE2Uyf8NebJV9//tHP3w3s/+/Ddt558eLsmR7ZNq3b71ReeEX7dI8+/OfDUcy++4uE7b7zyklP79Lzv5isvvPHiM05MrVWnroSSYHkln89XXA9UC+WvfvTl8Fp16ze48qwTj3zkrpuvHvzh26/ZeMdKZJGAEX4vtdcCfZVqNVIvP+O4Xk/cd/sNusZjW8vW7SWU7dmamkN4kNeO7dsfe/Gtj2RgfmznZnWuOPOE3jp+3uXX3Rw5j4qVq1RVRsX4Mb+OVqmtZ9/6aMjCuXNmnn5Ul1Yn9WzT6JgOjVOnhxl416xdt57EnYD9R6F+LzzpyK7nn9ir02+jRgw7/fxLr8pNfGrUtEWr59765Iu5M6dPOatv97YD/nvv7Y/de+t1EpTOv+K6f4ePSeKWxuSYhvd/+pV3Tjjt7AteeOyB/3Rvmpr40/BvvlTmTl6ZKBIZJLqI0V3XX3rOPTdcft7WzZs2prftuEeU0f2atGjVWvefNG7s7/pbz/oZy7BZt3rlilsuP+fktbaX4FZcz51+IAABCEAAAhAo+wQQLMr+M2aGEIAABCAAAQhAAAIQOFgEJECozIxMtuVJoQwKCRT63ZESFCjCfRS0yu52K/MizUKChYQK7fV3AlkWux/b/Nkzp2mf2+Jyt8N7H6MFY503vUKZKv/YtHidlZmRsWXTxg3OyZZt2ksccs2cMnF8btd063Vkn6lWSuqkM86/+Ig+J/zrvn9fddEn77z2gsQAZUuoP+c6CRXK8PjgteefGvq/D991jk+b+PefSxbszqqYMv6vMbndZ3+PKavCyk11vPOai87SfZx+uvc6uu/s6VMmrl+7OphB4mwXX3vzHXrz/+E7b7hizozdApDDzefzesPbNm7eIn3j+rVrrrrlrgckDvzn2kvO1pxnTZs8waa9q3bd+mmR49biv8SPyeP//EMCz7xZM6ZedfYJR65asWyJ2m621A/nGmVTPPbyO58og+Xac0/uEy6uTPjz919szb9inXoNlGm0Z9M1j9s1EpFuveK8U3dY2oxO6to3Bjzx0I/Dhn4e3l6iif6eNnn8XxJAVMrqiftvv2HgGy8+k52VmTl90vi/dD4yu0TH2nXu1lMCiASgrz4d+I6OOZk2lgSyFys9A53/eeSwodrfeFf/x2z4FW+65Mx+v/44/Ntxf/wySkJapH9KJD/+hgAEIAABCEAAAg6BPE3GQAQBCEAAAhCAAAQgAAEIQGAfCajck4QKlXmSaCEDYgkSVSwqmFjhsZXPPV0G5Ge82we6eqjNNturlJRCfSkjYK8F0n0cT5lovnTR/HmaiFUBkufHXtsxJ56yJ9NBpZhym7AWr5csnD833EC6Tceu3SU6OGJI+HXyulC2gBasb7q7/+MfvP7C0yO+HvJpbn2rFNEt9/73qQ3r1qx+68WnHolssz1sYb24HoYyTa648Y57v/jk/bf++v3nH51+NRaVbfro7VcGhN9LPhGX33D7PWN+/nH4j8O+2rOw39z8NdTOGOzlrSFhKMWuaZHersOZx3RtLZFA7bRov3Pn9u2OWBB+j06WgSIxo2fvPseZBUby5acf12vnjv/PaAlvKwGhY9eevR6/97brF8ydtZcRuZMFozGHX3PG+ZddrXk/3f8//5aY4pzTM33z+ScejmQrDl5vTs6mDevXvfbx0JHffj5o4JCP3n3Daed4UeQ2l1vufeRpCSwqseW0T2vSrIV8UObPnhEUz5zNklGCDMVWGSBnX3zl9U/cd9v1ptMs0vGgWXeE2XtxfQ/oBwIQgAAEIACBskmADIuy+VyZFQQgAAEIQAACEIAABA4qAcuGkDCh8k6tLdItJDqYIhEs7aQyURm24rvDQqKE3g7P8XiUfBHcllnMtlhtIQVDmRm6Ppg5UN43vd2vRer6DZvu5WGhReejj//XaSuWLl4oRjXr1K0fyUrig7wVrGTPXiWS5Csx0zIGtKgdeY0yEXRMmRUb169b+8Zzj/fP6xmcc+k1N6r0kN7y14J9ZLsaNWvVsZfyvVOstFRxPcdrb7vnoW1bt2x+4bH77wzvs1uvo/ooE0GeC+HHz7jw8muSKlRIfu3ZRx90jmvx/eKrb7pdGQpOFoRzTl4TYvv2S08/GnnOukmxW2+KnIsEgh3bt27Vgv3zj95/p0oh5TZfje+Sa/995+L5c2d/Mej9tyLbmD+1hDpXVlZWpnNOY7niptvvXb5k0YLBH77zWmE4tunQtbuyQ2SuvX3bli1PPXjnXmWs6jRIk7eMa9nihfPD+2tr3wuZpCsTY9fOnTucc/LZsIpi234Z+d3X4e2bt2rbXmKYMlr0XHTPLwd98LbTRt/JbcZLYk9hxk0bCEAAAhCAAAQggGDBdwACEIAABCAAAQhAAAIQKBIBEyv0u0LZFMqUkIFxHYuKFlqklGihTIkVJlbsCrjdOhZcvAx78VqChd5y18K7Mirkf6EMjYqhvos0vrJw8fIlixfWb9hIJuZ7tsOPPvZEK79T6dVnHnlAB+XnEDnXvv1OO0uliv4YPfJ755zK8yjrQiWfcmPjGFbLZ+Hlpx6+Nzs7Sx4k/9jks3DupVffqIXsYV/876PIBhJL5GExe8bUSeGL30V5HirHJCFlyMfvvhGZwSAeWhiPFEdOPuuCS1UCSSWddG+VgnrWfBaqWqmiJ++/48bw8agcUzVTWSRK/O/9N14OP6frJHSsXLY4mD3gbOJrSRmtdd0icxv/5vNPPshrjn0sI8am0OjDt15+LjdPj+q1auu/HZf8Ipw+JEqJ4+eWISHxpyB+GqMlyLS1xJDsY086/exnHrr7Fj2j8OuatWzdViJDeJkwnRcrlYxySkHp2DW33tP/RPO/eKb/Xbc4Bu46ru+RvivTJv39pzIwZFA+4JF7bw/P5Ekz9UdCS0Fj5jwEIAABCEAAAhDY828rUEAAAhCAAAQgAAEIQAACENhfAiGfCZWa1ZvhEim0V7aFQtkVWuyWn8AcW+FUaR0ZQKtdjBkOO7fVm9xrLVTqRgclfKRZSLhQP+V+W7l86WIZGleuWk1sglu/08+5cMaUiX//8sN3X2uhvrYZH0SCOu28S67cuGHd2r/MS8A516Bx0+Yqn5SXYNG0RbpKern05vxP33/9RV7w23Xq1rNKteo1fvxu6JBwTwunfYcuPQ7X54l//fFrcT3Acy69+gZ5Tnw2cO9MAy2eH3Zkn+OXLlowL3yxXx4N8vD47svPPtYYuh7W++jPRo6d0qVnr6Nuv+r80+fP2bscVJqxUbsfvv3iM2W2hI+7QaPdGS7zQp4izrl6aY2aSCTQ3++98twT+WUT9Dv93IsktHz/1eBPcmMi9irTtG7NqpXO+ZPPNhHBRKNvhwwaWBiOLdu06ygxqa2JUjIBj3yGElgaN2uRLp+NyP569D7mWBl/S5jQvGRsrsyJ15559IGvB3/8fnj7ug0aNk60+lczp0waf9FVN96m8lzy4HDaKPNG3w+JOIUZN20gAAEIQAACEICACJBhwfcAAhCAAAQgAAEIQAACECgKAYkVyRZ6M7ymhco4OQKGPBX0m0OChMoFeaymfdC0Qn+bh0VWqCyU6vXremVVSKRQSShdq32iiSLl3ntvxdJFwbJPWkTWXoJDrz7Hn6RFZJViWrtq5fI69uZ++INUaR8tXg+2xf3wt/nbdthtyDx1Yu4ZFo0tW0DnP/vgzVfyW3zv2fuY49Tux2+/HBx+X+dz9yOO6qvPkSWacmtb2GPHnXzGub//NPK7cB8HXSvzZ2VMRM6pY7fDjtD5DEvxePeLEb+9+b9vf5K4ckG/I7uE+18491emgD6P++PXnyLH5BiVz5s1fa+F/ibNWwV5SRgy8WYv8+vwPlTaqbuZmf8xesR3ymKI7D82Lj6+Y9cevSwTZKLDXSJVVzNWHz/mt9GR2RB5MWvTvnO34DkTcZ59+J5bI9vVb9i4qQSWyHkoo0YZLBJ9Hnn+zYFDf5k4R+XEbrvy/NNUHiuyH2Vp6JjKX510xrkXvR5WckvH5YOifeR9CvusaQcBCEAAAhCAQPkkgGBRPp87s4YABCAAAQhAAAIQgECRCCizwkLig8QKeSdo0bapRZKFsiqUGdHYQtkUKgslwSI7EPDLM0EeALNtUXaO3+9TqZrKFg0t5IHhZGpIwFC/8rKID92rSGMuzRc7JsaOYHH8KWedp/mM/HrI/7RfNH/OrHppjfcqGSVjapVikvAQPvd2nbv1VPZEbgvgMkluaIv2MpoePvTzQfkxUzkgCSG5CR96i98xBM9LGNnX56HsA5VGUkZJ5LUnnHb2+ToWmTXSvnP3w3T84QGvv1+jZu06/W+77rJzT+jVcaGlSeR2fy3m67g8JiLPd+l5xFHKdJBPQ/i5JqGMlO8tiyO/kk3N09u0lyjxt4kPud27c4/Dj9T5338aMcw537Fbz156JuN+/3lPhkxB3Fqbn4bafGdluiIzSHTcKfllft97CS/tQqyuuOmOe488rt8p777y7OMnHda28c8jhw3N7Z7NWrVup+MSxsyi5NfpkyeMC2/3/4LFPzM5CpoD5yEAAQhAAAIQKL8Eyv2bSuX30TNzCEAAAhCAAAQgAAEIFJmAzLRVonBV9yIAACAASURBVEhvpeutfWVFSJiQqbayJlRCR/4VKq0jYWKLLXBL0Fhq8Yu9AK7yT3oDvlaoH8fMWFkaEitUnkelorZYSAT5h0F0kWdQSjpwjLXrWRkeDflfZ51/iQyQHU+BhSZY9LSSSMoyUPaBjLPl6fCReSVEmkTLWDkvE+xGzVq00gL5H6N/+D43c+lwXBI2tOgd6SWhNr37nnhy1Wo1UmVaXdjMgIIehcatNhP/3LvElIysjznh5NN1Tl4V4f1I4ND9H73739do4T3cXyG3+9Wu2yBNxzesWyMD+D2b7qGMEgkikeWvJESo4chvvvgsvzk42RtzZkydnFu70869+AplVvw0/JsvnfPp7Tp20ecJf/1/qaWCOJlg0VVC0lsvPvVIbm2bmr+Fjs+ZMWXS3qxqK8PJNeCR++744pP33izId0RCjdgqu+Ku6y49J/JejZu3SNd88ppvQfPgPAQgAAEIQAAC5ZMAGRbl87kzawhAAAIQgAAEIAABCBSVgLIrlEUh0SHDQpkRypSQ2KC9QtkVyrxQaRj97bf1SwkYEiYkQmi/zmKDGXKrD71QVcXaSMBQtkUlC3leqEyU/DDK7bZs8cL5mnz9hk2aauFbgkS4ufOiubszBhwPhlvue+RpGS0PfP3FZ8KhyVS6UdMWraaO/2tMbjBbpLftoOOjR3z7VUGwZaodaUDtXHPxNTffoc/FWQ5IC+QSRySChI9NYoWECJ1Tpkn4uUrmo6DsFIkABYkVus6aV9Niv1k4bA7vp9fRx/XTfEeHiQnO+Rbp7TqoLNLMqZPG58esuply67xVjtpLDNExiTvKahjz84/DV69YLkEvuOl5a79y2dLFBT0PnZdnhMo6qdyVI3JFXte0Reu2EiOc75RzXqz0efCH77xWkFihdsp4EZNVy5ctmfT32N8j76MMi5XGXp4chRk7bSAAAQhAAAIQgIAIkGHB9wACEIAABCAAAQhAAAIQ2CcCIaPtKLtIgoWyLLQ5QkWsfdY5K+XkjnK7XbVMgFC9fgkVAcuq0ELwBgtlYuj3iFfHrd6+rgv2YW2s34D14VY2ho4pW0OZFuqj1G6TlyvJJOjpIWb1djMKGo0vsfB3qCdtJvdt04b167SILkHi5DPPv2T92tWr/vxt9A9Oa6f0j/wUzN6iSqfuh/d+5qG7bpGvQniPbaxckMo1TcnDv8K8IIKCxdhfRo0oCHRiYlIFG5bGv9fW96TTzlKZIB2cNXXyhIL6Kez5WmYqvs6EgfD28oW45ta7+69ZuXzZquVLl0SKEinGIpJBfvezikwJGeYJEtnmvMuuuUnloEZ+++VeWRTyEpGx91efDnynoHmob7WRn0Zk2yv//Z/7ldnyyTuvvhB+Tibrum+kgJLXvSRk6VxeZZx0Tt4TC8xsPNKfRKx0PsfuV9BczAIj0fFM+ejtVwbk1l6CRXGVAytoPJyHAAQgAAEIQKDsECDDouw8S2YCAQhAAAIQgAAEIACBg0VA2RVadJegoJJQDSyUBaGSUC0tWlnYYnzAa4uiGpPECLXVQvBKiyUWGy1U4kmZE/KrSAtdb+3cEjKcDA15ZCh7Qz4WEkJK1WYihdvCYyFxR6zESW/ay7NDJXhkVO6IPvnObdG8ObMaNW3eqp+V4Bn62UfvhRtpy5NBi/UqIXRH/yefl4Dx2cC3X43ssE3Hrt21+L3UPCxyu5nKG+nNe2UMFAQ621bStXAd3k4ZHHc+9OQLMgLX8UUL/ukFUVC/eZ1PqlAh2evN2ass2IVX33jbpHFjflPWyLRJf/+pa1W+yeljl6WZmE4QFAoKsykbID4kLDjt5V3RrddRfb79fNDAzRs3rA/vp3l622A5qPFjf/u5oP43rl8fFI+UBRHetqkJCGdfdMV1f4/5dXSkEbj9h+aWkBEVHb3Xy4Y65ohC4X05gsVfv43+Mbfx6PlIYFlgtbwiz4uVjjnCSn7zEW8JXyqdlZs4IqFFoe9sQVw4DwEIQAACEIAABMIJIFjwfYAABCAAAQhAAAIQgAAECk0gLLtCIkIjC9XYl3+FFuG1MKyQQLHDYqHFIguVwNGb+FrUHW4xzUKLtzo+3UJloXZnWthmGRa2TuvRbxUt7GqRX+ckkqjfErspgyIsJFTojXVHnOgY+qzyWCdZZFvMC/Eq1O8yvRUfZ4vv1cyn4stBH7wdDkICgcrvnHTmeRdrQfqpB+68KTcD6I5de/SaMWXi35Fv1zt9qezS7OmTJxYGskSS7r2O6hsbGycxxqVF9UdffOvD6qm1amvxXceU+VCYvgrTRp4aqbXr1nMEic49eh154ZU33Dr8q88HSQSQv4QyRL4bO33xuZYRoT6XLlowT0bazhh1TAvt/U4/58L+z776buR91V7zcPwmVPLowWdeeUflpt58/smHI9s7fhCzp08pkJnjGSF/D6efJFMQHn/5nU+ysrIyH7vnlmsj+1++ZNECjbdDlx6HO+ckVjz9xsDBb376zSidC7+mVduOndesWrHcMWmP7E/ZFTqWW7kozV3nHBNx51rd+5Hn3xxYs05d+coEt8bNW+p77Ppm8Ccf5PY9cwy3Tc+QQMkGAQhAAAIQgAAECk2gUP8wLnRvNIQABCAAAQhAAAIQgAAEyiyBkFjhZFeofpHq62sBVKbbyoTwW2ghXiVl5FGhxUqVf1INe2VUaFF3rIUWRiVYLLeQ8e9y87DQG/lB0SIQ1C2C2oUW/JV9IdFCn5NsDLp/Sd40Pnl39LS40+Iei4stOlsoE0VCjxipNJZ8KX6zkH9Hgdus0KL4Lz9+/82alSv+IQRsMLNtiT0/ff/1FxP/2tuY2um8SYtWrXMsNeKxl975+Nb7H93L30IL0ipxNMUW/gscjDUYNmTQhzVNQHjpg8HDzrjgsqu1gK7F+OFDPx80IZRxYGvrhcoeKcz9xo/5bbTG98CTL7557W33PPTSB58Pe/zeW6+rXb9BQwkw1cwj4t0hI35bvGDebI1BfY74+vNPlVXw4NMvvy3T7PMuv/bmIaPGzXj0xbc/yu2eznVqL9Fj4NBRY80SotGTD9x+o8pwRV7TrFWbdls3b9roLPbnN4/pkyeMU2bDdbff9/C5l15941HHnXTqe1+M+K1h42Yt7rnx8vMjPSXU1zdDBg3U/uEBr79/4mlnXyC+b3727U+6duAbLz4TWQKrZZv2nczkei8z7fAxOWJEbmWpRtn3Jse+HHc/8uzLvY45rp8yeV4f9PUP73058vdmrVq32x7m69GwSfOWyvD54pP338ptzo5gUVyG64X5ftAGAhCAAAQgAIGyQQAPi7LxHJkFBCAAAQhAAAIQgAAEDhYBLUCrDJAW5bUArwwCZT5oEd6pza8XoyQ+aO8IGRqfFuYlZGiTIiEhQ9c55aHUb/hLVSoXpbe6nbfLJWroevVdIraQL4XGEjQMt2hjoXlIsGgemp/ECYk32iujRIKOfD1c+flWRE5Qi916m/2D155/KrfJ79i2batKFj3733tuywuOvXy/tHffE/6lBfb/XHfJ2eHtZKKs/n/54buvCwP3y0ED3z725DPOUbkkhUSDrwd//P4T991+g63BB9/Ab9CwSTNlPhSmv4LaKKvksKP6nnDquRdfoXE+89Ddt8hMWyWwdO19Tzz/+uvPPd7//VcHPOlkkPw2asSwX03g0eK7Qu1kjn3HNRedKWEn8p622D/584/eef2si668TpkFylx5zESRYUM+/TC38YmZFvrzyliJvOa/d9545csffvH9XSYK6JwMtq+74NRj8yopNX3S+L8+fPOlZ2ViLpFJ12hMLz3R/+73I74H8i5RpsnG9Xv7loSPweNxB//72rxpk4TEvTYJLy8/+fC9tz3w2LMSg3RS2RovPPbAfz59742X5KXhXBBndaM+fOvl5yIN0J3z1VJTgwbjs2dMyVM8Keh5cx4CEIAABCAAgfJJoKS/nVQ+nwqzhgAEIAABCEAAAhCAQAkkEPKQUJkmGUa3tjjFQn4Vjjm280KUPAS0IC9BQiWi5lgMtVBd/cUWjiihbIM0iwstjrWQAOIxJSPgdgWsjVt+ASoXpcXVXyxGWUy4/8IuEjlKxCZ/ChuIhBX5UWgezSy0SCuxYlNo7H/bfrKFXLeVhbJn2xfBQhephJBZDQTduyM3lWLy2Uq+DLrzgqM29dIaNZky/s8/It/Or22pBCr18/tPI78rLFyVJGrbqWsPs31IXDR/7qx1a1btKQF0wZXX3/L9V4M/ifR9KGzfubVTBkmaqSGZmbt2abFfb/K/YgKAVaWKv/3qC06fMv6vMbldp8yDajVSay4x7w6VWSpoDCotZYv/qbOmTZ6QX5aAsh7+GP3D94U1xd79DCskt+vUraeEh2kmSET6cuQ2NgkjzcxfRKKUPDvMasMR/vZq3qZjl+4LTdgyX2+VZPvHpnJXLVu36yjRJi+RpW6Dho3NK6WlyjnNmz1jWrhXSkHcnPOxJmhY8k0D8S7sNbSDAAQgAAEIQAACIoBgwfcAAhCAAAQgAAEIQAACECiQQKgUk4QJCRTKIpAnQy8LZUAo60JZFvp9oQV5p6aTDJIlWvxq8YnFBAstpjumyMpIUDmpvhZHWEgESbSiUFFmZCHxQybAWpxXjLMYYTHSBItcF+wLnEQxNAjLqFBvGqM8PGSgLYFCXg4y0ZZ3h7JAVO5pdmj8PhMngnWu2IqHwMlnXXDpPY8NeFXG38qKePze264vnp7pBQIQgAAEIAABCEDgUBHAw+JQkee+EIAABCAAAQhAAAIQKF0EJEpIYJBvhQQLLdDLx0LHlWEgEUKChRbq9fa3siLkUzHFQkKF/BokQGjzhUIloiQ+LLFQFoYW+lVWyhE0lIFRyUJZGmkWEjeqmnhySErbhokV+h0lgUbmyU9aXG1xjIUyT5RJoQwFlRCSyKIyUHsMxUPzZ1cEAjIel6dDfzPD/uitl55TV7OmFWx6XYRbcikEIAABCEAAAhCAwEEicEj+oX+Q5sZtIAABCEAAAhCAAAQgAIHiI6DsAQkIEg+qWxZEQ5MnKptGIcEi+CKUlZjJtoo9KkUjIUKChcy1f7eQ2XbQe8KyI/aMyIQHx3xa5tupFlrwr2XZFRIpJH445ZaqWd8Job6n2vEcu3at9aUMjoO5aUxioCwTfe5joTJWP1tImJllMcNCpawkygT2teTTwZxMabxXg0ZNmj3z5kdDqpvBtrwfNIer/n3XAyrdVBrnw5ghAAEIQAACEIAABPYmQIYF3wgIQAACEIAABCAAAQhAIF8CoYwGmWfLv0KRaqKCCQxulYhysiHskNspBaWyUGsstIgs/wZlTsiwN7Ikkhb1lWGhthItVlk4RtzOmNR/BbNKkIlvS4v2FhI2Eg5GpoWyKkKhcTS2uNjiGotzQn9rXsqikG/FXxarLcioyPcbtX8nj+hz/EmffPfreG+ON+f8fkd0/nvMr6Obp7ftkGVmEAvnzZ65f71yFQQgAAEIQAACEIBASSJAhkVJehqMBQIQgAAEIAABCEAAAiWMQMi7QiWfJFSoDJRSJGQsrUyLCE88t2VhBKracSfDYpF9VhaFXpTSwr4EivBNAoaOb7RYZiGD3jQLiRO6p/rXNX5TQ2IthcMyOoL3ViaDBI6AjW+XZVpE9lvcFCXMdLO40eK00Dglwmis71t8YLHOsin2MtQu7kGU5/76nnTaWU+8/O6gv37/+cc7rrnwTBlWi0e7zt16zps1Y6p5jUskYoMABCAAAQhAAAIQKOUEECxK+QNk+BCAAAQgAAEIQAACEDhQBEJiRaL1r7JH6RYyxVZ2Q4oJCB4TEHRrLdIrLAMheEALySqJpGwJeVioFJQEDJVvisyw0HU6Lt8KtZFAIQFDfydZd7HB+/y/MCKRRAbXtS2U8aF2EaJJ0WlEeFVIrOhvcbOFyl9pUxbIm6H5qByUymCxHSACTVu2bvvoi299NHXiuLG3XXn+adnZWfqOKKPH3aFLj8O//2qwDN3ZIAABCEAAAhCAAATKAAEEizLwEJkCBCAAAQhAAAIQgAAEDhAB/V6Qn4RKMXWykGhR3SLG5fcHdksFwTJQwcwC85nYaWvIEiqWWGgvsUIlnzIsC+If2QfyszBRRMeVhSHhQj1q8V+CQFVbkVa3jj+GbhBjx+raMWV6KHtDIocWr4vl7fowoUL3lSDSweJsixt0wLZpoTmNsv1vGqtlVRTLvUP9s8uFwF3/ffqlnOyc7HtuvOJ8R6xQsxat23aoUq16DQkZgIMABCAAAQhAAAIQKBsE8LAoG8+RWUAAAhCAAAQgAAEIQOBAEFBZJplht7GQd4SEi2oWMuB2NifDIdMOKKNCRtuLQ58lPuRWCip8rOFZFsrMUKkn7aNC2RW72+7O5lCGg8pFHW7R16KJRUUTPfb4aBQDBP1GkijylMWvFhIsnO1z+/CkxWsWQRPxYrgfXeRDoGaduvU7dT+89/ChgwetW7NqZXjTo4476VSVgvr7j19+AiIEIAABCEAAAhCAQNkggGBRNp4js4AABCAAAQhAAAIQgMCBIKByUBIsJBLIwyLFQiKGx8QEExr2mGzrd4XHsitibS9RQSbUMtJWdkW2Miny2kLnHPNtJytDpZ42m0ix3fYSQryWvSEfCxNH3OpfY2pkIRNsjS3ZRIvi+G2jjBJ5VTxgcV1ozBJgJLwMsfjU4kcLeW6wHQQC9Rs2aarbzJ89U9kte7ao6Ojof515wSUTx435bdvWLfq+sUEAAhCAAAQgAAEIlAECxfGP+jKAgSlAAAIQgAAEIAABCEAAArkQkDhRxaKihcSLcD8JpxSU9k445Z022DGFDLELNKK2NrpeooDeoNd1Kgm1wQQLCQOKLaZV5OwuERXMtNC4ZO6tTAgJKRVCY9vvh2jloCSEHGvxvcXVYR3NtM9nWNxhocyRPVkVVg5qv+/HhYUjkLFzR9AfJKViJRmu79nOueSqG5R98eWggW8XridaQQACEIAABCAAAQiUBgJ4WJSGp8QYIQABCEAAAhCAAAQgcGgISCHQQr4EAYkE4abZjkihkTkZEgvt83gL7fXWe4FiRdi0lEmhDAt5U6RZqNyTyknJ20JjaOh2ueMCu4egklQSURwhpUi/a0JihTw6vovArKyKx0Pj8ppAEWkafmieSjm66+zpUydtWLdm9UlnnnexykJZMsWmfqefe+Et9z3y9MJ5s2eO+n6onhEbBCAAAQhAAAIQgEAZIVCkf9iXEQZMAwIQgAAEIAABCEAAAhAII2DllSRUyBdCQkGw3JOFjmkvEcI5pmwDiRUSG1QCSmLDfAsJD3ozvtCChWVZ+Oy+KiG1zEJlmOpaRoVEEo1Db9f7VBFqt5WFS79jJFaoJNQSixUWG+36HaFsjbDZ5P3RhAr1XceinsWAiJbD7O87LeSpUeh5FOrGNCo0Aa83J+fBW6+9dMA7n341bOx0fb+Cm4SL+26+6kJ5WBS6MxpCAAIQgAAEIAABCJR4AggWJf4RMUAIQAACEIAABCAAAQgcdAISJJTF4JRqyjEPid0WEv9f/skpLyvBQpkQ8ptQOScJF8quyNwX8SA0Qy0+y3BbC9MSEiRUVLeoZfeP0Rhsk3jgt88Jtm9gY5KfRZKFSlZJOFFGRoFbSKxoZQ3lV9EzdD/nupvsg97cX0tWRYEoD3iDP38b/cNZfbu3Pf28S66sVbd+g+VLFi4Y/OG7ryvz4oDfnBtAAAIQgAAEIAABCBxUAggWBxU3N4MABCAAAQhAAAIQgECpICAxQtkVEiGWWEiQkFohsUBZCc7mZF5ISXAMuXfZ5wyL/X3zXfeS4KHFaPUrQUIZEMny3bZNgoT6z7aQqKIxSuQIjtmyLLwFCSUmVqjEVVuLVy3ah81HH0+yGGWhcbCVEAIrli5e+NKTD91TQobDMCAAAQhAAAIQgAAEDhABTLcPEFi6hQAEIAABCEAAAhCAQCknIMFBCoEyGWpFx8RqkV8ihgkWbo9lNjglotRO5Z9klK29hASJBvs8/dA1ul4ixBYL3UNCSCWPx+O8bCXBJM5uX8Ht8Sj7ooVFU4tYCwkcwTSQvDYTK9TfdRZjLMLFij/s744WIy0QK/b56XEBBCAAAQhAAAIQgAAEik6ADIuiM6QHCEAAAhCAAAQgAAEIlDUCWvTXb4XaFspEaBgVFZPk8warLZkoEPBadSYJFRIXJCyss1hqoXJQKstUFHNqRwBRn/VDYD3WoeMjIcEi2u22d688bpff6+1s4oXaymtCmRm5ig0mVOhlLXli9LN4OuyBabyXWvwV6gO/irL2bWY+EIAABCAAAQhAAAKlhgCCRal5VAwUAhCAAAQgAAEIQAACB55AyHBbpZYaWPSxONmiks8nsUI6RkAixSYLiQRa3JdgIaPsBRYSLZRpsb/loDRBiR3qc07ohjVs38HctuVnoQEoyyPaPCzcLl9QW0izkAfF7NB1O/OgVM2Op1sMijh/s/09wmK7+VUgVuQBj8MQgAAEIAABCEAAAhA4GAQoCXUwKHMPCEAAAhCAAAQgAAEIlAICIbHCya6oYkNuasJAS4ssn9drPhGBdSYcbLTjEiyUzSBhwfGsUIbDytDfMuLery1UFkrqyLbQPVbZfraNQX2r5JTEkF3mZ2ER8EdFx0hcUSaIsjEqWUTZPMJ9NlyWXSGR4zyL0WGD0rj/Y/GdCRVbESv263FxEQQgAAEIQAACEIAABIqVAIJFseKkMwhAAAIQgAAEIAABCJRqAsrAlhdEkoUyG2pauaWKFlmmDchXYrvL7VYJJcd8W0KAQr8rNljI/NrxvthvECHRQqKHyjupz3k2BvWvY8rA8Nrf2RaB3VYaQZ+NOqExJ9s+zkQLjwkVbgv5W1xr8ULEgM6wv9+ykLk3GwQgAAEIQAACEIAABCBQAghQEqoEPASGAAEIQAACEIAABCAAgUNNIJRdoYV/mWvXtWhj0cAEihjLqlA5JYkFjtG2shMkDOiYUxpKgobKMTntiuJjIRzqR5kcEiwyQuOqavug6XaIl8fvDyZzaNytQmOWj4ZECAknFS2etzg+jK+OP2jxq0WmZVYUdZxhXfMRAhCAAAQgAAEIQAACECgKAQSLotDjWghAAAIQgAAEIAABCJQdAsqUUBkoiQISLJSZUN0EC8thcNvvhoBCi/vysFDJJmVZaPFfYoLECh13siuKQwRQHyoLJQFCZaEkXKjsU4qFkyluiR/BW0nAqGfRxGKxjdiTWlVJIq7GFjLZdraF9uEhiy9NqNC42SAAAQhAAAIQgAAEIACBEkQAwaIEPQyGAgEIQAACEIAABCAAgUNIQIKFPCBqmDeEPCFq28J/csDvl0xhqkDApzJM9ofKQklIkJ+ERAqnFJRKRUk98IdKOhVpKqE+si3zI1gSykLiQ6pFcwu3jTFYDsp2Npxg1kWKfa7l8bjrm1iR1KB2pTQ7dlbYIP6yz5dYLDKxoiim4EWaFxdDAAIQgAAEIAABCEAAAnkTQLDg2wEBCEAAAhCAAAQgAIFyTiBkUq3fBsqckHBR2UIpCvqsTUKEykBJqJCvhEo/6bPqMUmwWGIhM26dU+ZFcW66zzQLiRXKopBwobFKdHAMwp0xxiQlxFZp0ajGyUkJMb3CBqHyT2eYUKExskEAAhCAAAQgAAEIQAACJZQAgkUJfTAMCwIQgAAEIAABCEAAAgeRgEosyWxbvhRtPVHRx1hmhZlYB2IslWH3MNweOx9ICpluq5ySI16ssM8qtbTVsiKChhL7spkptporQyIomJioECl4SETZYjHXQsJFukVdj8cTtTvJQuMLGm/HJsTHNateJam6iRUdwsbwin3ub/3KD4MNAhCAAAQgAAEIQAACECjBBJzaryV4iAwNAhCAAAQgAAEIQAACEDhQBCy7Qr8JZFot/4paFl1jYuN6mSBQwz5Hq96ShceUgXj7W4KGxIrNFlst5C8hwUIeE8rA2N/NxBFXNwtlT+S2SZXQPaZbTN19f7dEDgsN0OQUjzsutVpKWsM6ldt5vX5lgLiyc3yvWXxqH+WxwQYBCEAAAhCAAAQgAAEIlHACCBYl/AExPAhAAAIQgAAEIAABCBwoAiGxItH6l2dFS4tGFil+ny/oDaEIbkGvCL9KMMlPQlkOynZQeaWVFk7mQjDNYT82CQ8SKiSQpEVeH8raUJaFRIglFqMs5tt49mRzmFjhio7yuBrUSnYlxMd4oqM9SbsycxYvXrl5yrhpy5d+96uGywYBCEAAAhCAAAQgAAEIlHQClIQq6U+I8UEAAhCAAAQgAAEIQODAEdDvgRSLmhbVLVSOabPPm7PdBIFEj9vKLgUttwO7TLzYZlkWjkAh8UAChQQMZVvIfHt/vSv0EpWUEZl4B+tD5bJJLJGpt87LM2OdjWezjSfFxIqYqpUSPelNarjMv2LPpfMWbxi/duOOLK/PX9EOKsNCogcbBCAAAQhAAAIQgAAEIFCCCZBhUYIfDkODAAQgAAEIQAACEIDAASbgCBYy2ZZwEW9CQJbf79tie5/LMhdsk2CRaeJAUCiw0G8IhUpASayQv0TG/vhXhOamMUgskaG2Sk79Ywv1LVHEEUY22njWWmTXrpHi7tqm7t5ixZINi1dv2J5tYoX6rap5WTbJ/maAHOBHQPcQgAAEIAABCEAAAhCAgEOADAu+CxCAAAQgAAEIQAACECiHBEIL+CrHpE2pCQ0sjrPQAr+EAacklNtKQumYvCtWW8jLQpkV8q9QWaiiZi9oDPLPqGSxKJ9HkRW63wLbp1k0ion2NKtXs+IeISIzyxuYPHt1xradmal+f0DG2xqbSlg5Iss+m4KXw68GU4YABCAAAQhAAAIQgMAhI0CGxSFDz40hAAEIQAACEIAABCBwSAnot4DjX1HPMirqWqRFR8dWtcyFZAtHzNAiv0pByfRaAoDKMimzQqKFBAuVhyqKEKBrZaY9w2Lp5OXbXIrIzbIsnn+cAQAAIABJREFUVDZKZaGU0bEwPi56tbIrqlSUX/jubc6i9f6tOzJj/QFPos1Fvhzy5JAQI8Hl/+tFHVLs3BwCEIAABCAAAQhAAAIQyIsAggXfDQhAAAIQgAAEIAABCJRPAhIkJFioFFNTEyjqWXjNu0I0KlhEmYeFPktQmGkhQUEihUpDyWjbKQel0lAhd+79Aqmb6KYSPlSWKr9N9/HGx0ZvaFinckKztGqOqOJau2GHa/O2jCifzx9tHhyWFOJ25ibRQqWhYkIm4/s1SC6CAAQgAAEIQKD8EUhITExKrVWnbkxMLC8+lL/Hz4wPEQEEi0MEnttCAAIQgAAEIAABCEDgUBEIlYPS4r/KLCmdoWpUdEwr28ebf0Vuw1JmgwQFiRMSCdRoa+hYUc2sZaitsk4qNZUW6j9PNFEeT6BCUmxMcoW4ZCsJFfw94zdf8LlLNrgystTV7s3mE2M7lZpS3ypxpXHiY3GovnTcFwIQgAAEIFCKCNStn9bo3SHDfx07d82OEX/PXv7XgnUZ73/5wx/9zjj3Inspgn9PlKJnyVBLHwE8LErfM2PEEIAABCAAAQhAAAIQKCoB/dB2Xl7yWfmkuKio6ES/z+vy+/3KTgj275Ye4PfpN4OyFXRQ4obKQCmKarbtzEEqg8y2JZ4khe6T1/x8VgLKWzs1Ja165ST5bQS3pau2unZl5jieG8Hx29g9Ni+9DRkTKm8loUVzzrd8VagcldoGs0Y61EsJppywQQACEIAABCBQfggMePfTockpFSu9+/Kzj2dlZmbUrt+gYe8+J/zr0Rfe+vCsC6+49o5rLjpzw7o18vZigwAEipkAgkUxA6U7CEAAAhCAAAQgAAEIlAICWpBX2adUizq2oJ/ktTJKtsDviBXBxXq/1VeynYQELfQrS0FG28ssVlgowyJozl3ETfdS/ypNJWPvOAuvhAMTC/bqul/v5v6sbG8Dy7K4zDnh9fr9q9bvsLH63aHxB9WWwG7hRf3W0Bwtllust+wSb8gPI9iF3ccRbxyRQvvDLPpYjLTzv9k+KFpEjqeI8+ZyCEAAAhCAAARKIIHW7Tt1bdoivc1/rrvk7B+HffW5M8So6Ojoi6+5+Y7rbr/34Y+H/fz3FWccf8TK5UsXl8ApMCQIlGoCCBal+vExeAhAAAIQgAAEIAABCOwbAVuw14K8yi+1tDjW4hRPVHSasivCNokIu8zPQn4V+iE+wWKqxUIL+VgEsyssiiv7oJL1VdmipoWyLVR+KrctOS42up+d6GWR4/X5t8xetG7Btu0ZaTZgCTDKBAn6Wvi8wflUMM3iBJuHMjckhIxOTorLGTV9jb9qpUSJGcrAaGzR2UIXdLE4wqJN6OZ32/5Ei+F5jIfDEIAABCAAAQiUMQL1GzZuun7t6lVjfxk1Mnxq9m8L7/uvDnhyxuQJ455/939fv/HpNz9e0K93l21bt8jXiw0CECgmAtRcKyaQdAMBCEAAAhCAAAQgAIHSQMAEiwQbp7wdjrQ4w+KkmLj4mOxM6Q9W92l3OahgZoVlLMyxv8fYZwkWcyyUpbDdQp4WOZapUOQpWwaDhIOjdWsLiRW/W0gU2SujwdpJiFBmxdvOTddt3PHM5NmrPaZc9LZxNg1dHyx1pWwLjyfKZSaZrpycrFlxsVEjrYzUj/VqVdxkokVcdJSniTWTOHF66Lq85jLeTnQXEzIsivy46QACEIAABCBQKghEmxeWZZ/m6dPVs/cxx7384Rff/zZq+Le3XnHeqaViUgwSAqWEAKbbpeRBMUwIQAACEIAABCAAAQgUlUAou0KZBhIGqtmiviJHv8eDvg8WWui3TeJBgv2tkk8rLVQKSr4VEitUIkpllYo6HOd63VBvJipr4lyLtDw6Vn2oi8PPLVy+6SfLslht41yrMasEVFCosHnERO+u8BRvORRVKyVUadW4Rp/0pqnvV05J+MvEil/t5LsWl4RY5DeXH4trovQDAQhAAAIQgEDpIJCfWKEZjP31p5HvvfrcE0ce2++UPv1OPbN0zIpRQqB0EECwKB3PiVFCAAIQgAAEIAABCECgOAioJKxC6RQqodTAItYMHyL7loggc2q9WejUitLfwcwKi6CqUUyb+lKJKY1L2R/VLYJpHiEDbO2lPqRbSNQIbiZUDPD5AhqLM06ZhwckukRFeYLii8fjdlkJKZdlVFSOjvZUi/K45dlR2E2MbrJ41qK4Sl8V9t60gwAEIAABCECghBN4+8VnHl21YtmSW+9/9Bn5W5Tw4TI8CJQaAggWpeZRMVAIQAACEIAABCAAAQgUmYC8K6papFk09Hg81W1hPyqUVbGnjFLoLsqsWGKh7AUnuyJoWF2M2RXOhJbaB2U8DLXwx8d4YtrXTfZYuE2s0AJADwuVinK2mZlZ3nd3ZmSvtgMqH6UMkFU2j0y3x+PyW5aF30y3patk53itJJQ/dsfO7Gi/P5CXN4bTr4QTlZyqa1Hf4k0LHWODAAQgAAEIQAACexHIzsrM/OitlwfUrls/7diTTjsbPBCAQPEQQLAoHo70AgEIQAACEIAABCAAgdJAQIKFjK1lMt3SzLZV9sntCBZB/wqrCmXnlEkxw0JG24sslllskVhRnJNUQoR8IUyY8NmtZZjdSWFagwy4o9Zsy4qx47Xs83kR933NhIhFlmWxyo7LFHyexUwbv8QLv8/nD9j/c1kGhmvHzizX5h3Z7rUbd8St27RzfnaOb0kec5BA85bFAAuZjStybHwBjRH/iuJ88vQFAQhAAAIiULFyFb1EwFaKCXwz+OP3t5vr9tkXX3V9cU2jboOGjfPrK6VipcqK4rpfUfopaKxF6Ztryy8BBIvy++yZOQQgAAEIQAACEIBAOSJg/hUqs6TQb4A4EwuiZVexlwIhDwu/f5udn20x3WKhhRbud5hY4ZSGypdaeLaGBAn9HQp9DpZ6Ch3XOOQ5oQwKlXxSKagGNoTYhFhPVI4vELN5l1clq9qEbqihajzHWwxuVa9SdoPUZGVMrLCYZSFxZYaNXyKG3xw5XOZVYeWgYl2N6lRydWtbL6VmtQrtY2Oi0iImoOuU3XGzhcSK+Rby6WCDAAQgAAEIHDAC6e06dvll2pINvfueePIBu0kROlaJo/+N+GPyMSeeckYRuilRl8pv4vNRf+nfN4XaTjj1rPNvvvuhJ/JrvGvnzh0/Df/my3adu/VUpkWhOs6nUZsOnbt9+8fUBc1atWmXV7MnXnlv0EPPvfZeUe9V1OsLM9ai3oPryycBBIvy+dyZNQQgAAEIQAACEIBA+SMgsUBm2xIBOnqiolIDfl9QTAhmVtgWMt2WCKBSSzLYlo+DQl4RBW6OYXdImJAIodBvDu1jFHZOe4kUMv9WVkWS9pUSoiU6LDMFpVG2N1B19dasil5/oL2NrIGZaI+w/fVmSXF6tQqxv1hGxqaaKXGuC/s09ydnrd0R792+OcaXsS3Kn70+xuPfXDUlPlC5UoKrRaPqru7t67vq10qxue09fCsbNcqOXGlxisV/LL62LIq1Fj4no4KsigIfOQ0gAAEIQGA/CWixV5fmZGeVSJG8YeNmLZqnt21fuWo1vVBQJrZjTjj59GRLTSjsZG574LFnL7n233fGxsUrQzXP7afvv/5CGau9jjm+X2H7zqtdp+6H99a5Hdu2bs2tjZXz9LTv0uPwHdu25Xq+qPffl+sLGuu+9EVbCIQTwBCG7wMEIAABCEAAAhCAAATKOAHLrpBoIKFA3gxdLPpGRUWn2CLJbnfrPYKFzKr9KgelH8GO4KDMir0SMZwsighsTgaH9vqd4bwcpWv1OTa0198KCRYKnQuYAOHdmuHNskpO52Z5fRPs0DcmUCwzT4pF1SvELEyIicqsEBclg221V//+wLxfXWmetVEbvckx/oSUijGJyUlR8bHRzZrXjY6J0fD/ua3dsGPd4pWbXzYD7sHpTVLXHNasqjJK2CAAAQhAAAIHlUDTlq3b6oYzp04af1BvXMibte/a43A1XTx/rrIuy8Rm/6bwbNqwYV1hJlOpStVq1WrUVFlKV9Xq1VNXr1guv61ct/Fjf//Z6lH6uhx2xNGfDXzr1cL0n1eb1iZkbdqwfp3MvHNr07hZy/TEpKQK0ydPGFeU+xTHtQWNtTjuQR/lkwCCRfl87swaAhCAAAQgAAEIQKB8EZBYoDrZWhyRYJHgD8iUevfmZFnExMa7sjJ2KKNCZZGmWcgfYoeFhILIzclZkPjgfHaEEb2J6AgWune4OKF+dPMEC6kK+mz6gjvbRISdfl8gxZI+OltJqGHJ8dGzqyRGu22v3y0VQwPICVpUbN/gWxLbJKV+h2qNq6xZlpLQpMMFUXEJLf3enBxP9G6xYuf2nS6ZcG+zKW3YuMOV7fe4tm7f5fJl56RHeXelzlw2ed33T90RdeJdz+Y2v1ymzCEIQAACEIBA8RBQyZ+Vy5cu3rpl86bi6bF4e2nXsWsP+/dBYO7MaVOKt+dD15uyWewdjYicy9zHI8HCOWMveeS7fpqVmZGxeOG8Oc1CIlRRZti6faeu+YkR6XZe/c+YMv7QCxYFjLUoHLi2fBNAsCjfz5/ZQwACEIAABCAAAQiUcQKh7AqJA3UsmtraQ0P7pe6xNwH3lIKykksSLbze7Cz5QehNT8dsWybWGY7ZtlPyKYTMyahwBAv97ZR5UukpiQC7LJTZobJPKaG92ksEkZChLduioo3BnZocN27l1sylJlicYMf+qpwY/UV8TFR0Ro6/ohlsx9mFmeu3Z1fIzPGmBrzuWr6oCje4qqa0rVC1/p6n6LHcCuePrK0bXGvXbnJlZHld2Tl+V6bP7fL6PRVdHk8Tjy+rUaxv57qqOxf7F93eLrvO1qlOJomTTRLMBIl7J/8vSNaVexY+9mShFHRNGf/KMT0IQAACECiAgJVljGraolWbX38c/m1JhaW355cvWbRghzlKl9Qx7uu4sk2wSK5YqVAloWJj4/RvmuBWGAZLFsybc/jRx564r2MKb6+MjtRadeoO+ei9N/LqR4KGBJJ5s2fqxZJDthVmrIdscNy41BNAsCj1j5AJQAACEIAABCAAAQhAIHcCJlbo3/tawJeAIMGipukC+uwxc+r/Fyyiol0+b06WKRa/2PkRdn6OhcSGbBMrgv4VIV8Kx7Q7PKNCp50yUPKkkDBR2UKZGvLDkCAh8UJj0duKyqjQ3xqX81nXVKiUGJ2xdrt7iWVXHOkLBO5dvjnzsNhoz0y/P1DLjrU234lkKxnVMXg7z551hL0m787YuiWweVXG9hUL4rZv3lllp7+CGYkHzDzDa/ONcUXFJMfluOKrxvgzGiZlb1qV4N1q+ohn5/a4GruSs9ZprBIuNC4JEH4TJJwSVpGQI1kEMYVdE2yPeBGJjb8hAAEIQKBRk+Yt4+ITEmZNm2wlEEvellQhOaVBoybNRnw95NOSN7r9H1FOdk52larVa+xLD6YN7NqyaeOGgq5RpoyeqbwslJlSUPvczrft2KW7jk+fkne5J7WZPX3qJJ/Xq3+vHLKtMGM9ZIPjxqWeAIJFqX+ETAACEIAABCAAAQhAAAL/JBDKrNCqvrIbJCBIFEixsgaxPl+uv3GdzAcJCfoxv9wisqEW6R3TbMdLQr8pHMMIZU2oHJTu6fhWKJtC4oUEEJ2rYiEDT41H7WU2qrcdA9Z5wLwqLMPCt8QGE20ixXk5Pp+uVYZIcLM2W+2cUx4qeMzjzdwclblla/Sa2Wvcs35Y7926Pi4qkNwqPq5GlQoxNUyd8bqi/Dmu7KgE1w4re+ULxKRUzFiVWmP7nOax3p3Jfpdnuc8Tq8UI+VkoNG9HlHGEifBMEueY5qi2jjCkueSYSBEwoYMNAhCAAAQgkCuBFm3amfjucpVUwaJlm/YdtfA+Y8qEv8vSI9yxfevWhMTEJNMVEiVE5Dc3eVLo/OIFhfPwyNi1a6cyH/ZXrNC9lNWi62dOmZirr4m8K+Rh8cl7r794qJ9LQWM91OPj/qWbAIJF6X5+jB4CEIAABCAAAQhAAAJ5EdCiugQCZVRowV8/zDMtByC48G5b8LrdLwEGP0fbMbWXIKGDMt/OsfOOF4UaSZjQeQkN+i2h0DUKCQtavFeWgtpIkNBxCR8bLVRSQvsKFhItNC5tukb9BszDIpCaHDtr7fbsBjuzffLa0LZHrLCyURvNiDvDMi28MS7folh/ViBu59pdiasnb4xd8uemjLVLPDuy/Mm+2CoVoqPc0fGBTFeSd4vL7Zdgke2K925zeaJiXLHuWFedbdOSqu9cWC/Ou6NSjD+rcrQvc43da62F9soMEYMECSc2cS1aSIxwykZpvOKhNpqvI9KIcYaJFTqmTcKFrg2+aUm2RYgKOwhAAALlnECrNh06aWHaBIuJJRFFy9a7BZUZUyaWKcFi88aNKnXpqlipSpXMjJX5ChZe88RS29nTp0wqzDOSCCLRojBt82rTrlPXHiotlVcJqvR2nbqonNiMEmC4XdBYi8KBayGAYMF3AAIQgAAEIAABCEAAAmWTgIQGLfY73hFacN/u9eWYk4MJDSHBQsJFQDWTdi/KO8LD8pTE2C03ndZWx5zFeSerQGKFQv0rdI3u4XhW6Ae+BIsmFhIlZlvMs1AGg85p0d/JwNhin7V4oL51LC4pLsrbICZ+SmaOP2PTrpxE868IJMZ6RmV7A61TEqK9MR5XWpzbv8Xj3ZURlZUV49q2xhvIXJ0V8G7f5TaXipyY+KisxOQYlz/R5I+oQKI0GreSN3IsZWObK2Z7psttnt01ts+tkpSz2cw8sqvF+3amRvuzNb6VoZCworFWtws1F7GTKaoWNxwmmocjYqgUloQY7bdbOIKHI+A4osV+lYiw/tggAAEIQKAMEbAMhk5LFy2Yt9NWpkvitJq3btdBC/ZzZkybXBLHt79j2rxpQ1CwUMmrgvrwmDKgNoVlkJhUoUJhvC7yuq+EiFZtO3b+YdiXg/Nq08YpGTX50BpuF2asBfHlPATyI4BgwfcDAhCAAAQgAAEIQAACZZOA/q2vH+Q1LVpaqMxAZxMqokyh2DNjt9vj8vt9yn6YZaFa2hIY1h3eppZTFkmihEpLOSWS1K88HpRFoI4kXug+TokoLfDLL6ODRSOLdAuVNtBbpGpby6JeqE+JBLqPSkJVtdDiQFXLtKhuwkWKxUIb6ia7c2O7U6zt61hh6CouX3aUy+ffGfB7PQHz5HYnVXUHarWoGFe5nr9iTk60O8O3zZfhXm+VoOKi3K5kn9l1KJPE7YlyWVaGjdqXsi2hdmtfdOLKpJyNq6O9lt3hyzDBwW2lsAKay565yS3DJqkxbrbY7edhezsuYUKCi0QMzUvikMbviBPi4fQjdo4fho9MC1FkgwAEIJA3geSUipWOOfGUM1avXL504p9//Oq87V4WmGmxt4UJAj8N/+bLfZ1PVHR09BHHHH+SvfU/cc2qFcpgPCBbi9ZtO8w3U+fsrExlW5aZbfPGkGCRXLBg0bFbz16auP0bKVgaqqAttVbtuqtWLFtaULu8zjdr2bqtsjRmTM47q0W+ERs3rFu7esXy/b7P/o4v/LrCjLU47kMf5ZcAgkX5ffbMHAIQgAAEIAABCECgbBNwBIS6Nk2VV+pt2RQ19jhth+bu9phg4c3ZYecW2SH9AN5Yq0piTocm1SVGOCWglDmgTQv2TqaFzmmhXv4Y8qTQfXRMmRJdLSRUpIVCZtupFlrk1+cWFupT/hbKxJBIIKFD53UPp6RSrCWAqHxUI7ur7mO/XwJ23h3nioqNdSekxLiSq+8MeLMz3MnVktw5Wf7YjG3+hPWrfIlROTtzsj27TLSo4M7ONt8Kvytgc7XsChXEisuMTq5j3hVRll3i9eRk7IqXkuNxx0a5AzF7pJmQriN9J8cfHO/uclq7x6exyktDeyfrItEaxNt5ZZ04oo7EHi34KBtD4QkZeeu8H/HCKLBBAAIQiCBw2FF9T7j38QGvxcTExq5fu3pV/9uuu+zP30b/UBZAyXA7uDC9H/4QDz/3+vv9Tj/nwlHfDR1y57UXn3UgeEgsamhj/HLQB28fiP4PZZ/6Lun+FStV1r8t8t26H3H0sWpgX0H973iBW6069RuMG/PLTwU2zKOBPCF0asaUvLMn1CY/QWN/772v1xVmrJWqVK327JsfDVHWyW1XXXC64wmiezVp3qr17f2fGDD00w/fHfntF5/t6/1pX/YJIFiU/WfMDCEAAQhAAAIQgAAEyicBLa7LV0KZC8qwqGzlDdx+n9dSDZxkid0eFiZWKEtAWRbZ0VGe6Pi46MTN27MyKyfH6feCfqgre0D9OakZOqasCJlzS4BQ1kQrC2VOSFhQ6Lxj+O2IFEvsmISJZqFzjlm3npD8I1R6Qpkejv+GFvUlBiiTwfHX2OjyeJJdMQnVLCpaQzOp8Oxy+XK8gaydWa6t6zI827ZkmNLhSfBG+b12KCsnJ+D3+22alixhJhiB4MeoaG9UXKWs6ApV3e7AEo8/J0jGsjH2Ktu0x+FjtzgT3OyesXbcKbclwUL8lIWRYOec8lESYzR+zUWfNQcxlpDkiBnZJl7os26DeOEAZg8BCJR7AiO+HvLp6BHDvupxxFF973z46Rdf/GDwtxec2Lvz/Dkzp5d2OOntOgY9mmZOnZSrsXJ+86tSrbr+d9e1eOG8OQeKQ1vzUfDYVlINwYsybycrpUrV3Rzz2pTJ0u3wI4/RebEo6J5WYapirbr1GqxYunhhQW3zOt+6faeuymiZZ5ktubWpWadu/arVaqSaIfch9xUpaKwa/8lnXXBpp+6H99bnVlYCzfFDkYna64OG/lCtRs1aK5ctWYxgsb/fmLJ9HYJF2X6+zA4CEIAABCAAAQhAoPwSUBaAajUvsVDmRFNbpdeiuxbHs0yoiAmu4Pv9WnBXO3k0bLP1/F2VK8TlmFjhZFIEyxlZKMNAAoQW3yUeSISobyHvBi3eq/yThBG1kRDhhJ6A7qvFAZ1z/CoiFwAkgkjoOMpC3hcKLcjI/2JB6FyaiRMmjlgX8qWw1/WUXeHyZue4YuJjXTmZ2W6vRebWXTFJtX1J8aZFJGVmb3e74nb5cpRB4fV7vR6f1xsUSqK8voxY787NCTlbt8f4MiQ05Okx8f8Sj64MbupD85YAo0wLMXLKZYmNOEnE0CZPC5W/cvw61FZZF6pdLrFDWSVO5gXixR7EfIAABMozAS3e/vrj8G+XLV60YPCPY6decfMd9919/WXnlnYm6e07drH/HfLOnTl9yr7O5farzj89tVaduksWzp+7r9cWtn2HLj0OV9s5M6aWKf8KzSkzI2PXlk0bN1SvWat2fjzad+5+mEQItdECe0Hsmqe3ba82s6ZOUmnN/dokZMkvQ9+N3DqQ4baO709mzn4NKJ+LChqrLnX8WaaM/2tMuA9IlKlBsXHx8dnZWVlD//fhu8U9NvorGwQQLMrGc2QWEIAABCAAAQhAAAIQ2EPg0Y/HaxHdMcM2bSKgkk++4Gr8HrNt6QUBn5VEWh0qB7XMDqyvnBy/08pBaQHdyShwshwkKOjHuxbpdbF+wKtL3UclofTjXwv1ef2w1wJ/fiaXup/6kOeGxq9NoosW9iW46D66v3lZuLdaakjQqNQdEx8XSKpsxyx9JDsjyzQYX3TAl2kVHHKiK1X1RVXw51h2RZTfH4g17wu3L8e6zMo0rSPHBhrIUUEsryc2JicqPjban5UT5fL63LtNyIObM5lwJcPJupC/hQk8sWojrCodZX9rS8j2B8UZx89C8xA3xwtExzV+7bUwIZ767MQe8YKSUc6TYA8BCJRXAosXzJ09fuzvP3fvdXTfssBAC896i35//CEydu3aeSDFCvHt0LXH4Srfs3Du7BllgXfkHOSLYi/3y2srz00lyfSPp8KIFeqkY7fDjtB+f7NSEhITk1Qq7H8fvPVKXoOSSKAx7U9mTnE+x8KMVfcb8fXnn8ZYTbehn330XrgHjT6f3bdH0K9DxvPFOTb6KjsECkxrKjtTZSYQgAAEIAABCEAAAhAo+wRMrNC/8bU4rsX/jhbyklB2gx3fLVlYxJt3hQQEr/0YX2F7vampLIZ1V57YalfNKrJi2CNISLxwPBqU9aAf+Sr3pMwAlXFS28YWKj1VlE1jlg9G+EtVupf8MHpYSBQJGV8GZIC9zkSKHFdCSk13pTr13HEVKrjiEuPdCclxMUkprtjY6OyYmOishOTK3sQqNfwJlau5ouISrOBVrCcqJi7oPe6yP3JiKlTaFl+r9rb4mtWyoyvE+91R4WWqcp1PuIghFchKScnjIrg3oSIYtjmikSMciY+eg8pnyc9D9bMlaigk5GgvQUPz17WKKCsZVeCbnUWBzrUQgAAESgKBmrXr1tNb13mNZd6s6VPlO+C89Z5bO5XxyW+BWefjbJW0sPNVW5W+adyspf53tNBbfvMwMT2uWavW7Wbuh3+FykGlNWkmD6gCt+joGEf4L7BteAN5hmhhfNmSRQv0Bnx+F4u1mO7TDfajcUHPdV+7NMFiWarVb8rvut59T/iXjM3VpjCiRdfDjjh6uTHbumWzslVz3fJ7Ji3S23WQGfv0yXn7V6S37dB52eKF87fZTQoz5+Lm5tyzMGNV2507dmyXAKOslsjxrl29ckVJFCv297+bwjwP2uwbAQSLfeNFawhAAAIQgAAEIAABCJR0AhIQlIkgM+vuFkeaNqFSBfH2xmTwt7fCSjI7C+EqV7TOQkaU8rzQcS3aaxHCefNfPzb1A9nxYNDCu0pAaXFJ4kVTC6fc0/7yCY4rFE4fur/monvpnprbSmu20VYQfDYLW+B3B8yUIjsYMfEx7qTKiSZaxEZ73DnmS5ERsBJRvuwsn8+Mt3N27XSbwbjb8iKCKRH+mMSUzNjK9XfEpVrUSM2IqZjsd0cX6TdSeCZGCLCSL/RRJbWUgSKhQoKFRB4JSp0ttBjW2HSOevaEUm3FT+kKAAAgAElEQVQfXlYr1kSLOItoxIv9/WpxHQQgUJIJJJkK8eXPE2afffEV1+U1TmeR1tbT9/gJOW1l4PvaJ0NHjpu/LuPnaUs29AiZJUf29cBTL7319uDvfnaOS4h4+vWBgz8bOWZK/2deeUfjcM6pj5Hj56z46Nufxw35adyMwT/+Oa1+w8b637pcNy0OX3nTnfeNmjR/9bgF6zI+Hf77JJkORzZunt6mvRZFp0+eMM45J1+Ca2+75yGNodcxx/XL6x4PPv3KO+9/MfL3/ESCo4//12ka6/jFG7O/GP33TPke5NWfxnf9Hff9990vRvyma66/8/5HVK5KQs2CfLxCJBw9+PTLb/8xe9W2sXNX79C8I++hxfe7Hnn25SP6HH9S+LljTjj59Gff+viL8y6/9uaCvpOFfa4F9RN5fvWK5UutqlaeXOrWT2vUqGmLVj+PGDZU16qEUX73MI/yyu27dD9s7K+jRubWrjDPRNx1rePzENmPRJNW7Tp2zut8ePvCcFNZsUeef3Ng+Hda36vLrr/1Lv030fPIPsfnNeeCxprbdZWrVqt+y32PPP3ukOG/Xnf7vQ/nx/OcS66+QeMIb9O0Zeu2T7zy3qDbH3xigDI8Cnrm8mF58f3B3/5i//dg9JRF65589b1Pz7royjz/70thnlHXw3offf+TL74p0dG5v/4buuu/z7wUybKg8XG+YAJF+sd4wd3TAgIQgAAEIAABCEAAAhA4WARC2RV6q1IiQppFR6se0Np+bGvRJMrKP9nO1vf1/1uNJNtJoJCvgjIlJEg4dZMd/4pg3SgLvWWpTAv9aJdwoDc8lfnQyaJ56NiBestSY9CPU70Vq3FJPLHP7qomOkgEyHbJh8MTle2OS451JacmuyvXjbdST9nujM3b3aZWmJG4z36I7zYNd3ts8SHKFWX+22ZqEWvG25Uts6JWVkxKjeyoxIpWHirenLmD2Q2h5+awKNRjDE+HcMSL0F58nHkkWTtlXOgZaQFM4lJzO6ZoZqFjOqfyWGqn5ynhJtFECwkYMSEBQ6WjyMAo1JOhEQQgUFIJZGZm7DIdIq5O/YYSp3PdkkxNUDmcyDfYO/fodaREhbRGTZsPeu/1F62rXfc+8cLruXXSyt5Qd4737nviyYOG/zZRC+pJySkpp5xz0eXWhXyYXCpV88gLbw6Ul8Cbzz/x8M8jhw1t2iK9zd2PPpdruR4tYL48cMh3WvCfMmHc2C8HffB2i9btOlx89U23R44j3TI2dMwRLLTQLUHkmlvv6a8xvPDeZ99oTv/H3nkAyE3cXVzS1uvFFRuDDQZjem+h9wAJNYQSSIBAKKEECCEhEFIgkACBUEMJfJTQey+ht4ReTbNx7/b1skXS937aHbNe7uw7WmwYwVi70mg0ejN7d/t/8/6vp/7PmTVjOgHS6hJipbTeT448/uTzrrzxzq6Ojvabr/nHRcsuP2pF2u2prTXW3WDj20RS7HvwEcfMnDZ1MtccduzJvyUgS/33iuqC8msHDx02HLx32u0H+91/x7+u+0CeC0eK9MBwurTuGuusv9G+Pzn853vs9+OfmuP7HHTYUZAVkBYny0h9+133+EFv492fce3vvJ4xbfKkocNH9EpYbL3jrrvT5uMP3XMHe8iXRd2D+pBQLzz1+MPl9fo6JqQJa2maP683026IBdRFi/Ov6Ctuu+6930EUQ5BBiJz196tuPPbXvz+bcbnwmlvuHTSkZ5+PxfW1HAPmOHPtx0cc90tSZx1+/CmnQwj1hCk4Qmwc8vMTf23Oo3K69q7Hnt9pt733+9FhR/+C84saD+YZxN7w5ZYfdfXF5/35pn9e/vctttv5e/sfeuRxPV3X1zE6+OgTTtnrgIMPH1X8OQFxx332Pfhnx4Dl366+KSK47PblIPBVfan4cnpnW7EIWAQsAhYBi4BFwCJgEbAIWAT6gwB/3xPYJsBNCiUC33X5PBYKUVoD/VsInweBz0FUFR+pSLUQkRcFRqOwZ4MsoEBWsKIMZQABJRQBpFOARCBNFAH+Xg2ri219GTv6YtInQVbk9VBNYiCyjldJQKHaJQ3G4NG17uQ35rrtc1viNUMHVQ0c6gexhJ/PdMX8nLgXP++EGblVyNcykpDEUvU5r0JkRaoiF6tMy8siH/ezeWkwwKFc9fF5n8MoV6Lri2DRZ0gMo76Q/CPy7OC+mHajfCG9BGPDJZBKxsyb90hmsiItfHldmDH7vP2z11kELAIWgf8JAhADM5WnR7HwXtP0DBg8ZGir0u3grWA6OUxL4QnQT5k4/uPD9tlla8iM6VMnT2LFM6veS1Pn1DU0DkBRce2lfzuHYP25V1x/+0fj3nv7pMMP2EvXTGQFeNO8uRD4zqZbbrfjgEFDhv7mmEMPeOju2/7FMZQIuVye34Wf2U49+4LLN9586+2p//A9t99EheVXGL3yAT896vjL/3b270u9KtZab6NN2ttaWyaO//B9SJBLrr/rYfp/6N7f3VK/vhKoPX5w4KFHvvLis0+V30ip/7Pz5s6e1VPaoa122GW3437zh3Puv/2m63534pEHy7spkLH0cNIIlbcDmfKPm+57nD4cfeCe3+W5CVhffN0dD5qV9W+/9vJL5dcRTAbvRilCDtlrx80x5eYZUGeMXX3tdVEumGsgLHj92n9eeJY9aaZO/v05F0L+PHb/Xbed+ferbqDPvC6/T3/G9fNMWPrJ/EBRY4yhS9vZaqddd/9o3DtvTSoam8cXo7DYbpfd92aMX37hmQXqHdrrz5iAz6K8KThPm+++8ep/e3vm/uBWPj7M1R2+t+c+EHSkNEPhsNk2O+x8103/d1X5/RbX19L6qBJQOjAfzzntpGOee+LRB+9++rUPfnPW+Zeec/rJx4Jzaf3Rq6y6OoThM48/fT/HGaO//uP622crhdQFZ5128q/PPP9ScP3zqSce3RMOkGGn/Oncix+869Ybf3/S0YfqI5PleX567EmnvvrSc0+XX9PXMeLzAXGij27zxx+8F3m7nHHepf8cLKXKb4877MCd99z3R5tuue2OI0auMJrUYJ9nXtprFkbAEhZ2RlgELAIWAYuARcAiYBGwCFgEvgEISF0RBexV8H1gTwC7Jp5IenkZTRfICjY3UhgoQDRBxx7TgVdUICwIxGAwySJWQz4YpQEBcwLln6gQYGdlorkP9+2XCuELwM33FwgS+kKf6vVg9fKiqIocr12XFFF5p2bwCHfgqI54am5XvKbeSaRqHflaZKUqSXfNnebm5011Krtniu7oltLEd91cVzyRaa6ryDYPkMLCF3GRjQW5mJJNoSyhIEepF7khEsNpFbCtep8pIgqRA17gRzHEhDHc7vVxF4yIWyBFdBPaivKOq8FKHazmvjxrsa467cwtPjuEk7lfINLCEBiQFwsCel8Aa3upRcAiYBH42hCYNnniJ4vyFVh57BprffLxh++Xdui35/z9HwTRf3HofrubIL5inRDAjq9fcqV1N9h0i62VCtF7/eUXnzv7kmtu+vC9d948/Ie7bEOefeoZsoLXw0csP4o9ygPTxqXnnnl6T2AQIP3+Dw74yTWXnH+2ISuo9/ezz/i1yIlNy421IUtI66MYagVqAwKxh/9w120MuUK+/2WWXW4htYK579g11l7v3Tdee7m8H1p4X0+6qw/efeuNP5x8zGEEh6kDFvm8GPqSjeDtOZdeewv+FMcd/MPvm+fm9/69t954LYQFBFJPK/kPOuLYkwjannzkj/eBrKBZgss94b2KCAyOQ1CgUKB/GI3/6sif/JAg8s9/9bszxQnhtfWZrT/j+nkmKB4WXDdsxPIjywPmA+XGvfb6G3/nHyKawITxY6x6uw/pvDbeYuvtn3jovrswRDf1+jMm1CXQjUl1b/dZdc1118esWrHyN3ur0x/cRFqtO3P61Cn4dJA27KiTTvsjfhOXn//nM1DLQFj0pLDoS19N//BbOf+qf92F6umI/XfbnvnJ/CP4v97Gm22pzFujy/GnX2besGee6J51h/1g563EK07YRp+3Xffc90DaKPlbNbolHi8ohF77z/PPnH7CET8x5Oa6G26yOfd9+rEH7y3Frj9jNFydReHywJ233MDnY9udd9sLsuOknx24978fvOcO5jiEBZhZwuLzfCo/e40lLL4cHG0rFgGLgEXAImARsAhYBCwCFoH/NQL8bW8UD3F9kSO4HpNZxQKyAh7CVUokV37bsoDAj2KiCumgCNj4px6wfnjqAaEhH2gPNQNtcp7APatPuaZVBeLgM7nEv1IQICWCfOBkO+l74KRrGyKSwlU/cpkuR4baTiyeduPJwU662vcCv0OvazxUF6mUV12RVNWck+ue66Q6pjjxXIfjKU2Wl+twY7mO6mTQuawfejWSYQT6JpyQy4cvMDIiEnzRAQ1CJqceNOlYh0onpIX6EeWa0nvIAxOsgMShj5AK4GmUK8BTSE1VIEGi1zxWsQ0UH0pWFW0pHUyJZwLjiExSvbhaS6tBCBva5n6oLkyqX45lRF6wX3BPERhfh/rlKx1627hFwCLwzUYAlcOW2632vZ6ekpz1o1cZu/oNV17yN3MeRQM+Exeedfqvpk2ZBJkebWNWX3Md2jJEhDlOgBQyAPUE6aUO2XPHzcvrmLqG/Ij8Hz5DD3zaQ1JBnXTG2RdgIHzFhef8sbTvb7363xcppccIqEKGPHjXLTf+/OTfnanY5rL777zl+qVKEIkskigwynGAmBFns+6VF/71T+XnSLVD28cf8sPvQwZwHj8CrVZf46Vnn2RhwoKN9DekFzrvD78+gRRTpefa2lqi+7731uuvlBslk/7mkKNP/PXzTz72UKkqYozUGlzz0bh33y5taxWNA6bKpDja+0eH/Axfhf2+u/m6pn/qXo+m4P0d18/zqVCgvkBYSKFTHjDfbpfd9obYMuQBc0TThb93etx23++gQxkbjekNpRX6MyZ4U3Dt4hQWKILKCTBzz/7ghpoID4s7brzmCq4/Xsqc+fPmzL7gzNNO5v2ijKf70lfagAy44Oqb72EliSErOL7z7j/Yn+A+Qf//PPfUv8tBZd5wjHlG2qh9DvrpUX8+9YSjICsW9O3TFTgLXf7rP513SVo/LM6QsqJUibXp1tvvxHuIjM87RqiSuPa5Jx55EGP6E08767xH7r39ZsiKxWH2eeaovaaQg9ZuFgGLgEXAImARsAhYBCwCFgGLwNKPAH/bE9wmOE0goLAisKdQdUFAwWp+0kehmIj/9kcbdIis4DjBdnM9fhWkliJATiCDlfucM+XrRS3IOWHLTCec/u5AJ5Z0vDFbin3RY2fEHcz6MOE0SPRRPdAN89lqGVSMdpNp3/GzgdM603Hb5sRq57/vpVo+cHIdE5yKjvEQFYInpsRPgRPzu6viYabK93H6cAn45MXtpFUBTiNSUAi2KEVUzHNSet0pxgGyoEskAoQBuPHeKCsIiKACASuj1GCla0RgqEHSP0FEcMxcg8tIZC7CHYtSjSr4jOg4fJMbqWdol+vmFa9l3Lk/BAbkksn9RX9RX+Rtyqivd6rau1kELAL9Q2D6lEJaJlZClwdlN9li2x0IEr4hdYRp9aAjjjupef68uTfJq8EcY0X3dt/dba+rLz73rPK7kwKnXQF5AqB//NWxh0My9NbD/z7/9L9Zvb35tjvtYlJC9VR3930POnTosGVHsJq7PMDfU32ThqdTQfBDjjrhFMiWCR+9/56pS1sQDZM/+ZhUjQttBHLB5q3XFiZBMMje58eHHfXsvx95oNTIG9UHfhOkiDINVcn84sDDf34ChM4t1155Sfk9qM+xV3pInbOXSAeuv/TcPy1QmnBvfDoIBNOmaY9+jlpx5VXuVDohSJ1DjznpVFbvf1Q08mYsFTIfWk7ocH1/x7V/s6xQm3mDwqTcd4NzO+++z/6oDiZ/Mj4aA1JGVeq5e7oPxMZe+x98OO09/+Sn/hX9GRPaNd4q7775OorXz2wE+AmYP3DnzQuRIqUV+4PbyquusRbXvvzCs09CJG2/6577nHjYAXtmNIk5vkzR3wNPjfLOLK6vpj4pv0iLhvoJZQXHeQ7jTQEp1hMxN2bVNdeeqFRckGm/FBn4wbtvv4EnjGkXEpHUcOXqijGrrbk2qblQNpX7gHxHqqEPlXqqlKDs7xiNWW2NtQ1m+LLgJXPeH05d4FFjTNx7wuzzzFF7jSUs7BywCFgELAIWAYuARcAiYBGwCHxTEICgwKB5WZVttUJuU6XEqPRLUm4XPSxkX5EnqD1RZbwKQXYC6tH3SRVDWKT1GhIEYgPiAnLDtM+X3a/f7FnkgUL3lU7LLFEH2dAZsSbdCMPWWa7bPDXhVKqL1YMcN1XtOq1vueGMcZ5bURu4sYTj+jnX09MkqtNO0Jl2vO56J2yTcCLboXM8PmIKSRikYdAXYYiKaItIA6Git7HogfWPlBds1TpYoQLxEPoiE/S6jnMStXgiF4ZLC2KIinYRDahSIBSiNFtKN8UVkA7UIeUTgYLuomqDNrkL6o3uiNgQs6IOQFbIFNwRrRKRJ6TiEL/iJFDT6DXEEkE4CJDSVFX4XECOcI31uygMrd0sAhaBJQiBmWIs6A6qg/KUKtvs9L09CByLSHiCOgTWN9psq+3+77IL/mKCrCgXLrn+zocmKW/UtTpe+mgElkePGbs6QUqC5vfeduO1i3p0UuWgTNhmp133KPW2KL8GU2kClI/cc8fNfYFydZEmBFox/B6v/Eg3yiS89LqVxq7GLzWHdFXl7a253oabsEq8PFXT1jvusjur2W++5vIFxA1pncjjf99t//q/Ul+F74nEIK0N+BilQ+l9zOr2nnL9Q4Dga0GgmWtIBfXXy6+/Da8Pgt2l7YA1wWnIle/vc8BPUChcccHZfzB1MAPnfPk493dc+4J5T3UYgzmzZk4nJVTpefpFyq7z//CbBYFoDe9c/C56agfDakgP0oGRrsnU6c+YcA2eEATo586eOaOn+6wopQF4G+zL6/QXtzGrFoLvb732nxePk8n26/994dmnHn1AaojCtrzc59njrVJ+r8X1lfp4YYDNrdddeWlpu7vs+cMfkfqqcO/PeqSQ5gky5fEH7749Ih9FQJAuzaQ447qR6ltPKZf2O+SIYztlHH/bdVddVtpnxgelBib0pcf7O0YQKZByzcqhdvDRvzjlun9ceG6pQgnMmFcSe/F3td2+BASMdPhLaMo2YRGwCFgELAIWAYuARcAiYBGwCPwvECj6V0AoDFVZRmXtRKpiVa3HT4qdKHZJ0X6lglJsPacvf+SexrjREBbmi7Yx2Yao4HUU4FYhNdSqKlurbKGC8fbXv3kx103Xel6QjXnNU+PO7I88p2M+7hxuWNUYOIkKNAjSmYi76WxyvJlauDp3fOi0zHDdfNYNKgYEfuMKYTh4JSesW9ZxIThEZvhuTKxB0ukQF9IdVnX6TqI9cL3u0HfySBuK9h+RR4SIgjAnRHKBLlPKKJEFpKSqEJmQFlHRKFVGY+jJdyLmDE/EnBVUh8IX9Kjo+hW1X0n1xmq/mt5jYL5K8fxI9T4qajMqYjRG5MNI5VItMqROI9ige9VpcBrU7lC9HqX6y6mdZVWWUycxRqc+8wCiiUALKhpj7l0p8iKpElPxVFwVh2I3i4BFwCLwv0LA+EWU+zcQYCdfPGmIjIpho8232g4SgnzyKBL2OuDgw2959IVoFfdRB+yxY6mXAMcIkkJW8PqfF5/35/LV2T09M0F9rtn/0COP6+k8aolRK40ZC/nBav2+4LbG2gXCYq31N9r0nNN+eUxp2hquX2ns6kXC4u0eCQtWiROULb3XJltuuwNG3C8999TjEBcnnH7WeRf93+0PvPz8M0/gZ1FaF+KH+/e2Un+dDTbZjD6VKlm4nqAvq+XBm/cYKd/yyAtvbLDp5lufeNj+exrlhLkXq915Pe6tN1494KdH/wIsS9NerThmLL/3nAkffzCutH/9Hde+YN5bndkzp08TN4Yf14INcoVURQ8WjdY5MV/YQsr01M6PlV6L+rf838Jqlf6MCe2uusY66/VGRnAe7xL2vdXpL26Mj/Eu2W7ngiqh9PlWHLNKj+PTl75WKt/aiaefdT4qiVIFAqqbI0849ffmMzzunTdeK8cUwojr8Wk58LCfnwBpWGo+X9fQOIDUZ+XzhuPf3W3v/e699YZrylUb39l6h+9ynzde+c8Ln/dzw3UoLGR4/vIOu+6xD94w119x0XkLYzZ2NQiN3lJ2fZG5+m291qaE+raOvH1ui4BFwCJgEbAIWAQsAhaBbwQCIitYiU8gBnPmgSqkLghz2e5CWqEFZtvktE5ImOB36tADqsOXN2PgHBl0cp0K7VFY/U9qpMgXQYXvDpAi1OVYZLT5tW6K8juVir+LeAlbZvvBzA+7vBUHVrjLjEWxgHV1UfUBaSELiHjcD93E7MBLpp1UdTKsG5bLdA9N5dzainRXtxPPdDp+Lu+0J4Y4ShzldHkV+Y7EgPE12dkt9V3Tqyv8poGyJx/sBU5Sp5tECIADrE+lkJorVUWzjg0VkQCJkBLvESEookNppiKlhWQRSh+l61WvNvLCKOAq5qVori2Fht6jrugs4ryQ34WehHuiiGnSxXm106V7NKPq0O1qpP6okJIjEKkRqE0NejQ+jSoQFFxnUjpwb/DhftSj3YiEMaWEtECFYTeLgEXAIvC1IWBSNBnDa3PjXfbc90esLkctYI6tu9F3tiBIjyLgwmtvvY9rIDT+dMpxPysNjJv6pL3hNdc89sDdt/Xlof6r/PqkOvrhjw8/mhX05UTB1gr+086j9915a1/aY/X4amuvtwFEC319Tavay69bWQoLVpN/LGfl8nNrrrPhxk8//tB95cfB4p3XX/3vYcee/FvSPWEQjWH0VRf99cxSQgQM19lwk83eef2V/5SaiZv2MI+GMCF9T7m3B/egXpdAuPqOh59Zd8NNN8f74YBdttoApchnn2P1NVG+EIDG+6JU/UFdVryzL1eS9Hdc+4J7b3Xmz50zGx8Hcx7ia/cfHnjIUzJmnif5hTk+Z+aM6ayu7wl3CB7Gvzy9WF/HhDbBB0LoHgXbe+urCIvI++Pj9z87L7imv7ih5Pngvbff2O/gI46BFChPzcX4yEaluXye9KWvhx9/yukoPo4/ZN/dSoP3zE2eE9+HHb+/9756loU8T3iOlYuEHXieePqZ5/1URtulmKyoD0hh3ixM6EHEQYiQgqwcw8232XEXjr356ksLERb9HSOeCcwOPPyYEyDgSj8jzB18YZ574tEHv8ictNcujIAlLOyMsAhYBCwCFgGLgEXAImARsAgs3QgQJkcNgccEaYeGawFlY0jEHK+KYgg/lGN0MT0UKaBIvUHqAVIU5eVfwaJLQ1QQ8Dbpg4zx9vI6hkKAL/fco1mFYDgpor4+4sJIHeqHTw4HzJ3pVg9Mi8AYLhfxAZ+SFeoR9YauNkUPPMdJ12dkzu2Gyaq4iItkS9De0JxKDY8Nr3f9qrXcTNMsJ9PRJmVFUg9WHbTFa7obOye9vcLc56cPDj+OVfjNyViQF+EQ1gpNyAYMtwn4Ay+kgPB2qhX1T7qBUwWBIRpgkEBswf9Cg1Oh+pXqUkp2GzG1kSw4bRcGTaQGCg08MapNqidUHJFsJJKOyLvCjciFdh2PFPIiR+BXKE26xzT8NESaBCriVpzBeg8RxRjOx18DckOv8bkgHRXj1qHpYVYE++qDSV0VeV4wJ0ReQGQE1vsCxO1mEbAIfNUIKCNO5CkxbMRyI829SBv0o8OO/sX777z5emmAf+31N/4OAfY/XXjl9Rz/3QlHHtxTGiPTzuhVVluD1w9KIcCK+L4+y9UXnXvWJTfc9fBuCmTf9M/L/156nVJSbUtQd1Er40vrj5SnA2oR7n/ROb//TU99WFmu2ngnlPthDBw8dBmCvW+8/NLzpdex8l++0StQNtt6++8+fO8dN19+3pm/MwbFpXUJQmOm/GqZ8bCpg4oFUkUr0Re6B+fBm/3vz7/sGtoG7/vvvPn6coWIaWvlVVdfa8JHH7xHyqzrr7z4/HKyR1CsRgD+k48WVlj0d1z7Oo491SOV1+prr7fhguf/7vf3lBP1sDuLRtTmOKvmBfMwfDdK02jJlyMaw2sv+9s5n3dMuM6oUd7vQXGwAE+t7v/4/XHvlKadKr1nf3DjOUYp3dKbUhzgwXL0gXtGCoTSDWKgnBToS19Jn8aYvy6vmadF/Jg28WbBsJ3j4iIm8wcnCozy+zJvovm2wcbfeeWl558u9WTh+KeExcIp076juc84lRuoo7zYdKttd0RNU0q+9Odzw32N54dSm9Vi1H7L/12xkP/LciNXXAlce8Lsi8zRb/u1lrD4ts8A+/wWAYuARcAiYBGwCFgELAJLOwIEsQlEE5Tm7/tVtIBzgL4PRtHuiLGI3Jo9R54WWcUjIBuMP4VZkQ8GEBbGw8KkhjJqitLjECSR74LaVVA7LKQcctEXlMg5vkpUh60+360aOMFJVyflUQFhAnGCNTXPkxeBEXcal8s4lfWQC1kvUdme81K57s7Oqub2inBOqnpAumrZiq6KlZyWimanu3mu0+ErJZRX5ead+MA5NWMybRVDXxjR9Gr70Na324a2fhDEndwyEfcTKuDvOm0QDHpHmog6oZzQ+7ju3KhzI3RsuJBokaKiTggN1zUcp/GUhoGxSooWSEihIdNwxxejQGqphEDGd6IwCmZEUGzoXrSlenFUG5xXW7hzN2uAGnWc58SsG7uNOSI45utNRsdn6hhEC4qQCvWJR0BxgadGDs5EB1B3QFxRIi4lwrCorMGwW68XmIIXzy8YXavE+Conum3bIvDtQYAV+ZgXDx8xcpR5anwTWKV/wk/3j9QMZmNl/Ltvvvby2b898efvvPEq6Q0XuRnD3EfuveOWxdUtPf/C0/9+BFNsVt6XEhYE/gmuYrRcmvi2FeEAACAASURBVF9/UW2vvk4hOP7AXbfc0FMOfsypSbv06P13fUaxQQoprn1TUdyFcRgWKQQeuOPm6y/+6x9+25NywtQnSM3r8nRP5vye+/84Sh/13luvfcb4GbwZGxQsTz5y/92Le2YIIlbJj11znfVOPHxhfwvuQUqo8R+Me7fcR6O/49qfsSyvC2GB8TckDQH0g3527EmYNb/4zBOPltadNOHjD1lBz9gY5QspmjbdctsdwWLc228ulNoID5a+jgn1jJ8E5tI9PQ/9U521pAy6vbfn7Q9ueEMwf9eSJ4rMxV/Dl6S0XcykSbv04F233lh+v8X1dZ+DDjuKNGpXXnDOH8219P+Mcy/5ZyKZSJIG7fhT//gXFCzGe6b0Hswb5tmue+174K+O/MkPy+9PqirGCgKz9BzP8uLTC48b53eSkgNSrfwZ+ztGo1dZNSI8IQVvvPqyC8tTzpkUZ+Vz4YvMT3utNd22c8AiYBGwCFgELAIWAYuARcAisLQjQBCalf54FqyksoYXS2gVJ1mbivIKnpDV+k5EVlDwoPikMh2fMaiugu9/hqCAjIDMIBjPinxW4+NzASlAOiiOQw6wF2kRTnby2XbxFCPkBVFdIC2++s2tH9bg1C1To/u9L3Ji5II7ut4U9WmO3g934skKt3rAQIXfJ+l9u5/x/eausCrrJsNUpdcRi3lSNaRi3d1xZ166wslk8+IQwrgbiy0fuLlVZjWO/c+cxpWbKrM7zj1w3E+alARrUsgTd0WKB91WqaFcB0NKSJ2UDqX1vhJFQ/FYXKQAypQ1dYwAXGSgrfRQw/Sa9yN0HIKpXWoH1DEQP6SWqligilHLCGXIhAVZAR0ED+WLQsC0G08LIV4rZQem3/QjI6KCtGCdqhrT+dmqP1Vsw5SIs3IjcgLChH2gOtwfxQ2KDI7Td45BUBgiAxIItYZJZxUpL1QgNkwqsa9+0O0dLAIWgW88AphdL6P8Tjyo0sRXHXnib37PquVS414C+5zDTLovZAVtrbLaWusQQIfk6C+I999+03XHypiYoLBJ/YMKhKDvdDns9rU9PC+oe/v1V1/e0zUEY1GUEEQuP09AFmwopeeUTSgi6x+657abFkVWUIdANPupkyZOKG9/o8233s6s9O/J8Jv7oKz490P33rm45yV1DibVFPxCytNLgRvBf3AtbevzjOvi+rKo85hpQ0TU6uEwtcZM+qzfnHBUub8JhBXtrKi0YoawOOaUM86i3uXn//mM8nv0Z0y4ltX7UfqlsrE17bKin5X9H8ssvqfn6S9uetQo+E76r6MO2H3H8jaNiqEnxcfi+rrr3vsdNE2fCdJMmXb3PfhnxzC/zv39Kb8g3Rj3nza558/NSiIsmKekqOopZRp9m6Z5WOpTgYoCBVK5uoLUa9vstOsevh/45Qbf/R0j+sXzLLv8Civecu0/Lu4ds4XJqy8yP+21lrCwc8AiYBGwCFgELAIWAYuARcAisNQiIP8KAsz4V0AmEGgmuNwio218LCI1NUoLV8vyld/XyXZ3zdKhV1WmJOJe2+arD8sNro98SEvNtiEsuJ5SUFI4zjQVAv8E2gmsQ2Dk1HBKxIAMuV0F678mdQW9db3BCuqP0SvIl+gBoi0klC9KwY2jFiCwrrRMGXk7xAYlEzGvujIhEUamvSsWNPtuUmmkYk53d7twyQmAbicWdISV7tysm+gSA9Fa3RCbtsqw2vcGdW83eFZ1OHuynhifiVBURRBMcfLBZCfrVuv1bKczbOeoMMdLo5hWSfs5ekfqLYyxIQQyGg7SVw0naZXeQwoxTqSJkl+GU4lKQu2kta9X3YG8F8mBP0VeJEVC79NxT9egzeBG0maAvKQVMvZwEiIsaBOvC1ev8TVpIEWVpkCN9ig4ZquNqbpmmtppFSGSFtnB/bNR6ihX6agKZASMF89LAU/mAWoLkz4qSqtS9L2gfrRJcbHgtTlm9xYBi4BFoC8IzFC00xgMH/rzk35D8JtV/aVBZALMtJXro9E1gXPSKd3VQ377vvTJpGFilbUhLEh9w7VzZs/k53ufttXXXn/DuarfG8mykgw5aKg88MqxtdbbaNM3X13YNJjjn2KRXazpd2VVDb/Tnbkl/gy8J2h/4mlnRgbCeA6gfCh/IO6D/0dfHtSsRid90U3X/OOi8mvI9Q9pUe7T0d9x7UtfFlWnS4YcnCe1GObZmFD35CNBii5SWslCZDP8F9bfZPOtNtlimx143VMKoP6MCfdfYeVVVp3wYYEU6WnjPMd7GpeF50DfjN9NejTwL1eT0J4hLOSH/hkflUX1ddToMWNJTXbjVZdeYD6vG2y6xdYnnnbWec/++5EHOI6hNumYXn3p+WfKnxWPleG6nuOkEesJC/pW/jlQtqmI4Jwlxqf0GtK45SThgdzEt6X0XH/HyGB27203XNuTRw4pziBRyr1Mvugc/bZfb1NCfdtngH1+i4BFwCJgEbAIWAQsAhaBpRkB/p4nEE7wOhaRE647P/Dzg7W4LF54Ly5CqZuUN5uV9G9p2f1/pC6YWVeZnL/+mMEElw1ZQTsE/01hNSZBf77UE+gg2G1W4FOHeypc7nHd16KsKBko3T9cVgSFgujewEiCwBbmqlVEZkCikLIq7zthtpb3kk4ka1P5+Um/o6UzbO7MOHVditKngsrOeLxripiEZhlwd4apcH6mMjazqjE+efVKt6W52pvTHHOzQ/1Ycng8nsWXok2lJTbS6YqtUDDQJq2T/uumdF4t5QNHcwr8D5aHhOdIgSLDbjwu5D2hktb1qDHAEOKHwBcExhDJFZI6B+aVGrrB2g+L6hewDkRAMAZVeqpaAY5iA8VFVqbbqC8SRRUG9yHllBgVJ63XVSIzID8aRFpITuN0iaBgle4ktTpLbczX6ybdoJ3UUjqf0bEgeqYCiYH6g9KuwpNBipkUUsbrxAyNKwLD+GBExIVNGVUya+1Li4BFYJEITJ8yeeKW2333e6xoPuiIY0/694P33EGws/Sizo42lH8OqWf6AqdRDqDIWFx9VquT6qmUVBDhH/2CkfUEP++ijTQ37CsUZC1vU+nsx7S1traUGjfTLkbHj9xzx83lK/jN9ax453V5oJjc+Kussda6j9z32XRWnR3tRSwkE1zMZgyQ1eVK0iGZ6gccetTxBGRJ0aPF8eN78kngPvLyXuw9aNMYnD/58P13Q9CUd8ukzykP0vd3XBf3vIs7n89mIeUjv4TNt91xl8vOPfP0UpNocz3pr95+7b8vbbTZ1ttxDLUNWF1w5ukn93SP/owJ1w8ZNnzE808+9lBv/R2iiDznJn3y8Yc9369/nwczPrddd/VlPbWH0odn1u3eLz+/qL6uutY661Pf+E5ALvz1H9ffDgl52vGHHxQ9q5hD9qUKCXMPPFZQRTBnSLVVfm9IQkr5vDFEnPixBZ9PWcXUY0L/0N23/mujzbfa7t23Xo/SnKFgIkVUf8aIz7ohcW79v6su7RmzsastinRa3Fy053tGwGRHtfhYBCwCFgGLgEXAImARsAhYBCwCSxECUldAEkBYEBgmoExaKHInc2xBqh59QeOpugI/91Q85v27uiIxbtiAqhkrDq9j5bxpg0BEYTV+IYhOYJwUU6gY1lMhf/Y6Kqx+gwzgPCQGX/ghQgh699nI9MuB2ZVZdWw1RY6iNBfRFgaDFMFfUQqL4Y6XGO146TWdWO3qTqxyecdNDE3EnFFV4eQRA7L/HjLEf0qyg7f84cnxzrqVDzibVF3vbFDxL2+19MPptSruXWuV9BOHjki+tv+A+KS9007HQTEn/2shTV7mX6vsJSJicwX1N1HBsHJ77dcV8kMrD3YSFfc4YfoEJ5bcFQ5FGAUOK1OnF7EiZdVsFY6hXCGtFCsZSfdAgIAUXKxwfU7lXkXFHpMS4gXt31J5TfKHF3X8KT9wXpHyglWZ4xU647r3RWhMlGKi2fclvNAMEFGhDFcaT09jKeKDY9rSamdFPctmubyzg64hN/zu+mK4mQgLVnISUIDJYvwpECdgDLGCKoRj7JkrzJtIIUK7KswLCu+ZWyU5yaJ7280iYBGwCPSKwNTJn0wgqHjOpdfewqr2c04/+djyyhwnqGlWPZvzVdXVNQcffcIpP9Fq+dJrIAp4r1RLqAsXue31o4N/dt29T7y04Xe23IaKEA2HqE1y1muV9gKvjCkTP+HntLPuRt/ZorRB3t/88HOv7/bDHx1cehwSBFXBKy8++1RvHaAOgfA5ch8vrbPa2utuQD/KDYipw+p/9uVYKKvWqJN//5cLMSM2bY3/sKCc2EKEkDm2zgabbPbzX51+5ovy6qB/vaWVwscBZQT9MNcSXN5lzx/+6HfnXnJ1aX8NIdGbooXV6NTXEPL7b8HW33Fd3Fgu7rzxzzjsuJNPIyXTv/552UKm6qXXP//U4w9DRB31y9/+kdRe1152wV96S+HUnzHhHpq2tag7eusv5znXW53+4sb4MM8evOuWz3hUcB+C863NTfN7Im8W1VcyM3F9szoKSXjVbQ8+RbD/mJ/8YNcWtcc5TZ9o/ugjHBFtPc2be2+98VqM6T9zXv3qad7QV46Tpo098/jPF//zXw8rTdrQ4SOWwxuEsebz8MTr4yOVUH/GaOjwZZdDGUKaKpMerLRv3I/PBsbei5tz9nz/ELAKi/7hZWtbBCwCFgGLgEXAImARsAhYBJYUBEzqHYgDzDR3jsUTW6Ku0HdE+TPodGS8HRkfxHSsUuqKynQynhrSUJFdaXhdaVCZPNhRigtt+FOY4LRRUlCX4DPfH9hHig4VUlHxxZLjX73KIsz5TnZ21omr77HqQkA8lI6A5/QSco9I6suwBB+unCCiLa+MUFMDN14vB4h6JU1KV7pOezyW+cSLuR/G3HijIzycRHyyLp/kBIn5rh94yXi+MxlzcrKGkI7CdWS2HeRcXz4f/BeXwiDurK6mm5UcyaRJws6adErzFbafED4sIiHnfOLWOt3pHyuoHzqt0ivM8z9xmvPP6ZqU04UKIjLqLqgVII9adAyyyKSJQrkCCdAsRUSDuIYaPZX6HaWAiuVloq12k7pnhDupo/TQVdovp7fDdbwWF25XGhO9jgiFiLvS9dqRPqpCSg3ICwy/I/8M9WeoSIu5ui4rAqNJ7wmixHRv6nWj4uBWOk5/+eI/T8dQXhTUNp+mEIt8PVSypabdVm1RmJV2swhYBHpGgPz0nBm10pixJx52wJ7lwXtz1UP33H4TygAICvLir7PhJpvtfcAhPyP90+9/+fOflrZO3n0UBQTdF4f7c088+iApbCBMUGSsuta66xP8/+sZvzpeMdZWcz3qCQy5MV4+5U/nXvzMYw/dh8H0Ycf+8rftqkfQtfReq665brT6fNw7vee4R1WiODI/WxfazIr4VddYZ71ztWJ9n+03WdMEgCeO/+gDjH5/LMPomdOmTOb6LXfY+fs777HPAQSy777l+n+axl565snH6Pcvfvunvyo7VK1ix+mDfnbcSSg+LjjztJOvueux5xV75Wf8ZzaCvzvttvd+p//loisJdC+v4P0PfnToEYxT6T2isVNqIALCpT4GpQ2a1eqYK5ffqD/jurixXNx50gVRZ6gUDBed8/vflI5v+bWPP3j37ZhFs2p/xtQpkyAsemu/P2NCG4q3z9tmp+/t8fSjD94Lngf89KjjH7jzlhvw/zDn2TNWr/3n+WcY2y233/n73914teUNqdBX3Ei7hEfMPZoXPakcuA/j09PYLK6vc2bOjIi23/3l4qsaBw4crL8TQjwyJpYoNSZN+OhDUirtse9Bh76iz9czjz98v8GReYP64Y4br7miJ2x7mzfgDVlw4OHHnIjKYvvv7bkPaqDLzjvrd3c+9cq41//zwrMX/vOWeyET/3DyMZGxfH/GiH5xza3XXdmjugI/FkiL3jBb3Dy053tHwBIWdnZYBCwCFgGLgEXAImARsAhYBJZOBAg/E4gm2AxhsaF8KlbJKN4Raul9MT2URAdB6MW8jDwrnFQiFq+rSiblW1GhPYEJvg8QWEaZMbwIAyQEK+VQbBg/BuqY1fSlaH0mHcaXDmWoODikBIxA0OXkc3PjMTcZ82LiVSRfULYrxdbhC+htfKEV/UGYc7NBRywRVBSi+m7CzXny3fAyjhc0KY9S1knE5HENLSDpgktuJXEJTkz3lCW1F/MToigSC5IcFWiaGh0ZFCXHIkQfKmAPccB/UEh5eVYkpZZwnXG6ThbdEb4zVP+T2GhnokpOxzJy2uhQFqpOf4bqKHmV3uuI0nplIlKAB4m8REQedJOmSa+zul1KtzVsTCsZv6K6hceXxUVk/g2JguKmEbeNSFSB64brNOpcLT4XXKNreQJXKoy4zlXrPtV6/AYRFm3FdFAQElN1Tb3an689gTSuCYuprWhroK6DsCiYdOta1SPVSCFV1qcppCKTb5su6kv/dNgGLQLfKAQwfM7Km4LV+U88fN9dvT3ctZf+7Zytd9hlt2NPOSMK6hLofObfD99/xQVn/4EAful1EAGPK7VUb6mYSutOmTjh4zN+efShvznzb5duv+seP8BP4pdHHPSDxx+4+/byvvzl9F8ee8Ut9z/xwx8ffjSF82+/9vJLv1X6m/JUSKNGr7wK958/dw7qus9srERnwwi6/OT0qZMnceyXZ5x9wb+uufzvhqww9TAzvvi6Ox4866KroxXzmFzfceO1V1z197+eWZqWilRPmEqffek1NxvcCL7/8VfHHP6RDJ0JhhtypLwPBJaffuzBe3fZa98DKZzHwPyknx24N2m7SutLIBM7/4+nRkRIT8+KQTJEVE+eGP0Z1y868dtamvHAcnj2G67o2TPB3AOcntR8hAw6/YQjftITsVTan76OCddg3H3a2Rf+4593PvIs7yF7XpCiw7T3qFKB7X/okcdhQM8xxpF0TqUKiL7iViWmCp+FKy/8y596wo/0Y/g79ORtsbi+PvnoA/fQb4gBVA1gUK4KArffnXDkwX+68IrrNth0y21KCQvxZ+nrrrjoPM33iT3OmyFDUHeK9FvYlB71BCTlXy677tZf/fHci/AVOfKA3XeAnMFTQxm3lsevY/+dN1+vlLTs6xiRQu31l1987uF777i5534NLfbLGm5/0c9k+fVWovtlI2rbswhYBCwCFgGLgEXAImARsAh8xQgoHRRBZwgFzEdXVNlYZXcpLNb1SbNdVFa4ij7rD/6M/KYn1FenHhpYl35h5WXrP1ZKqERVOpESiYE6Y4gKaYAgLUgLhcKCILvxKyAYjakh51FiEIj+2lLLhkG3k8/O8aWeyKOcyId+PBGr8eIxuBLiIYv6ShM6gcgbL/K4KNRran4u6G560KvMZZQyqc4XO+FV5N9wg9bJCvR0iLRocSoT85x4SlYNkjbgRREGbl50CUF/vYtKXCgkFfpHc1EI14MW3cEyO6kjurVqZlRIfUCQCkPIGaRm0p5jpIJ6SzWbxLtUSreRD5qdpvx/pWrQk4oUkPdGlJophtG22hugYw0qEEfcKalHQ2GRgLAoMks8Ka/xt0hrGlSLsICUQtEBYQEpNUTnIKXoh2gsJ+3FVEcVlTIKUUZkjaF2M5KYRP4buna2rp2lKpAYLZoAWak1QsETaV50ruBp4UolUkhzZcgNusVrAkPkly64exT2vlVcRFPSbhYBi0AJApjkkoJpcaAQXF1r/Y02lSgg+cF7b7/RGxnAinSUEz2Z5fZ2D9quVP6bUq+HnurSV7wNUCxMUMqlcrLEXIN5uDL71PWUUsbUQckhW4VMT6oSjJ4JtvamOKlTPp7V1lp3g27hRkB3UfhBGIyVJ4Y8tGfKyPkdCCL6gBKFtEeP3nfnrb3hgiG6PKqHskIdcmdxY9TTefrKCvjeDIr7Oq6f596l1xDQRiVy3x03XdeX1fH4IgwassywRY1hafv9GRPaJbg+f96c2T0pgVjBv9LYVddgP0Gimp7UIF8WbqRA6kQmJGasJ4wX19e+jAtp37SYJugLiWja04KcNAbbzL2e7lGlDxjzF9IT0za8Rn58xHG/vPvm667+86knHm3m+ecdo96eC6IRxdG0SRMnmDRjfcHA1lk8ApawWDxGtoZFwCJgEbAIWAQsAhYBi4BFYIlBQGQFf8NDKkAgUFZS2UBf/DbzYvHRYUCsXIyC8hh5rksan6aqdPKjkUNrXlp+SM24EYOqZ1Wm4h6KC33PMgqNlXUJKg1SQRHMNoQFTRHwhqiA3KA+29f2PSIM84rkdytWTn/1VLq1JyWFR2IjbV355jAf5t3qxACjs/jMWOWDrJMLOqUMiDnTWl/JzGx6obsyn817bn0iF1SkO7pnxtz2ebFkezu22JIxtDi18Zl+nTejo9JpysUlbhBh0eY5fovn5CTBCPGFqESZoD2pmaqjtEsmyVYh5P9pkaJChEC7QvWtEdmhRkRsoMyYpdA9+Zeb9bqJ9yIhpuvsjGCO0xpMEWXS6nSGLdqHTpXGEi8KFDUJ7eNRW6Rroh9SwMBPiXGQvCYiHmKSYiR1zIN20YG0CoSUTMoj0gM1BvvB2keKGky7F4ysLpIfBpRNd1E5MV+vZ6reVNWbKWVGRtcpLCD2IXTymk4QEahA5quvrZHSQ8bd2pNGhWfkPIEx1BaRYkQlsKTFZ6arPWARsAhYBCwCFgGLwOdAYMCgIUPPuuiqG40PzbbrrDikNzLzczRvL/kaEbApob5GsO2tLAIWAYuARcAiYBGwCFgELAJfAgKs6SfQTJAZdcUaKquKnJDaIoiW16MocN3QlyRgbioVm6H0T3MH1VWkGmvSy0hZkVQkOyuygqBxxG0UC+F2zB0hJ4x8waSMKvWu+BIeoe9NuK48JmLVvSo6uvx2N6+YemVYp1xJpps8GHIBXxF3yRz8TicXdkYkS5vTlp7rBfEglm9JhBk1L1lAMutkkzW+lxgYz2cHOgmF1itz88NB7tT84Nj41pr47La42z2twm2bVuXNbxJ8KB5IiVSv20AWDFMhTVRcBERMoXhP5/yITkhE6ZjkuSFcPRXC9mzwLRRyNrlSXmBeHkqhEDpzdfzD2DBngjdEagVfZIYv0kKPELwvH4xZUiyIvIjICvwrlOJJBAEkRp3YBcYwq/doPpJqOofagjtooAGgW3vIBPCMqR7zaJiOQXwN1L5K7AZtRD4anlw/OCblRYX2tSg8mCNKHUVh9WWnGsqIvOgUYQGBUiFSpErtt6tum67JQ7SoHmoOiIrWYvoqFEIQFsbjAhQMxRPBY4mM4jyxO4uARcAiYBGwCFgEFovABptusfWfL776X7JqmfHkI/ffveqa66xvyYrFwrbEVrCExRI7NLZjFgGLgEXAImARsAhYBCwCFoEeESCYjALCE0kxVAHg1RQUXk3qAwWVlf5IUWZ5VihCHeYlpJhRW5maPKgu3VKVjtekZSUdj3sYKLPqnVQ9BPEJQtOeciBFe5QUpd4UX1v6p88z3omYuqxIvVQUgauHN8oL3ncqvVN7fq4Xd1Jh3EsGXfk2V1kIvEqB0ZJrbnTzCZ1JOZXxlBN6MpSItTiZpGwnsrXOvO662Oyu0bWTs+t0D4pPmDg08cEnDbGpE/JOYlqdNzMTc3ME+xsUZgerUUJypMgIfCwYH875Go68wvLYcQ/Wv0N1BnIDkqJFxyEeGkUdQGYMIf2TrvCjNFKus6qIjpluIjK9lr5CtWXU7a3hPB/GnQ+DqaqTdOrEz6REZOBlQconfCsYW9ItQQBACtSIuYAwSOBvgTGGTkSpVvSesSc1Vaeunav3EBYVqk8fR+hkHQQE5AZm35xTPZm5OwN1DEXObLVA/2bp3JQMxEpBUSGPEadOKowaKS+QetA+KaEgOCBmoGyYc5Aq3J8CeUF/OEbfffldWNIimix2swhYBCwCFgGLgEWgNwRIy3TIz0/89VEnnvoHvCYw1770xrseee+t11+xqC29CFjCYukdO9tzi4BFwCJgEbAIWAQsAhaBbxkCSvvknnnjKwR2u5XWaUY+CKvDIFxZEeUqT0YEyggcmR8op7ecmIMwnYpnG2tTk5cdVD1DHhbD0sk4AWgC6qx4px2C2SYFFMcJKhPoNimglkiyQmSEAtwys/CS6cpYvR94fghRIb8KQSLjbC+eiLvJsDrRmK+IETcPPV3j61xbTXxQeybbFsv4+SHpZGVVVbrO6ZLBtpPsdjIy4iaeH6ZmOW6qzhX/EG/vrB4Q90c01semTYnFsxMyQXVrzq2YL8ICDFuLKZTmKLhPMJ6UWigfJHXRK5wgCmmbSMVUr7A8BEcB01AUhHwpNBLUVKg/ujKmo0lRDjV6v4xa6UBdoSt8VxSICIzV3PWcic7qzryw22kPO5zpwXTng6BFZEUe6275WmSidEuQFpAS3I/xpQ8VYhMgI2qKgxqKv4IcaJVaAuUFpALeF9Rp1R7VyEAUEiIfKsX6eKqN4TeqC7gP0lLhizFM0w5vjMkqmHSjouBpSEmFl3m11BfMqVrVq9O9hpK7S3W6dZp7kmYK0oK+oDmB0ECNAWmBzwXKC7tZBCwCFgGLgEXAImARWAgB/RVXfebfr7ph82123OX8P5160o1XXXoBBMYYebJce+kFf7FwLb0IWMJi6R0723OLgEXAImARsAhYBCwCFoFvCQIQFXpUirfuSoMSbZ3ZmKQE/rS5HQ0K/Q5WYFj+hRJViLRgSykSnZTSoqYymR1Qm25abnDNdJk+VKYSkck2q9sx60YZYEy2IxJEhYi9SVqE2oISpVJakjapSRTQFp8gWiHmJvSdJpbNBb4UBl4Qc10RCa6MqFUL14tY3PWDXJvv5pvT8eqZDc6y8pGIuZluf67kFsOcXKIu8BPpICsfb9EcsaBNKajkm9HdIrdtZVzyRqS6OtODup10d9LtbMmHKYLxqBQIpKMM4P1svYMogFyoiqywseaGsCBtU8GjArwrtYeiqNDRal1ZqRYYTJ7+jgAAIABJREFUC2y6CxRHIiIbTLon0kgpR5XOFVxFVojctSuc+TLEnih7j3e8AU6NyIt5YZdIhy5lvuoQ7zLPaQnb5MaB7Tekh8gAXValDkOoJCRIiUMqKNVTxBKISGDs23RMXtpOix6oQzmkWqiv65gjQ5RdqwGTbxqCh9D0qij6dzRG5IpMwiEx1N4UzcVmfDPoqpgNnEd45rTsVep0jyE6Dm5dIkMgUzRMzjwdow9s7CPChc2SFgYJu7cIfPMQeH0KYr+CFw8/m1RQ/kUm0OuMIEOh3SwCFgGLQM8IQFZccv1dD2Mif/yh++723BOPPkjN0WNWXR0T7vfees0qLJbiyWMJi6V48GzXLQIWAYuARcAiYBGwCFgEvlUIeB3dudSIwdX1s5u6hsxp6RquFE/LxRMp1w1yYXdO0em8L/8KRZ0VTU7EQ7++Otkq0sLL+0FlVTLRreMEhPArIHgeGS+roLJAXdGu8oqi7Kx6r1OcmaAR55e4TV4VNcVl957kE9l5Gaf59WanbaVqt2r5Ko/ncTNB2K00RbNE5ryfD2MTskHF/IZEOpuOVTdWJurFVThPtGWb6roz2dHZTGbN7kxydM4NJbpIFpQq+YyTaPhE1McshdEGDpiVqV+tMr/O9MHexHl5ZVfSPSIfiCKWBaaoQPb4Crfj5wBZQa28WAFIDVQDYFsQOGio9O8n2qNkGB6lh3IVqMtJQUG7pJFirJIiDBgdmAXC+FwV17GYs4aaH6sR2t31nalqZ4LsOibq+g+UJupjf4ZSNc0VF9Ep8qBTptdK0aT69C9JeijtsyIu2ouESuRZoVInQsITkTBHdecnXOcjDL1165EiN1bC60J4VsME8QgiMTDmhsEw8wojb8ZmvPbTda04CnVb/0SMm/4RgUEdWB98MdK6Fzih/MGYex79ounik0YIirTIS2nBnexmEbAILMUIFAkK8wT8NONnBwotfh+xkdpuuor9vC/F42y7bhH4OhA4/S8XXbnmehtu8osSsoL7rrPhpptroU/41msvv/R19MPe46tBwBIWXw2utlWLgEXAImARsAhYBCwCFgGLwBdCoKiqIBAexXrntnQnWzsytXOau8dIYbGhJAVbJhLx1XyFhGUw4MajkLmy9ijYHtM6+XgsSKYSsfqY5y7rh2GV9g0KGI9UpWVUzGpW44fB94KYTKoHB2Ee5YJ8COKh9AmFREVL3kagK+ySo3ZWyhKJE+qHVcYbqhOy8CiQCECWUp6joVPafWd8e94Vn9P13WUSrY1JryLhpWtH1q79yeyW5jkzOucmvc6GmlxbdWPOHTAsSE1UCE2CCQk4wpjSS1W2SCKQTWbbhu08qWOlhky+4QkdzVYkWnIy36YfECSE8Amy+/qXQnKnwoZyosCuoLjA0QLagTElUCc2RAoIN/KDwEibawnYQW6ghMFwu140RrXCd3WRwTcG3twvFll8Y+ldIU0CxMXQiMDIOhtodCfGq533w+HOdJEV01F7SIXhhk1Oh1JITYj6rD7pf+6TRTGhPQRCjQgEljVTIimJlBbzdKxbREWT6o1XFLFBJEW9jpE2DK+KNH4YOgcJRrqnyBBe5wWk+lDwS8EDo6DUET2hKcoWBSt14UDdvUrHo/ZUpqmQJsrgxPO6kBZF3Lg2sARGhKHdLAJLDQJFsoKfA3ym+bnJ7yFIVMhKCFrS0fHepoFbakbVdtQi8L9BYP1NNt9qx+/vve8NV17yt2cef/j+0l5sutV2O0346P332tta+XvKbkspAkvil4+lFErbbYuARcAiYBGwCFgELAIWAYvA50NA5AQXksUoelEkKwhoR8HpTM6PqVR0ZPID/SAYpYDvuop+b+fFkk5XV3tkFpAQSZFKR0vfw1TCycrjok2eFYnKdGIAxIWUF0PUFuoKgtFRth4VVtqzN0GkEXqdUdsyaQ61GJ7uFOLMS9omLwS30y/0vU5SgGGEvkq2lLzH6+NOenbMHZkJ3Mb5ObdxXFs4afXasLYq7qbjXmpoVbJ+boWT6Izn6mYHbY3TMtmBdX7Kq3CrAs9NK5uS3+kkK8nO1C7qpmlYzg83a8mkZ1c7DfM6w7q5lU6ziJ1cAcMCEQHhkNW/jB1boP8AEQcIAyRHCuqLQn2+UIsVKdbyNSa+lA9eIZWTXpM6ql7nCexXq1RE7fvyuSDVEneVZYkKBt6NerWimlpXM+cjhQQ/drMiKPIRedApf4sWXTUlmBx5YBR6EOh4oe/VOjBXRw3xgLICpUhO07NddSBXEnpfp/fMpZEiK0bq4ZbR+3Tk847ptxelfhqk1wN0vE3tZURK0D6z3NW4Fe5KmqoCCpGvRqQw0dzUfRhTgpbgAhHCZ4A0MbRhaKC8CIyCmoX5bn0uIlDtZhFYwhHgZyWf8xWKhZ9xk1RmFz/vE7VHYWU3i4BFwCKwSAR22WvfA1FR/N/lF/61tCJpojbabKttb7vh6ssthEs3ApawWLrHz/beImARsAhYBCwCFgGLgEXgm4OAW+JVEZkkq0RKiGzOj3dn85W5fDBAJESV1BVhW6fTnc3l0jnl6sHHuVIRevlVhI0qibg3Pxn3JtRWpmYPrE07len4EBEWrGAn+Evgl4AxK9xL2QjZYniDXVcWB3TEJX2Uws9L6CYjZ6ee9fllD1Ha3YTqjJHFdHUiWTutK1wvH4ZrTe0KlRoqnNSYdMPaymRLviGc3ZnNd4rbmZNrrZkWZFbawvVjjTGF3+MVU5082gDFyeM1ylYUm9fQmQm3aMq6s9ryA95OSHjguXl1IowUKioE2zojVMNCUL74uoYmooEKekmzxW1IHhVGqgdaYJxm6BVBvqnRsYJpNiqERtUjjdQgHZMlt6gJcSt6DRUS06xBeTFGjayoHnUrtN+kOnPl7vGRu6rzYjjUeSz3rNqW8TcEASmaitwUAUSIAkywjb+JrweEHGAuNKibKD9aRVbM13XNYgxyIitWDNF86IlJE6VzqCgaVXes6nAdhtwdBViizcwrfLkZRNltREQF1xQInoKfSkbnwJEV2PQBLHhPujLjdQF5gTk35IXdLAIWgSUIgaKqgp+Ny6mg7vtYhd9D+Cm9X/wcz2UvzwqrrFiCxs52xSKwJCOw/AqjV26eP2/u3NkzZ5T287u777N/uqKi8qmH7797Se6/7dviEbCExeIxsjUsAhYBi4BFwCJgEbAIWAQsAl8qAkVFBW0awoA9q/JNIcBDUCciLaS8qBCbUKd0T0OklqgTAZGs6NaifoV93TDhiMSQwXbKqa1K5pcdVN1WlY53qp6Mkd26ZDyWFFlBkJtSbqJdSkgQN8YjGUPmUmlFaRBpiZFb0BGi3YvaIlD1z0Ch2pp3vXHtbnJca64mHgaxtepjzWvWx2dWVyY6qtOJJpE7785uSryZydd2Op0jt/Sd9PC8IvEZf6YC8Dkn4wVOrDJIZmPhiJxXsXo8M2xeda5petLplLm0z3gV3CUK2HXq34J5LIQCZEYQKRcKJtx0zGRoN89gUOY91xSOQ1rkF4yGqzZjEZkwX+F7FA+F1F5hpL6oV0nqypSuqCimWapUjZTe1akny+rYMDEDK7gpZ+XUHs4bUlx85E9xJuffjBQdhdsEC1I1adqppcLzULL6h5XQ3TqubFvOHJVZOjNTe0zAh6vLjWINqgQG16bE+aDA4LkJVDZxvY6T7imQ3KKcDBNh56REdgzQibTg6dZ71B9tuk6Hnc6i2gJkIFZKvS7ixZRRkZLDKi4W/bmwZy0CXxUCZR4V/D4bpLKRyvoqeNRAePJz6xOVKSr8TLF+FV/VgNh2LQLfUAS6Ojraq6qra2LxeNzP5/nd72C0/dNjfnnqJx99MO71l1987hv66N+ax7KExbdmqO2DWgQsAhYBi4BFwCJgEbAI/K8RKCMqCLyadEylBAWkQuTRoAJp0ajo7mBFuoeKgBjuB+HyUk8MbaxJxyS0cPJ55T1KalF9MunUVsb9hupUWJGKkwIKsoOAs/GhYEUr7Rp1hfHHMOREafh/ISoA8wX9XwipE3IvoTCITH+VG7fC84C7ELXu61a8LtS1YcYPg/as701sDby3O2NVs9syw95tlVtH6DRvUO+1VlUk5o8cWtPa1N6dmNMc1ueyA4eHwYDhOfmOB3k9cHqalBZdTqoi7gQJv6bbTaw3ORzYPCC/3OwVw7b5KbeTMSMIB+bgi5k1SgVUAJAYqaLxNk9QofcE8goB+1KiwrwvJTQKmBdahUDwI8KCVEuFFE14WARSIxS8IxglFBd1KkP1vl7ERpVmUaGeMmfp2DDVX0fHPtQMeTbe4LwcW9b5ID/eme5PdPJhV/QczA16hqqBOQrvI+4gUj1wrGBD4TpTtH9P5t3zVGlNvV5BJMNymnDVmhaeCKUGYUwKMkx1MXX/UOfx8WgupokqRCoZ38LYwsGlxZqleeasH5EkeGcw9B2RQXdh4/pCyqxCP81c5hyKiwU0kCUviojZnUXgK0aghKzg8wcxsabKFir8DOD3kPkZ+bZeT1TJSFXxFffKNm8RsAh8ExF49t8PP4BXxf6HHHncbddfddmI5VdY8ddnnX/p0OHLLvfrnx+yP0rhb+Jzf5ueyRIW36bRts9qEbAIWAQsAhYBi4BFwCLwtSPAdyaC+iXpnsyXKILWBJkhJfi73HhKGP8DAtMKuIfDpKwYI5+K0fKlGNXamR2h9gYPbqiIi7iQy7QC6pEkQlHxuOtJWYEaI4lcgutVzOpV2idoRCFYbkiRxWNiyArVLPAVha+Cuk8/KITF36anGgqGO5350K+IudGj9qMVeXE47TLmbm3OhRXd8nyIe25FexjzxneG6enduWXUXuX6dal5Ajk+Y15HbUdXnpwkeDZkPGV58ttGK8WRYv21ScevkhVEmHPEfbjpqvxy7WFqs9eDladmM4l713ZeIEURK4lJu8XKf1KcEFAHfxOkQ3FB//FrqBP6+FF8OjpGb9C/r9gkkYIc6dSeFYaFe4oo0L8jtU9HFEZW+orQWUPnxmgva3KVhLOyyvKadfvItXxyYg3nQm+g82zuSfU9HpELqaI6orY4l3jGLl2f4in0P/O0Q3WatX+XvQqG3utpVqzhxWXMrZmHMEVZyyp1rALSQ4eYf28WyY/PkGWRKQUERoGkkpeK0yhoSEWVUyFdFmmiUG3wvMagvOAfUsA34raK8yRqrh9zxla1CFgEvhgC/D6DqPiOCqo+fJPGqaCk4HP6ePFzaz+XXwxne7VF4FuNwO03XPOPzbbZcecTTjvzXIoB4+5brv/nw/fcftO3GpxvyMNbwuIbMpD2MSwCFgGLgEXAImARsAhYBJYMBMpUFFFAtnisdBU4ryEr8CRgT4CVYI5Z3U5wu0rXLSuyYuVYzBuZiHkoLAYpxVNjQqTEwFpl+knJy1mRYPLrZHLRYvNoZbwitqX3KgfGeFf0Nfi/ILBUqqb46qmKQrfJVCSyIsCzQpsxXe5tsE2aoJQebqpW6r+jVf7zZAwxoDsIh8/qDlaa35Wra8+HidbQWeaN5nzdvHx6fDIR627pyNZ1ZfON+XwwSLgLe3EJuRonCJYTaVHphPmUzM2nOBX14pGCMJZxMyOaUslNX3NXen7lrnFvVXpNBf+KQuAcJYLpCwE8SASC7GkRC3V6ilRETzHiZjTwvABpcVALhdhNCL7nJ+YKKAm8MrgHPhm02qVWZhQtv+kT5BfKiKRqrFJMTkW/SCFFC/Xq0+6xYVI47Oo83X2jMy2sVM2KyBcDUoA+0X5hLhT8OSAsmGs8SVaSC0ga6hKYnCxmYk2V5YVjjYihgjiGdE+us4rqNus4ptv4Wpi0U9H0KuFwIv8PdS+BF4nqJ/VgpIySFYlToQ7UBlKW6BqTZorno0/gDPaYfbtSW0RPaJUWPU8ge9Qi8EUQKFNV4FOxocryKhCkkJwowR4t+dnA59SSFV8EdHutRcAiIHVxLnfswft8b6fv77XvRptvvR3LaJ557KH7nnj4vrssPN8MBCxh8c0YR/sUFgGLgEXAImARsAhYBCwCSwACRWLChJgNIWDeE0w15swmsAphUfA2KKQP4j3nSDE0WFGdFbUfJmfnKhVxFV5VTWUiWZlOOPXVKUdqiuipuW/M8x1fEVxeq8go2e3pb/1Fh797xlBNLeA2CnHnrzoPVEk/UFWoGNVJaQ8JmpuURQDBe5MmiPcYVb9dFXebR1XFkrO7wxHzM35dZ1dONtxOTKmKhs3oDgc+NzfvbFwda2/vzlXI3Dwm8qdGuMf0XZjAf8zN17l+W11EWKSkEXAbP3S6O7plsx1UBW5mrXY3ttr97iaf7Nz93PxqpxUFABtjaWLv5jVj26CRxsMCYqFAARQ2yApUEPyHJwV1PtVcFNJBLZSKK2rdXF0gOmgZ82zST/G+Xa/BB7UEhMUnqkGqqHqF86ui++QjdU+BMnGdrdBduIOcmopjnJd0firqDaWKmpP/QNYW3ZEPB6mh6Gdr1McgIiMaeV7dErwgCsZpGr6mcwQut1dZRd0bCHkgSxBZnTvLaIquDMY6h5/FXL3OmhBmkbRYwFsgtJA6xsWvRAQU/iqk2EpnA6dRr9t0f8YrrjYhLuhDpV7zvKSQghSBQMqJuIhSWQG2JS+Ks87uLAJfDgJ8lseo4FPBz5uHVT4qfr55P4nPozXV/nLAtq1YBCwCBQQC3/cfvOvWGykWk28eApaw+OaNqX0ii4BFwCJgEbAIWAQsAhaB/z0CJuVSwXD503RPkYm2CoQEwWIC8bw3ryEv6lWGqCynGK/qh3NFVkzHQLu+OllXkYwnpQiIlBVmgz9QeqjQD1wFaJXgp7At7m99s8q1r0qL/z2qC/cAcmCiCl4NpGJCSUBwjFW9JlAPvssp0J2rTbh+tVIdVSS87qQfT/vZ7OjWXDjk9mm5/Ighuc72rlyz/EFmCEqIDgJs+C4MFTsjAkGR7+5lnEyz4vTJeXKJmOEkKlw3m/Frw0TX1nNiFbNfjK/4+Pbtr7cWx5uegitjT6E/jAuv2/UqpVJQOEQZtqSIcKO+E/Cnz6RSqSySFDwPgXbmSblR9aeIMJqR7aQ2E+73ImIE7xKIjJzae18tzNarEWqRVdAjdKxGvUJBUas7b6v3G+v4HJ3/r14/GhvtPC4SY34w38kHE5WWqUVHacmP+tIiicV87euFG/2jny16zXPOE2yT1ZUdRSp8Px5HMaQKhQRlK+niwVJaTFPdN/R+evHZS5de0waYZYvppzxyQlGBdFGgK+VFtXajdHxZtT1TbaHwgLMDR4iiTh1jTCjMD47jceGLtLBGv5/OHvvKItBnBMpUFfy+Gq2yXvEz9rH2/OzkdxxqK36e8vPPbhYBi4BFwCJgEegzAov7EtPnhmxFi4BFwCJgEbAIWAQsAhYBi4BFYIGJNsFc/tY25AREBe6iBHcIIHPOkBoEro3PAcHqgSpjVUivkc3ltbZdwWupKYaJlEiLrOiRYJDHRdHPQqoA1+0tdRLXGqKiNC3HokiLJZXQAEOMXQmMsYEjhA9ExniViSooLsAzVx13c1UxN1sZd/M1yZgnQQoqg/T8bOjPD7ys1BUEtAmyv09bwpDx2TEWiyX8vJgAZdvy20coz1B7mBjQojX/7YlYwq2Ix2Mb+Tkn/n5suYYp8QEPHdL8OMF3k5LLEFYEx+lXswLtyYigKHhBQBRwDqohU9RQ8Az0zYwUz1kIrpeqKsodSHpKsoKCA0UC/eGVq3vEpGqQmbVeY9zdojZHqfWhUXIoeberblpXDNAxlBgNKBS8Ac6zQnGWN8Tx8+grIC2mqFPzIneMQvqlAtHC1i0MUWLkRSxAtpA3KlR6qLVFUAwXYVETi0VjNVAdS4qR4FpP6osp2ufwLFGdyK2Ee6st5r+nw56x0DQwoNpQSaixhAxLhuk4RE+u6HWCMXi7/mlTnXlqjuAphAbjjOJiQTNFZCFHAqu+KI6i3VkEekCgjKxAXXWQCj4V/Cx+TYXfc/rp4Lyi0iRVhSUG7UyyCFgELAIWgX4jYAmLfkNmL7AIWAQsAhYBi4BFwCJgEbAIfIpASRooArYEYktTQBFApRTSAclAWAXSotRom+sIP0cmFMU6kBUoBzoVpB3uec4yIiyWT8S9nlIjRZ0hcqtALX/fL45gKFdWLK7+kjrcEBXDip3jmXh2cCX4TzoSSAsIC/DO6yGzikh3S5niJwWUotox+YMku/JB4rVsUmvyfYLrrMRnHAheE7zfwvNitX5RuuBna52geUzgpad2Z+MTconKXIWUFkODIL9DPucObY1VzbyqYYeWnzY9SjvRsBTHlr7SR1YaQxY0qTCWmGZzvDAH5JseXeNGKZJyKryG/Cj4WpQm9OqJoCgfyU8JjoJdOe9p2XPmRcbaMRXeBzpCqihf/eB1QRM0VD3Ylj67gVMlxuBpt9qZ4aZESFSpKyPVnDJj+eOcXPCBkxdpEyW70m1CUT35BX13I4PtjEiIFs3ldURerCgT7gZ5kjBeyrWltGd6VnUN8+6m6PpCV7FmYSwphWPF5zOPyYBGIBfIjbSuYfxzEXlSeGLGtFsvMO2uUKPk029WXcbBjA2tmHRWEBmRgbclLgrY2s0iYBAoISv4fYVCayuV76t8qALRy8bPT372Gg8fC6BFwCJgEbAIWAT6jYAlLPoNmb3AImARsAhYBCwCFgGLgEXAIlBAQGQFQU/+pja+E6Vpezg+SGWwilFVEJBGbcFx0hiZ45g0E+RhFT7EBnUUNg4rRVKMUYB1oNJCQXr0uhGzpUv9HJullawof0yCZAS8KTNU8EaI/BGKx7o+6QgqpncFY5tyXmdrGGvIBW4qH7gDPmgLBlfGszO2+DRobfwwWNmvrQQi/EH8mpjftIXGOTnfi73ndeWyackDNNbhCqq7XaubZiX/cyUdNGRUpERQISAOocFYYTjN/UQBROoQkzaK+SAVRzSvOF9IHWZ0G9QKo/Mm6L74Yf9UsWHunNXdwapdrWDQPVZtjtA9WCFd6ElcfQqcHVXW0I221vl/eTHnFT/uyLNcSp5Kx0+sJ+7nlKj2gq3rYH00iibpEBA6MU5KByiN2VJdrKdTW0gDVOuL1hCkVaozSMoKlDBzJRQKk0knls3JXNv0ojgIpQKT0vuVcDmYexvSUB10MF9Pqu1K1anVver0WSKFFZeU+p5EnhcqEBnsu4sKDOpZ1cXiZ5et8e1BgM/Nmiq7qYxSWUmFn18QFo+rkBLKJKf79qBin9QiYBGwCFgEvlQELGHxpcJpG7MIWAQsAhYBi4BFwCJgEfimIlAkJ0ofz6R9IkBa6k0BaWHIg2X0Gj8K/u6GjCCwTsAHpQUrVKMUNsVjBMgJsBO4hpxgHbsbj5I7uXJMWKxyIqrYB/xL6/Slfh+ajKqY1B8L+SywUl7nYHZ6S1PV1/Z7q2cIgGlFnCGBCLqDIYFoguktTTm/IxuEbXk/L64i5mS9eNz3M14uyOXndCeMqiJaka9Cmwv0DETVUbBEe+lYgszghNs2tiqXaG6PV00J40m3QtyV7ulu6bne+L8P3PON49a+E0+KCJfw8ShAblbysy8YXRM4L6hi2JgHzBEC5nhaMA/ADBUCz4MawxiN0z/8KZh3VXRqwYwrpaxKR7dcV4NzRoEwQe2BzoJUSZPVS4i0Wh1rVBmgHtD+aJ2v0d0h3Bqk+HlW7zt0PEfirPB5HVUSKXeVAmFWcY0TtB/gZLyCXoQkUl2Cjvabij4TtYHvrCVCgfmfEpkxUF0drYeTQYgz3vej1FmkgEpHptrShPAohmEwqaHKZ3txwCQIiZBlY9gwbScNV4PIlrgm4sCiNz2fKHDs0HWkioIkYr7Qa/NZZT5kjWG3VBd2swh8mxHgIyZi1jlEZcvoZ1BBzXa9CmQFfhU2BdS3eYbYZ7cIWAQsAl8SApaw+JKAtM1YBCwCFgGLgEXAImARsAh8cxFQoNr4TZh16gRujPcEBAUrTFkFz9/XkBEEm7kGwoIAOsFaNmPATaCWFeXsCY5Sl3oQFgTaeV1Jlqe+cRD9wr4vJIVZtN7Tovby0LcJ9hvixXhKRB7L2UDcAOB4UXD9q9ggGFg1P6eIqUm3ZYgkkQmBDLXzWrEfkC4ocEPfCeKOG2QzybSXSXTmPnGq1/hz2PnxIdmge1C7/CoUqFYlGVUEgT+g4AlSIC3Y/JzvxHPLV+ebWxOxyplzgiC3jKLijO1YRcG3CMLgjb+9sftrqt98/Fp3he52Ufg8FHFhsCqkefqUuOAZKEYxQQCd/lNnSBT0L6Q0Yg+hgd9Fjd4zh2gLU21Dgnw6Zcr1Nr2NfBC1OUFtTFArlSrLqNWVIjrFl+KH9E2uUkSFzi7cSyqJCr3/bzRffV3bqfOdSg31WDF9k3rqbhY9c3fXYU633EHiblzz3BMpoHRUvggEsQr4amyoTsflXzFAJEKV4M0rXVRL4DrjgDl6dn22UA8ZBnDBI5gXxWeEETOPayZtZNItxEWw8MFUdq/o81aX0zHmpi6BsCD1Vr2ur9aezx+KE5POpl11UMPwGcWs2xBP5ueAY0mM6CNht28wAsVUUPyc4XfTriojVfDq4XNyicpLKm3Wr+IbPAnso1kELAIWga8ZAUtYfM2A29tZBCwCFgGLgEXAImARsAgsXQiIrCBQY0ohGU+BmCB4AzFBgB7Cgo2ANKvhV1TBiJRAMGl3yJ2PJwWpoLjOKAAgOUgBNbxYlzCsSRvVF2JhSQATMmaOQImTcker2SPCghRAChi35YKwJeG5xlT8q+gvGFMYAwL9n6g8WdwzVsv4YS6rqHmsLefGu8OE5yvi7uXaFcHuWi7m5DZoiM8jB3tzvPajUJYWsuFOyxQ7Pl9D/67v+wrOx5ZZEA0vPkGYr5AD9ai839Uw2YvPSacqvIEyXXDzGX9LVvOr2t+K/SBNVelWUDYUNkgGo7worQN5YdKMMQ94D4bU5VlRAkBWsHGeYHuFZmkSijHHAAAgAElEQVQqusrYeC8IqxdrlXXkM28LM65T16O0QOVBoH5dtU2gnzvRB+gXyIzb9f5h7T8oKj2yuj/1scn2w6fUgiiOouoi37aT0xkbrDNupGiAeJGFSPRZGCOH7sh/QoqLdfSA9B7T3jeL/asQSCnNK0+pnfJwDwXVkcBQTfOBLH2WSGkByxF1prABuId3Osf0j87BYyCtibxndIh5i1k4SgvIN9JIteg9Kb44FnlpqDAWkUE370VisI9WlVvyonQU7OtvAgJFsoKPEr/PICxJBcXvv4dVnlDhc8rPJLtZBCwCFgGLgEXgS0PAEhZfGpS2IYuARcAiYBGwCFgELAIWgW8SAkUzbbMS3vgImNX7hqRACUHQleOkACJgbhZ4E9QkMMu55VWi1eIqBD5RBJi0UCgPCFybtv/XMNJvEwc2aa9M0BxywqhL+C5BYJdUTNMUBB6mB69j5bpeS1kRtkjSMFGVO9UIaYYoxmC8r89IYB48C74Kn91K49Fgim8FudQnqUAUpKSuEGmS6Zjd3ebO7q7q6AjcfC7OevvQSfhZtybelB5V+QFjmE0OfjZw421evnWVRJirjsl6uT0MEqpe6eQlFSmkhiL7EumhVPI1Yb517FQv0e17Xvs6jhtWJVKxukxnfl21t30YhHP+/vYezx+7xl1RP6W0KN9K00WVnmPlMviyZ74wt4wiw8yrQkcKc4x5WKVRg1BgbqaFWlozqlCDFoyle3kPouh+2UH8JiDasOMG+0AEXCwyL0fzU6H2MMomeJnWkedUwH6ueCCIOa4tJJua6rj+E0KlMIvyMuz2YxsIyh85H/sppZCRf4WA2U9QrhxPRGmtKmKhs7rIiX1ERgwV3O/q3CyVpMivlOp2qkNxneOzkhKBkYrzhOq/XlPCogH3gvRkunbB01HHbFGOKT0PXdPhhD7gNWIwYiJRaiFGdDihtiBqICUp4MyzMRbm82HSeEWKjKICI2rYkhflE82+X0oR4CPC52BDlU1VNla5X+VfKjOkqoCktJtFwCJgEbAIWAS+VAQsYfGlwmkbswhYBCwCFgGLgEXAImARWJoRKJIUPAJBGkgKY+BrCAUC7gQvCRATGCaQTjDHGCsXzJILKWQgL2iDlamshudaE2xmlTarUgtZ/gvbkvK3OX2kfwRjC2bPhT3PQxoQXkOyGF8OyIGpihCLHHBqFOx1xViEXb4zT0Hhj5MKQ2vlPDjwvIWV+n3fICzoh0knRd8IDhszaoMzgfK3VCaqQKBwXbTAPnD8tk7lbvqoba47K1Mxuzv0uzwttZdRtiLfuaA2Ni8ckpxGvyLlQ7xGmZFydcnAHeiF+eqO0K9o0fNkXM9LumHMFQESLd8PEN6EXiw/f62kF2+f7LjvNnjJrhXUrlJ5RYqSzRU/nyg/hreL2PX41CZdlDmptFFmM2SFISwCPZFJO8azETgnMM++kmC/9qIEIs8LyIVGvZZrw4K5XAzRF5/UBO9LyQpDtRWO4T0xDVIhuq8fpYEyhBMpolaLMCaoH3M+VL33FeYvzH1PpZC+Kub6+gwF0BU61ul05e91sm6jDLVvcN4NcoIxcIbkA8cT8TBMV6diIkZ0+21FHCyj/X2aU4+pUVRKyirmtBXlKXwGG/S6RuBAcuj/T1Ni6ZqCAkL+IGojsiqPHkkcU/Hp8bkQv1LYiqxcXIRFrU7U6t5spA/DP8MoqSDrOtUQaaPAncsYI1JGUQpETWHe+ZAXlrQoImJ3SxUCRVWFmcv8XNlcZY/ivGf+kw6On7mWrFiqRtZ21iJgEbAILD0ILClfipYexGxPLQIWAYuARcAiYBGwCFgEvskIEGw05IRZrU7A08Q2TSooUjuZlD1RKhkV40dhcn2vqmPLFYM8BNELgWXHWUUFEoM2jN/DkoQpwVgICwgK+kfwmwDwPJXxxWNgZFLkRP4RAq49G4ZzRFisoIBvWvv5uigrt/C8iAueneAWbfVnI1gG9hBBKCbY0w6EkVG1vKPXr6iwJ5hG4JhnYKz8QARFxu9ob852xvNSfQReLBPKUCEeKOORGyiNU2x00s2S1oRnzbiJ1my84c2s3z5yqsr70gjIzcJvcfzqDWKJRCqfU1YjPSy8hdbnJ8IgtXG+ZY0XvGTT815iUr3oGsgDL57wVpK993rq/ai/vbrnu79Y704T0F7k85epMFBgEBQ385I2TDopE3yHGGCsmK+kokLbwDVZoSBnCQXsQ2eESqVmaeSKErXAiC56Y05zZ+Zu4TWpoCBGcJ/gmO+M1D4ppJfXvURDFIL1KviJmBz3lToIsdepDrcJ5Y6w08nGd5UVyCPO+2G78yede0yqiV3U/nZe4CwXiUHCKK3aRpo7k/R6os7NVeu0i7MGn6NGMQ48c7VuiHqnTuOCCoMNAQXNgE1Kr5kLnCpN6baAKTSVRS5FIhrecw32F0WIDGrgDDlB26ilmIPs+cyb1F+8jtJGWdKiiJ7dLTUIlJAVzPnRKujC+CxuovKayqEqL6rYNFBLzajajloELAIWgaUPAUtYLH1jZntsEbAIWAQsAhYBi4BFwCLwJSGg6KRZXx6txlcxptgErwmKEow0fzOb9eesuCbwznmz4p09xwjwsB+lwgp0SAlWZhM4HaZCGqjBxT3BziVhM6vF6QvPGHlkF7GAaDBpmfAVIAjN8xA4BzMw4P0sqSggLiYq4DtfJwZpOXyb9tMV/DXpeSAfCOoSVKeUmnBzXzAybZtAMAQE7VKXwPlUFYLGEBYUQu8YNENWfKACmcG19IugfU6KCH9O90Q/CGJVMSffHrqpLD0PCi7NCblZiFxhgf6CxElpL9msxEczM2G2Ya4cuj9QZqRON4jXSK0xyovna8PAKzJY8Vgs5g0Js3UDcq2r/tdLz3815zS7IiuGx1Neys8Ha8uoYS/XC7sue3/fD49c5eaSpES6Yx+2EsNurjVYgr0xhjZm22CB8sE4WHSrkzIQX6AUQnGR1lkJP/6fvTcBtiy5y/zOdve31751bb23epHU3WohIVaBBrFIwIw1wBDDZocJe9DgwYEdMIE9ROAwYyMiCBzhYMbjAeMwoGVYhBAgkJDUPVp7Ue9dXVVde9Wrt971rP5+eU6+ulWqqq5equp1V57q7HvvWTO/zHPuu9+X//9npIsy9oLFSh/jtatSLWkr51FyJ12vUP9lIi8DjWWuVKaLirSOV4QE6nBG77hH2KMnUQFzcMQ8BAckjaEObBALUvshHZl58+kXvM9lpzSmVD8JQd9Zj5QOKvAacerdIfHrO3T8n6qQ7gshINXxtB3xQYm9jH+HSeGkc+tQI8og0hBFEWg8sk+5KMLC9Lp5W7ZcH9CeSo2kTIHFYFD8jdkl1DqeBepms6JlDCvk0mFEEN8YgjOWrbhp7wvGoYmQGfO4sCiba7noC9sp7nW9IHBBZAWeSz+h8ssq+PFgrP3HKn/LuF4vdXb1cAg4BBwCDoE3JwJOsHhz9qtrlUPAIeAQcAg4BBwCDgGHwMsgIHbSegJY2tYQlCrWS8L6N0CMW58JyEbIV1I8IUxAVFqRg3UIFaxnxjef7TmJtECwuJQXw+vRXxeS4VaMsee+cLsl6SFXaQPErJ2Fbmenk/YD0QAxgegG3iNaWBNosGEbZPKhdugf0pkQOWgvhC0CA+IHogcz0yF3t6nsVsHTg2va9Fg2goI6lCmNPO+p6nqIPMyuf6m6Fr9jwJJCHRExOI9tI/U3KXyW4pP+6f6BsBbub0Vh2hODPZSIUChbkp+Kc47zer6aTbOv9R+hjnU5NIv2HiYyYFgJ/OyEmO4DEipmgiCYyjNdPlOz8oYfiSJPkmSm6O+sJcs3fy2a+YYEgcEGP8jrQeDvy7P8Q6rU0cFgCC6ILq9qGU8dpagL+hZyHNLeGsKzDpwhE8GCOAhewYoyEh2PAMd+jGE8LzJIfP0rRSobS2SlkXN3BsIH9S/7HoNvRApED8SJ2KSLSnSWVJ9fMPiVfduF1DfXEloSL3qKguD4MoUaXhl6F71bBtxPeY+nz3pzYepNSEH4XsQHiV1bFKnzHTrmmD53iX7QcfM6EuHDjNsyGMJblIgwo1MZEVErESvQGIwSlVc7IWLoc3lfVOsQMLQOzFITOVN5cst/JeA8Wmd8bNhdn0l7Rsoq2sG47+iAGY0Nng+8H2o956IfrFBpTdXtq3EUkZBhoj2ccGF647ovIuutX5GJhJI3w3Wv03WsAPcRkRW/WtWB+/k3VA5xn1zHerlLOwQcAg4Bh8ANgoATLG6QjnbNdAg4BBwCDgGHgEPAIeAQOIdAFVlhSXpLy9poCZubHgKdtBcID7tUIOchwiG0+QxJCfGLOMExMFyIEjbywtK/nJdt1yKiws7ihpS9ULCwqYX4DUA7IOhJ80Q7qSPtgliG5IaYflQFMcBEKqhA0EIS21nkrEeogJwlCsKKBkRi2LRSCBbgwXUg62+pzvFiVT+uS+F67ANGt1V1OKjXz6scVqEPmPHLgnBxWgVCnFQl9BHnYFY/daTdvEKs+Ztb+/yp+uY88kdx4OVn0jQ7nWWjNA+KWphHrX7YmTwy3Off2XmUdpceDWhZhZmYH/nhaJsfDncV4WiyyKIokMmCL7kjT1XVrCMyXNqGn2kMFPdlK3d/PagvfzmcekGiRn5/VA+mlBZqh0juH9c8/uC3H//h//AL93zsNed9r8SLdEy4sGOWPkFYsH3PevBnLEKggy9tJCUZ/QiO9BXiwy6DoJV6xmM5QL2UgpQPy3vevPO8e7XvJqHFNUK936Z96hD4+sRYOqJ1iFxEcgh6M3Y4C/dRWR+/FIlU2TC4XYJA7n0x08jIU6+tTFwP1WqqUerNaMD+uFJG3S+G/3Pa/9M64KCJcDiXVs2YYevkTe1TJ6pCAgbCRbNW/eKVCOLLuJuICbOUphYGp/E4EyNiamXlyV21VPsZdaHCRMYYpLniWgwSRBETYVWBTh8cUuG+KlNzlVjbe8gm5DJRImMRGLkTL9bwvqZvJFbQddwbPKd5Dt3IpDx3zHtV/u+xTuB7AB8ZnvVryw0u6lzTMeou5hBwCDgEbjQEnGBxo/W4a69DwCHgEHAIOAQcAg6BGxiBKqoCBCBMrQcF7+06IiYgeEvT3pIUZ3a/9VIgKgDCFdoTUnaPCiIFhBf7QvmOCwXsZ691tZG3EROQ9fydT31oB5ENkPrUg8gFtkHKPaOCJwXkHPvSdvanQEwhKhBRAZFvoxesCGONuSHBObedUQ4pDW7WLBvCmnPbFFtgg8hhSXtwBTPIMK4B1pwPshcyHZEDwYJjyhntZX0hunmlrziX8Qyoio0PsC4NZtL8MD3eT73bD+e5L/Itj+VfEeVhYzLxmjv6+cT2lXRmYSpaYkxMYhsukaKQ+DAosobOo6n54ehEkXY2eEVto+hrGW0rYIBp974un0u5CPJtftZ4XPscK/LmU0Xev00bp2SI0Go0wnuVHupommQP/9uv/OAzUS20woouVyZk+vC9H+f9K1oq4YJjTNslYFzoTGF8PKprEO1QCkRlmiPqABFZChlEUIxM+qaylG4XRF9Qv3MCmFJ+6RMm2+TFQlzaoTPyvqke2WKugV9GYPr1kF5XTRSHL3EjN9fta11Da5YU7oCgxbYQySO62zshi5Cv5Wdlfj3wGsq8dY9Si02bY2NFMhSGUPZ13Gd11EEJCPQ7C+T/KW1n3DU0ABEtWorOwE+krsrzuRlJODF+FWqRtplXc74yvVMpXqhdWlF+qjbyitDBwDZAEHlBdAcjC1FL4xIBQ+cOdF7GZQIOWge2jPGBjmfMMraJwqDenMoKjPRRIvHCRF9UbfKcgGGRuOqv9BHPdsY84uuNutB+ot9+pwKAMYto/BfgIoHCRrDdqPi4djsEHAIOAYfANULACRbXCGh3GYeAQ8Ah4BBwCDgEHAIOgeuLgMQKKxzYVFA2BQh/E7MO0hBCFd8JRAnIUV4hxZm1DpEFqQVpAxG/T4XoCvYfX0yOepWLRTlcbRBoA3W16Z0gSCH9qTt1RZSgXkRBYKD6RNU+2g+BjUBhoxWYEY7YgXgAccVxVriBcOU6HEOxngJWIOF6dtb/uJgDIctMZs4NrmAMsW0FFY7hmpyTSAquw75sp86IRJyPOrIPwgv7WMFkfGa07Yfioa0fyj/y2AezZ/t3H12INy4GfiEjcEkX9Xo7S+s7Mq+2ZymZW5RgwfFEzcR+1BuE7WO9fDS3LNFCJH0xLLLWhiKt7Zd6IVKebEQkGBp5fhTX/SCdK2oLs0FtuFqk7VERDRbjQbpZ3HbUaEdTw156t5fk75GAAZZElFj+2wgsqp8lrw0p+CoFjDXBooq+oF+4jh3bYE+qKIQKMAXrZX0GwxNClDFC9BCRK3WtT9REjscfAszBnnPNa/2j2pJV4gOYlb4YhUSnTH2bG7EA4++XtK6vq07oc5k6qqZxGJu+N5YQBkbWi+CvP+itZC8p0uIFb1M+lBBQeG8lAVQQeTUZct9D9ITWMQ4/qXMdkejA+AwlFixwHn2u64wT+mwinRSZ0dIxjLFpCRasrxtBIl+LrODaJm2WZWPt67jyWEVk0DXqxnNGGNXDxNfDxLh6SLAwkR+VLgK+WyrhwvqysG5FdWKshVXKKfqJ8WzHuxm7RF9ItHAksUH96iyKrqALiTji2cKz0qSEutGWKiUWHky/qLKjaj/fkf9R5UmVNSHtRsPGtdch4BBwCDgErj0CTrC49pi7KzoEHAIOAYeAQ8Ah4BBwCFxDBKqoCutNYf0p7Cx8yKmSkC1f2Q/iCsNsiFtIT2b6M8sfYpSIBFITIVYgCly4cF6IfF4RO67lYj03uDYEKLO7mcHOe5umCqEFUu6QCqQ1wgKv1lwb0hRyF/8Izgc+RDBYccJyuDY9lI1qgHy1hDttNumYVCzJZfwkqnMhmnBuM9u8Wsd+XAvBBIxtf0DuWg8Gm46KfVkHaW2Nuo0Zc1UHrm/6VwYEaySbBACt+/ho4mOnM03RrwdFpvnwNS8P6p2ldMPWM/HWiZtaL1ofC8361/ZwIJOKblzktWGRTG0vksltRTojr4KE2IqSSS7k4R1Biue7lCDoQbJQaRgN8jw4psurjsXeUT/181TbPe/7NcUfjwcrtIDDOE7j0SGviai20RcSLuysffC1Kbjoc8ZCadRdClnge7ISKGYrgYJ19HHpKWIluBJV+hPD8xXtsU/H7dZ2RZ+YM7b1eZfKQIVrHDCyBJEURG6UMR9Ey+xVMebUVV9Sx2a43ZhmP1Ec9XblPe/esG4MR7y6eltE/81KGTWrU9ymM/2OlIKHqzRPoc5bGpPonAKP8UXEBIEQBFbUJWbMSWwgvdicmjBZx5xbi1F0qpFS9ulayijT0Ist42IGx5gmlT0WkDJKnxF/eN5Q2EL0ECIQY4xnCvWjrmy394G9T6xwgWl3hmgR/5zaMTYinJBxya55pRtsH/Cs4b684ZZKrPhONfy/UfnBMQD+td7/qYoTK264UeEa7BBwCDgEri8CTrC4vvi7qzsEHAIOAYeAQ8Ah4BBwCFwlBCqfCkviQ9RCDNqUT1zVRgnAPbLe5paHBIewR5RgFrg11oZwhMwnogLjaFJB8Xl8sZEVdt04r3mVWro2A9te26ZNMjO4qzYgnlAXyFJEAd5DQtM+BAwIVKIUrFkyZKqd9Q1pbcUGCGWuw+u4SGGoVByKhTtvbfTAeJvL2fQlMW6Nom06KdbbGeb0FZgjCNm0OWxHNLH+Gbav4IntceMRCsW4WDFeCdUQQeTRrAjeVhS1Rp5GzZVi6vaXgv1PvX36i2BhRQOdI828aDD0s2avSCZEfeeNsKZUUmLMc+kZeF0Uvnyj/SwQnSzco1vytDkR1idfEtSnPT+dCqNgf65p9zrphOp0r84PMQi2iGC0X+mCZIohzwW9DxSBQdtiRVxYMS0rxZZXt1TCBemiwLBMV1RiRh+AL33OK2mMWNdTXSBv6QN8JlYrEaNl6lgaZpcpk0KJeIUx88aUe0XriMzYriMjE2WReXuqcze1/YSO5LxJ5RBARALeGWVf5qZetHOK9FDhTgkMgaIzTnmfyQfe5iLRfed7W8NMgkbg7UgVoaGUXN/QOftByzvmzygip6vzrHhpIetvpYsaSanI9UpPyUPbDL7lKtoBIWVGnhYdNaahbYgZIbmdcOpm4YBxgYD22pt5PNqClWtKXXUHajtRIBowpk/ZjlBDaqoJoj1U77aiPXLVJ9D/8MHoaduyjrPRRTybuOcWtX44+GnJZ8SyaAnK+vkSMqxO4qIwyi57tQvPdSLnwP5V32ev9uLX+7jKv+NO1ePDKu8Zq8/P6/0fKA2UTbt2vavqru8QcAg4BBwCNxACTrC4gTrbNdUh4BBwCDgEHAIOAYfAjYJAFVVRmgGXxLc1G+aV9DV2VrMlbCHvIY/5DJnL7H0iLSgQvcyWZt3u6pV9OA+k7vhixQ/WWTPfawE7RBvEEvWCxLdigq03xCmEHKQ/7UTAQHAhwgKxwhJ1tId9OZ5t7M97Q6JXhfMTvXC5dtnzlT4I57heK3RYIcKmJbJEOucGZyJC6DfqwvE2ysN6aXBtyxPb2b+Gk76UUDFW2a9JZfgLpYG6I0trDT+Wa3bYfsupdOd/XslmHpkKl2hnGYngKylREA+UHmrFr7VO+mlHqXwkLgRJEAQ1eW+Lh46GRrTwfRkk+PVN8qpopIM0DoPOsVonXlSlUrHmJvWPxIiNRV58q86hOvuP6BqkhgJnxALaHYjQNmS19rfG4YPv/7v/kP7N/A9Ia1EcAMgFNSIQynYHijEQm02So+GPbrjQw2Kt2Va40ArECxsrwSt9zEKbO9qSqRBNhBhHfy1V8gRRE4ouMRbahJfgU2HNtA9rDe2AZO9glG32882r/D2Mf8VTKi/qM6m+0jL2Qe+qdEx6R38jYnAvKlZC6Zu2K1Jiyvu8PC2miyXvrqLvNSVeTOtHbKj0UJPSi75X0S0bhNVXJWg8LNr5iC8f9KInvWHkpX6sQtoq2lHoVdpSZZw90DGLeGJoI/f4lD639D6qlbUqnTWo3tgwXxMwKvHCDvK1XSrxIlbPKGEY+gcpsjIJFOQPM2m59ArObQkjLZMzTUKN1vV0HbxDlnRO+tikQUM/0alWTQqrKhJH200fa4WNSjLG3Yq4uGTfV/3rXi5AQGQ93wP4sBB1g5jLvX+jLdznP6byfVXDiTL5qMrvq9hnw42GiWuvQ8Ah4BBwCFxnBJxgcZ07wF3eIeAQcAg4BBwCDgGHgEPg9UVAZDCEoP0715pPE3Vgoy0g6yGo2I9oA5teiPRJEPa3q9yhYvN4Q/pDptoUL5wHkseadV/YgGv9NzZkJmQlwsOLKkQJUAdmDZOGCDEA4ok0QNasGmKZddb82qausR4YkKFm9r+KFRlsaiGiF66k08YjHtjfRljw3p7Akq5W1KDerLOpccwMdS02BZX1qLAELtvWrnMFYoWXFPVDoZ9/FVx8pYQKgzBK69NbB16y48XebbNvmfxqFvmpkQVURDTniReOzgbN08tFPDuXx22MpXeH9SQsxIoXmiJviexSQyiioogm8qQzl8X9rhcOX9CYvCmqBSL8c857i/ZfEYQQg9N6D3leZpjSe31m/YLWgQH94a8ks8FEuLKj4y+cqIVpsFJs2u8X+fFh1spHXufWMtTDO9X82NLTwx+eedkc/JV4Yfh2iRe2P6g8hC2RNowhBBTGuB0/GKPPqJ7swzW2qbmIdjY1Wk+IMf6mtH6v6oNIUddIxNuCqKQHVEgr9Y3q/AKv6j1bA1/nKk276VWTsMmfVePaXq+Y8I4UC4pSWfbuUgzKjDSiIgi929VJN8lG5HvSnvdX2cD7RO1e7xGJFzldo9GeSV7K9Rnr77DQ6NepyzYWRsQoTeN9c2/TllCSUCSBgfuhrZRRZjGhDEZJKD+83PCnO02IUaloIFbY8W4sL/Q/rmPOpfc17WC8cgQ0OI0I7qi0D0RF7tl+FYVB39hII5t2zQh1Ei3oEyMmcmkJGC6NT9l9l1sQqxBHn1d5SdEENwxmVWQF445Iwl8eA+mP9P43q3H2cvi57Q4Bh4BDwCHgELgqCFzrH1NXpRHupA4Bh4BDwCHgEHAIOAQcAjcuAlXqJwCAFIRgRXSAcIS847ONloD85jPiBamQEC2ImIC0tGbTEPzvUIHEgcyCKL8wldTlwL4iJv916C1IShuVYNMjMcMdohlfAeoN+UlUBe2F5MS02s4ghvhkdj/rrIgxHplhUy1BghpD7SsRA2jXuJihvhmnpCuKdq31lte1K2xEihU2ONZ6PJi22jpUETTjWF8yBdSFWA9/ZHbU/OjiIekDx/wknvb9eq0I2/V+0tn6dP/eLXtaLxyZqZ3l2qV44os7DlIuLePogdI8NY8URTClmfozfpCL3C7p5UL5i8o4FRly59G0DLpns1hRGfX4gI6dVmRFUyeRebQ/lef5Tu0r826R86QuYr1UFLV2mCX57HI8O1xNJ3tx0eo+3nvH5LF4145GGO+Iw41JLJ4+yoYTaX0iDYpGUBsNp4t6c0Ls/YqXDJ9s//GpJ/NMwkEQKDIi6A3/8QYr8rzcsKPPrWDBaxnxUC7cA6uqL/eKId1VSAfFAumJ0MCCL8azalPpyeDrPpImpP1qOmJalLq930pT9WJsRnsp2vCP9EmVVAOcGlIdY+69oGiK5/TaLIbeLVGuezgwBtt1nX2mWPHei09GdsCLgj3ei8Eu1W/OW5XcVCjSIlBtokySZLGoa5ZW4rEQ576w/izcK5lSQynIQsKI7h+JFDxLMOPmuaGYGlVRLdc+Rg1gJSPcqEoUq0xUakOFHWCR9skcVyltflpR40bNIAJDRReua32rVJIMxh29H8qAY6gUUohZK9pOhAqCFvc7ODa1T50q6VRDFSNYScAwzwUnXNheuOgrfkSMaYS2Gy31Ed+L+FX8pAoiKe6+HxkAACAASURBVKIdkRW/psIYc4tDwCHgEHAIOASuGwJOsLhu0LsLOwQcAg4Bh4BDwCHgEHAIvE4IWAKVV4hVCHrIVkhX+EErWLDemm/zHsECwuqkCqQ9n8nlzUxw8ppbDwWb6/9S1S1p23K5nGBxpftdFhbocS3GoDrwfchWqE/+rkeEICqCdYgRh9lHhWgQSDk+WxGA2fJEZEDSgpk1PbYztK24wOcrFisurLh4eNvmceHC7lbysueMArim5X7HT2UxHcfvvPONXeey2K1tzHNSNX3dG422ZLX6Vl+GBcOkvu2l7JZ9h4a3PHdf7SxjpzQH93NI8bY8LAS3NIVotFCk7aNZKvtsP5iVmAHLroZWpgRBJGEsn/aL2oSXN6Vn9I76frYrk1G0IgKaSgsFga9Ig2K3zrCqeqzkeVH4Yagt/uQgbexYzWemF7ON+Wo+u9jPJ+9Q/qN9TX8wEQfRNu0pBj05KVeDHXkgU+8gO66Yjg15EMiPQyR2GP5dEAafFaxP69xHJc6ckkiDkHDRRdEWphtMV/zNWvQE5C1jCuwZG4h9jCPWI+QhUpAqyvphkMYpEk70H2Nt2YgbgdoprwidwcaQcI5StChTTzEGz81qH09qZOUsegKiP9QxG73D0oUakkUa/kCRUJKS1GZ6yFdv7Qxi772KvJhQzb6ou/4Jv+UdDKZMaiWu0tC6zDuodFHz0g7iyvq7MBEWRDWYNHGVJkF7RhIsZoWjMayXaNCQSIBmgUhhBjb3YoVRie35n9aeBtaQ2zbJ7FaNanODCQFuAxN6gSk568rTNbVbC1Ej1FNIY2ikt/jrHKkEilTH0RcTRugp72cbmYOYMcLrwhl0l90zvijCgO+Au1WItuJe59l5QyxqO/fzQyqkfWL5OGNK5fdUEC/Gn7U3BCaukQ4Bh4BDwCGwvhBwgsX66g9XG4eAQ8Ah4BBwCDgEHAIOgStE4ILICmuqbfLDV8WaFkNEIlpAUPH3L+QUptk3qZgZyiqYIWMYfIsKURaQhhCpnO/loiYgd6z/xYUm3FfYmivfjcokWQHJ/YVGLYhF1pM2hvRPULuQlTbyws4cpy2kdiIlFNstycx769dgoxsMfzpW8IS4quTVWEQGQoy91jdhfmE9XlO9ikLRAv4n5bm9u2h1tvrDvky0g30rxfQDj/ce/LP7Jh+BtEOwEgFcyFA6lPdEfbNKosiJBVUyLbK6jLKVzae2OkkEBj1oWHkx2xIVlNYIYUISBccEyWmJHZvk6rwNoloke1OZpDboPG1mzedFGHaHjeZKNje3lG7Y1ssnNw38qbmB356eihYb9WBYi4PpaFjENUV3eGGj2DPK0migIINha3J7nscm71HWrM9lQeO7szx4uzccnvXz5MsSUz4l0eKTEi2uJFUUzUC4sMKVHZhWTLJjrCTJS4IcrKznCBAw1hiTpRdDpiiL3NsjChSD7YZeEQZvNxEEiBblObgPL73Y0aBa+JMS3hSZIRhWFGmxW/rNJmX2qisKAyljh7a9Tz4X9+bHvEdlxP3RYKf3mBFSQm8y2Kzx31bUxQFvKT+utdiORBIqEC9yPEaU+SnRuUdG9OOqtJd24sE9IQEDnwmlAtPzROKFqjOQShA1FOmRXCaZ0PhgvnBgrw2cqvX2NNWNYG4PE8Whu1rCBs8yxFReuedtBBQppDgUodI8Igz+5/xnzNklXpAq6qrez5ftx/W1EeEM8Yfxt6x0UC97f6yv6r+m2tyso//XsTM8off/n8pzKmuyoTB5TRdxBzsEHAIOAYeAQ+DVIuAEi1eLnDvOIeAQcAg4BBwCDgGHgEPguiBQpQPi2uWs7XMihDEtVoFotlEVlpwzaY1UIEsRKhAsECog94mygGCVF4AhsKxYYa9xuXZyfohBCFfqcjHBwtZhnCi8kLe8JFF/4cWVs2aYpvlhTcr/fL1mstRYTwGiJuzsWP7O55x8tiQzs+yZIW9TSNmc97zadFk2LRRRFdec2BwXLy4H+muuW56NZK+M6fW7vTR5h3woFKlQm5HhwW0v9G67+Q+P/+zij23/PaJumLUuYSeQohENFFkRFmlH6Xf8rX4RtZUWqq2kO/vkvC0iXgEDvuAz0+jN/HntlovozoYKzHhJZ2pladEWrBPaoLFXbBABPdXLpgZLyexcmtcb3WxiUzef3Z1GnZk0aEwFtVq9qXPWxMynGmYd6SISOnLlj1LuqChr5KtZHE3HcvXuJAoA6OfTo9gPpr16Qymp/D1+5m8Ms2G7FfbPbvnUZ5/859s+QpuKD9/78cv27VjUhe0G9o8rIYPxUqZ8KolzMCp9Y0pz6IFajvQ0rXYTuSBxQRbZuu/0fk6Vb2n7Vsk6YZRnmHgTqXEyL/xTMuIYnicPXuQukagwkmxwTIJFLKq5p6vtKVJve1GXkXXDRHnM6Lqk7OooTVSev+htD+Zkxj1jEkjNh3PesWiTN1CqqDRbkmAhaaI47Q3zBUlMiANoP6lJVnVG10LUQGjBDL2vRmCKHerOwOeijEDxFXGiiBnZoNM35zlfG5CrqIuL+V7Y7SaVVNXWNd1jrO34ZyBasJv0MFJAkb6HSBc+kzJKQ8DYbDT0Sjor+jkizRSvVXooc2oMuqtaYdR9ze/xy93X12pb5d8Aac/z/q0qn+XaWu9Zkp731QKGBrM3A4GvdvEd9a9V3j6G95f0/qDad6Xp465VV7nrOAQcAg4Bh8ANioATLG7QjnfNdgg4BBwCDgGHgEPAIfBGRKASK6yvAZSeTfFkoyog4BAimBrKDGQ+kyrJpkZidjJpnxA1mEWN0S4RFXhWcA6Tll7FRhxYmCra8ZuSvrDelguPGT+W9/YcF0Jvjq9iCy7rZ619iiTNFiRWPKEEQo8rJxEz3WmvnelO7nHOx9/5tAVymegPa6BttxnyEuJfi52Jbb0jrotYcSEoV/Pz8ENbEGaONP9k4TEJFoeUb+gWCRg1ha5sjovGdz3df9vq3yx+4D9/9+wnIOaHftTtesHUySKeWc1T8X1ZfaOMuHt+EB8p0okdYq0b8svWqJE2JEdo+pL/Aj/PtM9IQB9XZITki5T+ujkIZCMtO2l5VGxdSDdPnkm27tQE/yjNo4lR0dqc5Y2WojTkWtBXrEZNrsxJ3sj7qR+mkizSkZj14SiUlBFG6t+jq6OotbmbTdWDdHR8MOrOpaO6Uk6Fkbwtdvuj5H2hly6kRRRon6/KvDv5yGMfNH0t4eIycQHf3AMSMjKJFggV4MfYQrBArDBjf6TAkoVwUkEL2aCepf2oyETs+6fywG9KYCA6JJIZxQzvtW1HM0921NJUhtL+86Ow9qReF6URDCVkJBIvMpxBiFfResPng6epVSQ/k2lFEzR0by9p7K+arEo7JSJ0coy6kRkyiZCZUkSNdH/3vWd0d59SxQ6I9c+l/gQIH+GMRAol7ipmZHy+ICGERFULEiMClVVFYigyQw1jDNBvqxIDygRVOlYVos1z9LVY3qZqVtP1kfnKquq9UQMq4cHGDtmIifL+M9vt/U8jL+rnbVdaCRGjbvvQUbqougQLM+AEzqTezmp/oqmI3uHZR/2JphpqPfXX46OMvhj+jJc2/90NKVoQbcd3AX2IgL0WXTEmVNBF7IegjV/IUonyG3dR2/heeI/Kh8Za8e/0/uFqnLxxG+dq7hBwCDgEHAJvKgScYPGm6k7XGIeAQ8Ah4BBwCDgEHAJvTgSq9E82moJGQlxClELWQyrxCkFPQahAgCCKAhNqPCo4FuJprwqEK4uNtmC2so3OuByAlyKrIL0QPi6cD36lnWFm70qL0Gzp8hRmNvUFZ1NkRRIn2WqS5S/WwuCFei206XQOVm2ypsnMrrYiBUQlhTYze5ZrjUeQ2DqalD+vOXLhSlu8bvYrHhMF+Vfixrd4fp1xMKdIi+9JvPrK3y1835nDvb3P/8zO3zKRKGH7eJAu3TXvFVOHi6x5k5e1mXVfgwDHcDvPpUuEQx0uHSxa8rXPRq9oTjcnvZeKPArTJFvOUv9FnWuzvCrao6TRWUw23LaYbkx6xeyciHxFKIShGHoZcasr8lziRJbWinQ1zLNB4CVxMxws1KPBsgSIofwOEsNRK+JCuZeiQdaJ55Ot3TPx1tv6xeSdqd/aOFCwhZyl5xS98MOjrLH4WPcd8/dNPHK2E64yJkYSLjKJFuPOES/bMxItrNeFNWaPzkQzzRcb22ZOh1Pblv323ol8sGku601KuNgkPr4jnEi3FMpkI256sWSBgiiBiLiLdjBs14rsZrV/qhu0hlrfa2Wjk5P54KTyacVxUOtI9ZEzetqfznqn60VqRAO1Wa4dRU933iHd9SN/RdEcI2+PxIoJcz1FQOiacyLz36akXvsVUfGS7vIZRVoILRM1gUCQSvxY1BNkWX4XPWGZhJI5CmJERPMr6qIvk+6R3i8r0IU4EdxjUuO+IXNs/b8vEUNG7KV/jG5ZZuwTrdXRD+0ITwqMtgl9uFAZYn1U3uPoENZv52VT0F34EDIG4KVAxtKQOfcmtXlaoT3btJ460ddEWvEcJAqLlFYITRyCx8XoRjLmFmnP829HhcVj9Bs4AB4RFJVgAT5EsBCNYKPVXvbeuBY7VPWnrq9IbNRxfDcSVfErY/VEzPq3Kks63xtajLkW2LtrOAQcAg4Bh8C1Q8AJFtcOa3clh4BDwCHgEHAIOAQcAg6BV4FAFVVhIwag+KwxM1ESEEoUyBiIKN4jWBA1AXkIeY8YgTiBRwWCBecgmgKCGhEDknB8uVi6psoD11xnfHs5R7q8/qWWC/f/pv1KfcIPRjKnGMaZPxiJR9XU6ShUmn9tqUcBpPkgTjNFUPhHalGwrAgLRBKINqIrbNoS2gs5CREFCWojK9jPChZcH3JqnPDSRPhrnwLqMphdm02+96JQ+HtRxg9KD7hbYMsJIbxZEsB3ZHl4+vnBW46J0F8WsW8mtPtB2vXy2il5WRxX/IRm3ftlFA92FczF19T8IiA11JCJ9uLd41rcXcLLISq8UVyEwZks95fjtL5xNZuOziabNnWzSXHgzbrocBISYVaQh0XSrfnDpUY0WqwH8VLkx92aNxq2g96y0jv1ozBJ6hGuBn6RZgqlCPIsy/x0e34kPjXcnsynW+OlbONDq9lqp9+YjNKgeVOUFfcuxXNPKNLi6yKsMWuWKuIVRFuQIuq3H/8gAoxd7AR+T9u+qS8QLRhPpIj6zMS93tHaxo2xF94lTv8eDaQ7R7X6zGohk/I0a0cSJ6Kg6Eix2VYP00bLT4p6nmi0ybnDL/yRsmlJjFB6rWLnQDy6UMiyem2nBJaTipvo4QdS1KK2kI1XkvaZZh4vSrToSSLKmsKp3k6Hyi11zM/yiDbpjtihPt0YRronSNsUKkVS5k3kfckSch1Rvet6d8gIFMRhRLp/Mq8rLFa176qiNlYkZ4y4O+QO089XJPYtqKwgi6h6ShmVr+ooaVPaR9EhWl+YaK1VdWBmRCzNyJdg0NIgUAowr6M26U4+F4oFoPXqiSFRwYSQUCzQ41EYrDMpo8yb889hHoaVWME+uoavC9X0pqZB1dKqWI8R+dyYSJBZ7TtFaivzfJDReHVB81yQcHHeIhHjTbdUZD+RFd+mQjQakShrZH2VKort3Nd85/Bs5buC5+d6IfSpzx7V9ZkrTeFUtfsuHffbKu8Y69h/offPvVLx4003MFyDHAIOAYeAQ2DdIeAEi3XXJa5CDgGHgEPAIeAQcAg4BG5cBM55LhsMLIHH36yIE8x6hWSHvIf/Q4hAoOAVktAKE0RWaB61OQbRAiNtZj3fUb1u0iukz5WkcLLErfV7IJJj/Lgriaqw+1SJW0zbxskvk9GFGd/LvTg7cbYfLnaHYjiVrL4uR2Alx5+dqPfbjdqiiMdjMto+rW0cj+BijbVJV8Isb15ZR30hIiHarMeFNVI217YCxQ0pVJguEGv7IxsWmx9bfFzD6u/lhN2QaHC7yoTm798ngMDxc82PLT35yweUp+iHZ7Lf+PiPy8diYsUropOen+xQGEQg8aLsPk3tN4JFpmGqPENe3lBgRKMxShuNotb149qKn9QTJYwKev18sr+Szk6upFP1YaF9Ia+zpFBYRhb6aa8RDE5PhkuHN9ZPH6p7w24jHA0bwXCoyAplHeI/E2JgInGaFZmtqAG5Sq94W2tHj5+Ot46e7d1za9PrNvvRhqgfznpBMlDaqeB2yQQHdDUbaUPkTfRbj35QNh6lGKcxZqJtqvGTV2KNwQvx4rce/QB5xNix9hHdk3q/WRV6QNX4Dh37oIbmdikRU1lQhBqE/XqYh81a0cgHsrLQsG0ojqSTDLyWSkOGEcNaE+Yct49aLkZdQoMEitrWYdbYmo3yNCryrl+LJhSVEiVFM5XYcbxRpPOK3ui2itE8AkazmXSjDempsJaNguVsVYEukLOzhGEo6kLaiHmWIPCRDm5SsAkQ+Vq0dK/UvE3qOvagvxVBIxK7FC8CmXmf9RvSBDqK3ugpDdVA0Qk9BUY0JaWclYgB9U9oFCbcei7oOiNFdRDFsKxrNATTJm3HGFzqjXluGFEIoUjRF77EijTLzH1aq1JMGa2CfrBPP/PQqJ4Wa8JFNX7LcXfuQWlCJvDfKI9BvGioNLXPlK6zVa+kPzql19N65VlBtEUhsYK2l9ctFwQMc543mXDB9wTfBTwT+V4hOo/IEyIraDvbvkuFsfKsymEV+tNG5Y0hf93e8j2I/wZtwCT7Shba+T6VcbHip/T5j51YcSXwuX0cAg4Bh4BD4Foj4ASLa424u55DwCHgEHAIOAQcAg4Bh8DlELDRCpbQh0S1JtqIBTYaoqQKS3KeY0jxgWk2JD5iBOvYn3WQl2yHhGId57uUWGHrZn0dIIXYF+KfUpoLv7aFepPOB65xLQVMprnZZ5eH/osnlr1TizRPakxLk8FVNk83VjfNtI5MtuvPtRrRGZHFNuKD3SA8rYcFr2tkc7VtXKi4MSMpLt9fIiz9P1Fv4Huy20vjjhfWNBs/vVdD7J9q3R8Nf3j2UU7xP3zwR9Nf/8MvdsU3Kw1QcBaut+zGajgVRFrgp81c93RShPReb7iltxB4R082hsmg2a83wpV+HkbxUAEyWST2HvGBLEfqmVowHE1G3YNT4eKL09H8yalgeUlhCmkYKCRB9iUa8aSgWovmGU8blutiJdvsR/UwVk6i7qnEb077QXc6ymKvEXQ3bIhO3qEIjRNisyFpidbBiB3SmjFtZpHrnIwXm0bMeB6wfqxM5nk+KWNqAktuDcLg3bryu3Xx2xR/sDlqhvLf0KCUq0RrrtYuFAjS7yderd30YfTTNFHYgoIfag3BjG2ITk+YgVoVSvtR1iUvlnpSI/ihnilCIpzJAYn9Aj9Kw9pWwTCniIyslzdWa34y3yqSk6Ke46iZp+2Z4fHJxX6vvpJsE6W7TV7os6pbA15fwsSkWrlXfhMTumsmdbEDasO8tithldZJTyHFVnWfb9A7OVxoz7p3hK4NJ2V4rV4IZgnvUDWPeEOlj0IorJtjywgLyG1m79Md5Y1ciqlWNDHihprT1b5EQIEtaZwma+qFONHI0goNDbPg2sHDolQhyrNcgUpKPxpVMzWwmVNJC5IRemSegdskYIy0SWNBKbV8Q8zbuhr5jEO5fHXVqhlv3JcqygDs8SOhj3j28j7VNkSA21S+VQVyn+8VnqWL65DQp2+M0HglvVEJMYxNvgft8j/rzZ+obYw/tzgEHAIOAYeAQ2DdIXBFX3LrrtauQg4Bh4BDwCHgEHAIOAQcAm8aBKqoCig1MwNZxaZdsuIFJBMiBNEUVoxgdjDEjY2i2Kn3zDolesKmOrJpoTgOMhr+jmNsdpZL8X6WnIUUgrSCwGJf/na+Aq7wZbumL6JSZGXRkGnFrIjmfHWQFKeXBv7JhZ7fHyXiZpXbRkURF153KIo3TY/ryk+0m9GTUeDTdshl6gfJCOlEKigKn+0MeWuivUY238jRFIqUWOs7RUusRbhIjBg2P9b9hmhhjGfvFJn/DlHbE8J7i2wlvl8dkTU/Cq8vUtf3l73+8zK9zk9pNL2kIaV+KVZFKk8bWwCDtIZvLneCIG7mXrRjkLfqLwSz0SFtC4qFHTO10xNRmNfi2rTf8ldk5tD1I7/vNaNR3g5Wk6losTsZrpyUOfa8HC20rA26oBK5LklaE3UB2x35ad4K+vPdIt1VC5LpUP4ajaA3ociNbYGX3hTW/I7GwoYsLZZIuWYsrQs5PfiqyDky10zuV0k0Xqe1y0ZFYii1UL4rDMNtQV1Ch+ffpj3u17H7mcWPdqNxO5BG4cszogjqhdJnyYhCOa+yIkgS2T0TdtEoIhJokfypLRd5pWySfbhPhqiiRkKtJA28tkIutCaRT3eeJnldkRZBLVSMSE1X9n1lhZKwERPJEU5lXn1WsSeyuiiGg6i+FEfRmcl6/6XmatwLBtlGpXHaJOECPwvZYug5MlQViL5IJWSMvBfV2wuKtuhra0N31kY9IXjOzEjM4NlTV1jMlCIisOROFHGRaGu3aOt900tSjRwj+OReM1AIjM5hUgnl0P2Zed4owMKYZPPcmdUrwkio2xusl42PRvVg0XkaxFZoW6IxJenCayjopKHRVIpUppsqFWFtMJz/vKlELDPWzXCUFqRzKECFMA7VITDeGy0qmWReS54pPEO1SV4e5bOEdHJWqEgVaWGjtYo3eLQFQg2C9v3V6+f1iqcM6x9UuYf+UKHPSRWlyKtvsh45H+zr8wmhhe8k0kK9KNGB/rroUokVtPlfqfykCkLa8yp/orKeokauD5Luqg4Bh4BDwCGwbhFwgsW67RpXMYeAQ8AhcP0RUG5qFn5gM/PMzrL0lLvaLQ4Bh4BD4DUhMJb6CWLNihXWNNuKFvytSrGpn0jvxHtLxPMeMgZzVCIo2G5zj/PcwrOCqAoWK1aMpz25VBtsnRAFILA4FzNxbX2upO2WELekr60DpsJn1f6zInanRBRPLffj5NCpXvPAsQUlxy9IA1VsmY0wrPD6gyQdxsnZM0vZU0oD9fC+rVMHlSKKeoEBRBXFpn2yPhUmfdWNLE5c2EGVWGH71dPnQqKFEbb0Xv9PlUinIIrik2L8d3nxcL8SAol6rt+t5DgddcxGkeSYOXz9c7UNZ9+TnF3QewkWIjwlXGRZPusHTZHcYsE1jR/unNRN8mdonyhaOw/WZgdn/Hyyk8fbonzU88VGx6NG3FLCqE5todWO+v6G5tlgIlhu17z+9shLnhG5jlCAswX+BvbeWJtlX6UWKge3GW2VHqNWRUWSNPxhNygy+ReI95eVt6pFrirumUZUD2QI7m1ME+VkUuSGxoo8DUwKrHmNTYjrltaZsJHK8P4eNeedatQenWOftt0UyDhcx3B/tWDE8zTXkM67EivAJVPFk2Ev+ZypmB/tGKXFaTlhj2qRL70mkDwjVGV6ISZ/Tz3wJur5qDUx7N+iA2eHQd2f9uUXLcONlbwz6vuNQd3PlU0qCWTxYVJSSc/Q5QMl5QqmksCfkvWLmpQnkjRW00Y4NdpQOznZHsx3uoOF2nKy6ncLUjS1tRNY1BQbs1tywqwiJjZIkHhWAsZhvy4S1zfp5GgX9udt7btV+5FODnNtiOxFBdCcCqbkDfFWLw32KzvXacEkc24hJqlGfzcNhdZZ9duK1/cT7zj9KOEJPM+S6U3dhYDBsiohJNb2CQJkEFDMNgmaaggDc1bv53S9SSQw6r6mtK31exnjM7asfTJvqogMBjshFfT4mjqsqA4JFnv1eVLnPiNlhfRHx/UZH28WE22jzzxnSB1ln71m4xtFwBBxD8lvo+/26T0iNt8bCN081xFqaBv32ddVHqHd56G6fj4gonOv8l13t8qXL1a1SqxAeCNy5OeqfZ7R62+q4FtB37rFIeAQcAg4BBwC6xIBJ1isy25xlXIIOAQcAusKAX688YOIH0jMyho3aV1XFXWVcQg4BN6wCFj+jAaME/08f5hJCrkEiUh+cWYjMzMUE20+Y5AKmcbftcyURbhgX+tpYUGx0RpXChLkImQPpBavNhXUlUZYjAsV9pjjlVjBRPNlCRKriqAoDp5Y3nxqOW52lTZHERSeIiggC/uteiiL4IJc+N+QkPHiSi8+E6f5saq94LAmJFfPZpPGpUoXdaXtvBH3M/0hoYLxdY7/9X2I9i+Kfr5DokXba0/tVASAZPtkl/LyvE/0+iRk9udqc393NGyOvjueV3hMslrz8q+IAkalkEDmB3nhd1I/nGDS/Wkx4AeCTrDYqu8uFFWRjlpBL5us1/3RqrwqTiiiYrCpdmLzdLS0rV0fapDFNaWA2ioB4C4R1bGY/hdVwaauG53nMDDWaxcaNLNJ1H0R+UkcSnmRmbjo8ojd0tBXbihtTbWqWhDjIhHtjSDyJjIZNes6GyqRgqikjsbeMR37oA77Tp1kVkIF92RLTt8yElckkJh1BBP9B8H+pMqndY2ntW5exy5oPEotMaKf4iN0bV/BBb5iJqRiJF7YqXtpvS2xYkO6smUq7b9X0SHvVBjEHpysRaAHc3m3vuh3RkO/sax6jgaBgiL8aLreDto4WQfSmqJEZ8JRW2bTeRFMD6NmMw5qW7pha7HVHJ6cbfZOTYer/aJf7FW0xRYiF4wQpBRR+nyzxIYNRd/bEUx7z0iGWVRtMaVOTWxBKXO11DnbJBnMaV2iLcfUphd07BF1cRrs0BFyzpHwofRe5ki/2CK55ZT2XZAg0SXPlXSFzFsVTg2TPqp0qSAdF8+3utbTKxDR4GWFgdN6fxa8pQlt1L6KYvHkbGP6zAgQ9uFiRKtKnLjcTW0fTJh1kypKN0FDp9msj3h78KyT9CPhqhRCzXO13M2IF7ZeNurijfL8QJjAv4TviK3VfU9EHkLUH6nwXOU7BZECsYK2r8tFQkNMZAVjRuUWvX/iElEWbH9I5T+qIOaz/D1F/Y1pgQAAIABJREFU+6/b9q1L0F2lHAIOAYeAQ+CaI+AEi2sOubugQ8Ah4BB4wyHAb1vC5JmZ9vsqzL5zi0PAIeAQeK0IjEdW2IgKzgkxBqkEiQcxSroSXhEhiHKAUOJvWAgoCqQqs90hZHhO8WqjKi6s4ysRGziWelAfxApeX873wmRgUbEpOjiea5LjHkLsCRG4A01D36EZ+SkG288eWawfPdOrdQdKk68p1OWMaF+pbuTEm+UrQRAckojxlMjIQ5qdPj9KUpsOCsHCpJIZqxf+FE5UvrDXL/7ZjoVz41CZiJQ8R/ba3l/K8byuTvh2sfFKCxWIXA72yFSgrvcdLxnuPeg1Dn4q2pjvzfutKS9b3pDHh6fypDP0w+2jIJKDhKZsi1E+WWB+UPNW86gVNDRBPhbfnOWr6uOD7Wj1yWYwmJ+Jzm6Zri2/XZ4Me2p1CSWe307z4haNpEX1O8QkbsCkqFIggo2mMI0qM/6U2oNtxznFT2EcEi4QUpiYrwGc9mXcvSo9jBRL5UEYHQTKFhTo3H5Qz4oMw/qOoiN0X/kidou5qBac0Ql2aN0toWrA9TLlElKkQ6rxPNQrhPoL2ueoXg/onJ/RuH3iF+75GOT72vJbj75fUQZh6Idh9jNv/ZSpwO9+9f31H1v8e8Yx99fkwK8fi4psUemfflCRFjvyhgZ0EYQT6bDd9xSD4dd6q37z9HJt4oVe0u74UTAVpt5sI0sn5AbSkCUGLLwMMoRhGqiE00o2NZFG9ZPDRn1hdn71cHNBOdcSyQuKtlB0A5B2dCd1lDKqrUqFShF1UmmfzkqiWJQYoTRZVe1CEcSRimrq9/RMAFSjqXgDwSilUduIsIh0/6cSVZUkSvbtYXGTRtSqdJoTXh6KQlZytyTvaZ/SCLylY3jG8YwwkVF0i+rFM85657C+ZyIwuBbqmIQLxoQeGQgdps9J+WRALcWjtcVGX5TPlipAp9pHF6P+Uj8QelTIWlaOqQ1aj7gi0cykpoLgJgqB+lEY4qMqXZRJe7Veoy0qfwq8jBCf+W5g8g2YI3yDMaI37SEFFN4ua5EHIvbHkFxXb/k+IVoK0Z7vyvPSQqnN3E/vVfmzsVqzzx+rnHdfrqtWuco4BBwCDgGHgEOgQsAJFm4oOAQcAg4Bh8DLIWBmRVY/iJiJxo+58d/CL3e82+4QcAg4BNYQuCAVFM8WS8xZ0QIiCZYIEolXyDoEC97bFHWIF8wcRaCAo8O3wqb3gMR5vRboT2vyzTkv9uwbF0FsmibSxtA2yF/WHVD5W5G7Tw/jlBQvUzIabitioi3fip3dUR4ORrEXic0kJVSS5uHqIJ1M0/TFMAye7jRrxzrN6NjmmdbpLTMtm/ZpPOWTS+3xMj2OZ0WZ+mltseIT/Wc8js0WP8TH4B/E84+8uA9B+z7Rl7u8QH7F9abIQf8DXjL6filDXzoWtZ5dKmrDWpHvnSvScGc2lJG2UhNFjdZApzylU3Y15V8pd/ysr+GQaSq+hCqR8QdafvbFerT6pU44ODIR9RC2ntHo+ifJKL9Hu5PpSCmovNu1HhHgBZWRtsszYm1CvXwnSq8SsiPpfSWqldPsjXJVhFFWhI0irKl95JQqBQv4aPJMmR1pd+7XU5H1qZdxX23TiXfqfFtVhw6pqBScYXbU2CxyTctHqFCB/CR1FCmkntPrRyVSHK0EsyNal3zksQ+Ca/7he8mk5Xn/8r6/OC+dEOt+/u1/Ef982SVsWyj+Jv58FccpMj77Xr3fJFo5b/rx0mQQ1GTdvWOnl9dkQf7EUtj5/PONHfVe0LgtDaJb8yzbXqR5Rwbl5emIPpCPeRbVt3fDaKv2W46D8BtbvMUDjaVYkRnm/lQ6q7LnpQbMFD3vLUqZtE3Sg2QFYT/pHZVPxQrBG+dl/PfNM2l3BeISwoX+TavbFUchsSNQBAaSBsYmuRdL5vJ87L7lHhEqwZR/WP12XEcTq1GanCvqyptUt5iIMnwnzNayj2rqD/pbZu/Gg6CnbFjyIvF2KcJkUyVYGZNt6zxB9EUVcGEaN54+rGxsGV0hiDKlqgKCKAqM/cmEuhhyn/NxPf7mG+l47gWiPeh3BCbqxnvro5NJvEC0WI9/HxJRYSP1aBsYIk4gbr+HtqpA7DOeiTChfSYFloh/b52KFowZUlsh4Gekf1I9DfZVKija9i9M559bvkdvn7X7XbDNfXQIOAQcAg4Bh8C6QsAJFuuqO1xlHAIOAYfAukQAEoQfb6R5gDz5LD+O1mVNXaUcAg6BdYvAmLG2raMlia0oymebVxyCifWsg8wlVzfbIJogVe9SwTiVfZiZjDiAoEG5mn/fwoRCEEEiWvPvcczZRlohZpxTT0QUPpPH/y+VzmkoMeIWkX+n4jSblXihnPqyFxDrKH8KY7KtdUorI9ECT4CiOCwAntK6fhT63Y3TTfkDwBOSAn9dEoPrdvxdpGLjfK6NTrDiE2TlE/D6TByXUPG93lRrh7cqrQgH7Lr8in3vXn0R7u8mozRM41o3miyOdTbKaWGlVmia/6jRlt7Rl5GDhmij6QX9rtcaDOK6nz09Xfh/vdkLPjtXGx7cWjvVUwoovlPlgqBZ86EsTFrRbXKg9tJRtkvM8g+mo/y0nLcPi3xnZjiqC/UzsQRVu+ROrQn2oe4DFA2mxGf12mo2vTX1GxO0gribxGtMd7PJDcoPdUjHTRjzaUVW6L1mnReMVXmqmHRJc4VfNCRqaKa/xqam7qcK+dA1+orM0LUKRTT5J7TvEXHkx8StEwVyUPUrKfgynQ51M38/SLhAtLhSIpt76Esq82rLE/pr4wHVB5J5RkLPbBjGqk2xUXf5/Vu8ZP/0oLc88BpHV6P2p0+FM+Gq396riIzbwyLd1grleRERM6DWyY47S4Pp1UZnp9I3Hdg8sfjl5kK8WWmgdguHbYpDaRFtAWEv9l72H7p3R97+fMU7mze8o/KreEGJsBZ0LqINWETviwQPRBrnIvNJ+FSS4qwnKmPGRMjkel7IeEM9s6B+iP1It/pWaQU4iNwi/eqw0kYt6PglbSNdFKmzVHQJIifMs1E4I+LyHlx53nW1jmt19choVcESvh4ZHBPRDiQqFnLL6XFy0aVarRRypTG4kNKokzRnFDPjmzIZhl5No5PsUczK51kMqY+vD+OQZy3PZRAxQqpECxaTOmo9RFxU0RWMQ1IFvkOF5zbfFwgWD1SfEQRp066qjbSL9jylQrvX49+8/F1OZOEtKnwvUl/ruUH9365ChIVdflVvHlPh/nSLQ8Ah4BBwCDgE1j0CV/MH3bpvvKugQ8Ah4BBwCFwRAvwQhcjYW/3Q4UczM+rc4hBwCDgELovAmEhhyWGbXMWaV0Or2RnuEEkIFcx6Jm0HBAzH8R4iyQoAiBcIFkRV8CzimUTucY6/MGWTperGoyBeS69xPvv847rj0Rec186KhryERILsYvb5U3hW9IbJtASLQMLEaYkQg94wVR59vydjZJGlIlTFLvZHyigjdDImiOfFmSgvnhtqVr4EjTNKGTWcm5mEqNKM+vO8d19Lm260Y8eFCptf6RylWxlNm77zJdQXhUhpuTuMsodEx0bytJiREfec12yzvpMrS1SeSD+oaTjUQ69faLiaWCENjZqsJyQwtdKhN12Mism0vyBG+Mu78+Gj92Wjw1E6uRpFe/r+5iPMYF/S/fLnGgaB0i19qMg0J1+Escyxt6oOW0dDEa5FoXvACAWL2kb98JbqM+tdOopsH8y9YMSskqgOSWWFFmZy/GS538iKSN/nBbn7STGFwNfWrpMaT3xukWZIjLUxhJY4wTgbisZeVJSFSHJ/mAyzka63oOgLoojO6ELzel3RNshs7knuW8a9jQTiXsgQLXi19WPQwZz+UhV9YQeh/93mHWT414pPS7TIlL4nENFceN+i+k36hpLXfSdRRcLFXCuPvVYSb5nLVodz4eojT3o3PbYQTd4qOO5SHMPuuAg3CovpwC9qss4IZPe92S9IIuUtb/KXDrX8UV8iQUpUhRh7BAhZgZvzc29PqZIbNWVj1qSKUnou9cppXZ820c8kbmqrpbSd+7KmXvDlY2E8KbR1RZ/7Ol8qweik1nDOVbVlVMiRRKJFGG3WlSSByEMDv4s0m/d6hZ4c2cgIUAgVnNsWrqogHokbvvYDf+I+VFf1W1PviS4zCKUCQMOQWJO1VHbjHhdVVAYPXwQWM/7XVFBEL30msEYhFy3CemSOzthCxDB+KtpuPRCs2Md2278IakMiLjjvdY66gLi3QgTjkogRFsbqV1W4h76gcliFfiOyD9wRyTjuiEQPtvE8T9ZLtIXqkate1OlDVV0/oc8IfSyMA2uyzedDKn+qY2irWxwCDgGHgEPAIfCGQMAJFm+IbnKVdAg4BBwC1xUBSAZIDWvYBynoBIvr2iXu4g6B9Y3ABWmfrCBhXyGDeI7wd6jJg161BmECTwpycvPcsREYrLtJhRmy7GNmgqtAjkHAcLyNxrDAWO5tXCh5vUCz57Z592kXdaE91INnJelTDlWFXOMrIvpI3zE3SrLWaj9eWOyOegurQ5kbeytZnjVEOEuw0FRmMZEYAxiCWR4WcZIdjsLgTDLqr9605fbktru/xXvuGw9f6Wz116vNb4rzVGmh6C8FBYxBWA5YEgiJvDXv6Uvt50sUCB+Rl8WqsvWrP+VG4Ad3KifSLV5vRX4qxitBNKd4zjRO/YWV3G9N1BUw4QfdFTkxh3IxTr2d8bDYkg9Hs0V2uF2kT2/JYyWYLzpF2imSU+/ptzZ/JkkLEvJ4X1TKpSUVjSMTibN/NMz2KdpCs+b9Dar1u7SOe0YeGIZ4hXB9RmVJ1WiLcFe9TWKgodyki7o/zCNx4IQElCmGCr/ux5r5X0D+M5MfAl0iiMwRZGwhoSKU2bfIacJIRM8Xfk+nORFnxTdEsS9LlEhVj1j7ipAuhhqupDOSm7fqZlJTFYneo0McUWEmPvcm17C+B3y2s9XF2Xt5JWSsjS+bPooV/vd4L0m0YOY795CSIpmohVnj/cBVQALUiApRap/JrB8/NHjmr5bCiT84Wt/YPh3O3HHWb79bYQ0y8S72trw4mmgWnSSp3dTNlGWpU3xxl3/meckzQ3/FSyRabJF4MVINJxVlMUEaJkUbBOrCjfKceIvW1YVxIFPus8aUW1AJAcYLteDet64yjLENWreRHEvaA5yQJvDgwevjjNQEUkchMjQQPvxNuuomCRuZjLfPqi4n9bqsa5yRBpbIvAMxirRQlRym80C+m7RFBhPfm2YM6LMRg9WNNQGN0MG6tomYqFC2Q796ONYrIeNc1qhK3o15ChuLdjOq6EeevTy/eW8eUTyuTN+ce2ZzFH3GYgSMSrhgv2vqcyECH5H73aZ/yugX6s9Y/WyFE2PU1B8BQK8rOoa/bxHOEeSYqMMxeLchAuzSdoQOIp041kB6HUUM7gvuKfqE78gvq9BmRBeiSezyfr15duyze+sQcAg4BBwCDoF1j4ATLNZ9F7kKOgQcAg6B644AP+b4scePImabMVvPLQ4Bh4BD4HII2Fm3NoKCfXkPqccsVgoLhBZkC6QQhIs1ud6j95BBEP82ioLtiAE2FROUJZ/P+Q+cq5E9DoHj9fx7l2tBOpoJyCqk5KBQR+pCW0w6FBXIRNK3QBZPSoOoK7qirQiK+MzycPnome79/VFyryIsptKsCDAikEBh3HZ9HI0LpaIp8kV5HsgYob/6b37u2+Nf0Ln23HLf6xUtcg6tG+SdPCwsdmORN+gSBgBl8jfvrCBl4iRMXxf5Ea3t6x3jFIHgHpX7tCvbF2U6MhHmWdqSgcLG4eJNOsnssMjl9jzwtsgKY7vsHmaKLGoW6famVzwk8hwCFMKTsbS08sSvDdp3/Xr2i2/9T97//vUPHNDxf6hK7NG2b1V5v1Iy7W10JD3EeaAIhyZjSb7enSKXl0NW7BEXvaJBRlQCggFRErXITydbQX/DYpI2h1lNUSCqapB0NNTqeWEEEFINYd4c1KSVQIYroiJhGDJrX40+qc1nZWQwr/fy0ZDNdBmPoggEXRm6WpnLjIwQmPRSkNiMeUukgyXEtRUswBXS1+KL3GCiL1RM1FC17fzRmOocde9prfz3OvIftOc7dMRDKveod7aaHip0LxaKhAi871SN9s2k3a9NJb2/7jSHXz4abThxJpo5KP+K9/SC5rd1I2kQeVxv1OJtQZHv0we5qi8+HoXZCR27WedtS7jYKePtm8LMiA66H5VmKdP9PZBoMfJ2KknYMbXkhISLU0oThV8FdR9fStMPO9ow5K5Jjgj07EokyuaSIXyVXFiBItuNaqTIiZoiZrZ6g2IbopN8LV6UfvmsarVg/gYrz6r2CsTEnF7H6P88ZyCqIeV5FrHJpsiDvG7KK92kC0tMB1ZhbdprLbTiXG3X2jF+s1R3SU1wT+iYujoNnw2uLSGrNAqvrk9bSIlHv9v+tX4XicQL089XO11U5eNAW0iTxLMZHBh/3L+fVPkWle9VQUie1f7/o15HEh8SvUdwQ7AgOo57HdGDtKjU/dtUSCVFmj/2WdD+RozhYtdYvOCeRDyhTm9TeVTln6n8CnWplv9XrydUr/WY1mqsmu6tQ8Ah4BBwCDgEzkfg9fwB57B1CDgEHAIOgTcnAvwQg0SELLR5fd+cLXWtcgg4BF4zAmNpoGwqEoiscbEC8ghizebcRsRAhIDwgcSF9CfFEzNh2Ye0F0RdMLMVoaOcs1wWCKgL00DRhmrGvGnOhQT/eHTCKyX/bTvs39Dk7IcAI9KDSBDaxvkhaiEOTb5wMJHJ9ki+Fflyb5Qfm++2FV1xe1H4tyqzU1P2AEasEAlsks7L2Zh528c0rVkpX4rRkeef4Dns7dr7Fv/Q84+66ArTra98IcKCoyrhohxDZgQYl2Y+Ik7wplSOykVCRjHU3HbGIeMTknlFxy0oZxdjfFURGB2FJvjTXtbclfTEJhetLAg7s7nyCUmskCG3Ihv0/ekXpHV6p2a/P6Wp8hICjNjFWAolVhhC8Rff+onBb37l+78qY5MDIoIRISC/H0qTYleaFpN636o15IPdCNtKZnS75IW9GiOxUjadkVjRJTpDURHtIJCoodROyajW6qYdpYOSPiG/ikJHKkLC80nqQ8xFnKOODbRuIBUiVmv7AmVB1zlG6intJQFCkSZVZATwlMEaJs4ho3IYWyvWpJ2lBTbTzORn3CvywtzXEMYIGawDczCjSBQx9wj3uN1OxIWZlW8jLfzvM31gidnni09qpnigKIXA+3aVh3TGnarChM6IKLBdn7dL1NgTqCP3Dk9+bm9wcv7J5u6Hn6rv7i6FTfnG+LdGUa0z8uodpWLbl/tBT/s+s6mx/HwtS09IkJhTjZd1zr56fb/ON6X3TbVF5uTeTJ5KZCJ1VKr9RnpOjWTM3fHO+A3hFFTRI/apYu5aLaX0RbqoGc6hQrTFWa1ZJqJCR9FmMAAL2rpYSSBFcLMCdXZ5RWQSS3lZ8jXZcZw2kRZYU2jAnhe9wt9qpAjDoNuItnqkgPWEHi9N7Ut2p1KeKutooiqqWpYhGGNPRIKHyr3KF0QLXdhEcOCdoe0SyExKsTJgqexvrsMznDUIFqBAu3gmWsNuT8KFFXavllE3go2N1gODv1ZBpPisCkb2X1T5xyq3qZAijWf5n0p8wI+FOlN30p0hTLDd+nd8Su9JXPYdKrQBcYZoJ855XMcz3s97Rl8tEaNKC4X/Bu3i++e7VP57Fbt8TW/+DxUb8TK2yb11CDgEHAIOAYfA+kbACRbru39c7RwCDgGHwHpAgB9kkCp3qNhZaq/px0/xN2vN4uew+WFX5a1eD+11dXAIOAReGwLjURWcic8QWIgUCBGkdoL84TliZ2CzH4QRi42ygIBhRjvEEeIFs9HHlzIFy8UXzsEM39czIoxnFc9DZjNbE9yX9J6ZtwgWFNpHeyHm+MxrTzpFV0LF4OzKsHHibH/T4uroDqWG2h2EUSNXeIWI4ipdS+l2K853BGGsY09q4+qpl+CkoNDhKc8nwy6Dgdt0EQTGoizGsIT3NQupkHhVP5MeSs4DUo/0uYw0RMQwkQzFU+qFQ6KFNc5U8rQj7j5qePls28u3bCjSra1s2GFKuxwuZDhSsvUENYhu3iJjiLfqpGcU9/AlSGTG6q//wZeTX/mJB8z34S/d/+eGCP2tRz9Abv0zaVw8m4wSUrzcJRFiPwS9oi3K+pepiOpKGzUBmyzBwjQBv/BEt1I/m/C6st1Iw5ZuiFTZqoIikD6DyYXSP5k0OEo3dEifT4n+RmRYUDldjV1LMHMtA0xJYjNGTVWFh3hubLhLChwzcmFhNiIucu/y9wNCj4nQULG+DObeUEEM4Z6y6aKAyhh1s/94iihz5e/zDhR/be4NDJEP6ozfrXKXYJ7S1Wrm7gvkg5MbUpmJFkfvGh7+WjNPDjzW2veppWCipvRbb+kXtSKPprYppAHh5Hml7zq5MVlJ2sHwtHr0lJJyHS5W5BExNIT2LgkLpcgamlRQDb3bK3HjJm3f5ccSLWdkyt00Qta5mezjhL915CkxwAdip861U59IQcWzAnIcAYfrpDo0lgiQ6h9W6p7UMI4bRYov8ZVUSs4hIyORxMa7BNP1VfUNWHJVnn2ci7EF/g1VCnGXc09W5trmeaad8SspxbkxscJ8vmAxCgR3SLmfr7RWddVqTufm2VxGfJTP7yqZlLlvrBjDZsh8u471pq8lXpgIm9cr6kKiAe3+IRX+biUKgvHC9wn3yoHqugf1+qsqP6KCJ9IHVX5S5c9VPiIxgHuAhbohSns6r01jeFgfbbTdP9J7xjmiBZhj5v316rrXwuAa4YV76QdUuJ/s9xBfGj9F3at0V1VzLv9SRaYwfhCfGDM2asq05WqJL1dUObeTQ8Ah4BBwCNxQCDjB4obqbtdYh4BDwCHwqhDghx/fF5AlEIqv13eHTZ1i5yC+qsq5gxwCDoHrj4DoSitS2OgHCCs7g5YKQlZBakEa3a4CIcLMVBZe2ZeUJpCckIzkpCeFh41YqDwF1tr6MtRaOWu9uu74vtTLZkRZI2G1Di7OruciF4vagAxiFi0pOCBYOR4yDIKO1FOQYbQFEQZ60pCQMtI+cWppMHj+6NLkkTPdPUvd0UMSK94tkWKzPCuUgkdpfXBItpUtJ/ZDln1B256XYNE//MyjRU10uDG2cMtrQmDNx6I0LcfcAT+Lsu9LJrYaB3IsULqkaiyUggXjXD4N1TrtLBqbsVsUWRLUasthUJ8v0jPacGa68DaJEq+hPJHbJ9IlNOizyA90Qf9dyrs01/drG2QC8HDsBc8cCZqFxBTjSWAjQf7lfZ/oibh/VuNjIEHhCUkoG6UMvFWRDHfpmjfleX5zox1NRrVyuCqhk5eLfg6VuCfP5Awd1zUQ22KlNTQzTeXXukGt42c5Mkp/GcNsNfq0Xg9LSzlda0rxKPxhmmRDtZ6sTxkIGS2iIqkt+BLWWIMmY8wufDSfUrRANJhC0dB5iRQSOe9PagMptcCW9E2kNBroDNwrHAOOVlzkM3hDbic24oLmSbwoJzi81xtq4gOCRc8IR573LpV36gx36crKnaVPsaIjMj1DUt2Hhbdn9+jUV4Z+7eAjrdseVyKvXfV2MO0rVZYCnrYfq2/6R91RY2EhmDi0Nzn5xem0f9xvScTJdB+mIrsT7z69v1e9D+Ffg2ZX3UOTECyRALuqK6eKNJjyDki0WFa0SaI1yVrExfl3LUm0xuPEZIxu0jcxrjDPtlGtpNlSlJXxuqjUIgE96cWhkhSpLlnxkgJnDqufTqkPoMrL8wbqCmliejUdY44l1VeZig9BST4dJkYGs/XC29yI1Ef6xGMIvYvXtYchx1dPUNuM8sYp9yv731PGKVN31gRav0FyGtE2iEFEe7B+Dr8eveK/clbrbRopG1lCuqjyfqpE2dcgYPA9g9k2Qhm+Du+txgjP655Id9MUkfPf0Au9+D0qD7FOy53sr22IFzzr1+qj96mOPaltf6H3b1Eh6g+hgu+AbSpgTLSDjbz7hN6f0v7WgL64CoQ/9wnCAqI+31H/lco/VfkMddP1SoP4l1kqkYf649+B0MNoQoynq01qQ7c4BBwCDgGHgEPgWiLwepFO17LO7loOAYeAQ8AhcG0R4Mcas9P4Qc0PGNJivOJlLKqC7x6IS87Lj1ezaLudLZ0r2sKJGK8YYXeAQ+DaIQDHayIBSv7cpkmyYgXrrDBgZ1NbUh9in/cQLCzQbOwLaUSucIim3SpEYfCcuFwUxcUabLm0C8UI85hR4dlCuTD6gnUmjU1VF8vNWbGD7URTMOMdEsfMWq7qOO5dAUEGWWVmj4vxXTy50F96/MB84+Rif+tyL35AARXvUj6efcq+s5jnqWZF+1sq8leYioVMU6V08UlL8mSeZ6d+7afftZYf/6UXn7hYm926V4jABebbFRUfVH1uXioRQyqDL1GCjjHCRBVt4YuSLscR44V9EnJI9f1wuOzXVhpeprz+RV/M/VSoqBhfh9V1ehlOxHU/WK55/jZ5XL9dHRuOdPssK7Bh6AcH92T904fC9kDCxRpJ+ssHvP7/sv+nXpBnBWPCz9LsOY2hO1XpfarkHfEg26f7cJMI9Y3yoGgrwsKQvho7fpGk9VHeDGK/HeWptINiKlmIN51NsmBeU+MZpyd0Dr6Hl/FTkDCSiIXm3qhDfEM265JlBqgxrcwAZgULq1Ocu2OIQzG/MZWGSE1Vaii8G5S2ilXmyVGaR8c6bztDXpGEQuoz1bWlrFLtUdEuuulktxkOFrbUjxM1YGbgS7wws/MlXPB3As+OZ/S3g1JzGVPkU6rtWSk0+7T3tK47rVYQ8bRRPTcrj4rNt3tHvnYmmTr9YrDtkTRq3JN74Yaw3WqNgtb+xdzfn3jRZOJHz8iI+9mt/uLZYNZbEPl/WhEoC0J1oHOAbNjdAAAgAElEQVTuVr0x5A4lGLQ1ChrqVlmT6Hk1UCqkwusUXW9Z2/p6OqxIvFiQ8LGqep3/N02h5pMHjrXlkwpDbUQeqZLmeYgvyJTOP6VPI63rqyyrmCgGPyLaR626VZEY9wlmyaj5kkYnTiYvKFEZEo16Dj8S7Q7ufbWj9LQQ5lW6KCsSYySOmMCF6beAnFF8tiqueXNONDH3h9Eqyn2MnkGWMTM+zVaTLqquMtTKEJ8Ure1oHwSMVV2nrWNJXcXu9COEOMS7FbpNVFNl1u29EuFCxDvjF/GBcU17IPKpLiLw/6mC6GyWKqXSY3oLwf9vVN6nwpi5XwVB7PdU/icV/ga2IgeH8nzH8J7nAILIe1QeVOF7je8Jvsc4B+fienxXkJ7pYdWP/jhPwnodRIxdOiffm9+q8rsq/4xKakEouegyFknB9yzCC/XH0wOc+H7jeYOguJYO7lLncusdAg4Bh4BDwCFwNRBwgsXVQNWd0yHgEHAIvLkQ4AckoeX8yOIH76sSE0j5JGKBH238mIQY7Nk0UJVY8YNax8yuJX3+I67n0kS9uQaSa82bEoFyRnVJyEDeQDTZaAi2kdKJWZtsgzhiOawCyQ+5Q1QF27j3Sa1xqwqihhUVXg1oluAfj5KAIOK5Y01gL/wbmG0QM8ygvjC6gmMhbjD+/awKhqy0k3pSINzwGuCc7IeoC1HUFSmHYNFcHSS74iS/Qz4VDyrrzr40iTnnCTG3XJdokioVlKFzD+kjosgZ0VqXJJxeDTDumIsgYOhWlVpd9K6GnYh+s9e5aAv6uhQsEC/KaAxDqKrQf5VXi3o3z5UxR1y77y8rd9CCXlvSMWRyrdw5YrPDIExkhLDcLvLJdhh1wix+W+wH8yMJHZxcF7UpZDi35YsTEfRr37si7Z/XjhD0XzDRC/JwSAY5JsDv1njbo9ehIjB6kgAiOUVvH2adiV4ws1mKiqa+T6bFIHgqnw4xHT6tsYbA1pQiwcx7P4uLsxIOprWe6KZOWFcKK03SVxyQESxMFAUVs+T1xQYUxLdqawUOiRU1ikh+UswYwULT/sWJK/wii2a6xfTGUd5op3nAvTkn0WJumE82VrOpgUSd5/v5xOG9zecgn20KoaEwACcj6vj3fvy0UkT9g94/px75igrE69uEy91q0zYEE/2b0VPq/jDM73/36Kmnt8WLT3zBu/NLo87E/UUt3NFTb7XrE4Kmvn0xmHj76Wj6hfetfvUFxan4/ox3POx48xIiHlcUw51KAbVPd+Wkzr9fkOxSc4WXRJlM93FfJSeWRcR8TTPvOyJ9M++gRsGSrn8uKRSxCVYKLcUA/pnoB2QxA2ugZ2fo7dUIY80xFZ4/Xe2DgISQKzlAaaNiXaujgIuOKrtd+96iUfwZva5KLEhNWikiWhA9FMxjBAGwM6mYVMC8qe41ES7aty1RoaV9jQ+7BKfKSuObOhrJDk8PxeGUu+iuCU0ojtYZAUPn07kmqK12oE0z+ryB0+o6M0JgXvVh/EH+s1Cf0kK9rBfRAkb/qNZ9UyUusYKxi+BtUz8xdviuQYDg2U311gSDKl3SIRH4P6f196n8vgqeFSw/qwKJj5MKx5u2VgKDFcDndezHtfovVfg+4Lvs/SrfqcKYp30c/89V/i+Vj6rwHbE2hqtrvaoXokV0/UeqazNGeFbFF0sDpf3YBsZ8zyFSEE2C5wVRISyIMM+q0C8IF3wndl8HQeVVtc0d5BBwCDgEHAI3NgJOsLix+9+13iHgEHgTICByn2c5P9D4gXdWJP95M7dehyZy/r0q/OjjBxY/dCDnLrmMRVPYfTgHx0HsIVSs1VH78gPqv1BhRhgz7A6pQD5Aar7sMjU9AyHqrSwv8QPrqi/Ts3MblhcXbCqbq349dwGHwHpDwEZV6NXk3leBPLOeDvYz9zv3JvtAFkHk8Bxg5iZpNhAsyA1PWg1LMPEeUdQKH5bSu1IIrCjBs4Brci67jAsW5+aCnyOFeTZBztiIEI5jP+rLTHSeeRBo+6r6WkKHWai0GTGG5yPPMJPKhtckzbuL3WE0jFM5G2eJmLoojEQCl7Q0GBgCTF4W4slT6sD5HhW2kEan+ytLTrAY68TX8+2aAfefqIuZ7290CBNKUApeZQSBLTZVDbqCJVZNKijtkWqdUiMVkQ5MEwVaKBfQSuIVhEkouiKfFXM7nZS5fZQeKdo8zLNGrPO3/MwQz40ijxu+7J/lrazPlGpOeznbXhEXJrKA8fLhe2cGIuwZF3iaBHmWy5gd8cv7ig6a0WkDpWJqriaTM0dG+/fOx5u/re/VNssmRUcHSZ5t6j7afegbD0z9w0utsM85Z3UM96q8wosFXXlJ51nS+ebyNG9qXVOITNcbsreooqokiEiUkDRjAQI/8x84nmODSwirUa7ajrJ6QxEUtaRoNheyjVvTNNK9XvSW07l36LCsEQy9XjaxS54btZVsbj7O67e+NNj/wrHh3qOT0dLZbfUjJzZGx7knrVgUkzJKokV85B82ntjZn+ceOq5qQNwyy/5dqs99ehqEVUyCF6XZzTcVp71er/Hs4/VbD/eL9rTo+YkRTiO+3wkbjQeGab3/Z1MP+h9YeQQiuKZ/dSEU60kXyVz7hKDs5aveLRIpvkXb3iE9alIYqTeEgYh8OZ9MBKlm2a+KmO+J/A68rt/2jiid02G/EyxKObr4xA9kDGuHbQc7cktinmXM1sengr+ZECHwwaALSLWl4aZJHoHI8dAbNd4v0eDbyyi34X8tdWRFHheRxo+2aR0RbniPMPY6avWytDQM1PEfCRRf09a6WcXaRGpnI2jqvTAw4XPEhNTVVlJIIUwEXqhixquiTEbCg1RY+KCE5pyJ189j/c2HqXhdkR2KEMkSb6jzb9JxTRP1kQmbsk58ZzBgIPh53vI8pn21KtIiU6TFZf++rTwmOBdkPM9qhD3EAcY3z/FTl/Jz0Pqhjv+S9sG4+hdVfqHqAqIXiLL4bzmfTSdlu4fXah1jb6BzkCKKULg/VGEM8r1GX9B/v6RCFAfiB5EXCB0Yda+JWa9SHODvZSYG/HcqCA2/oHPyd6q9RRFO6O/9Km9TAWPSqDFRyAjm1cLvCCJOEHb4DuI7zy0OAYeAQ8Ah4BC4Lgg4weK6wO4u6hBwCDgEXlcE+BEC4Uf+3GUJABj+nScKvMarcX5mh22vzkPYOeHxV7pwPD+IViVUnJdLtxIrCJvnB5xNsQFhyA/VK1p+43f+/R+ORsPhL/7sj2GYeFWXu+592wN/8Od//6UP//SHfuizf/3JP72qF3MndwisMwQqoQJCiXvVettYoYJXRAJIE4gnCDZjxFqtZ9apnd3J/Q2htEeFiAoEUbYjatjF5rO3BJWdcY44cCkhg30NqatyKWKrmg1v6sJ5bOoqPtMGG13B8ZA6kFzkOYeM4jN1pA7WjNiSpxA77GMjODhvPL88yBdWR0lvmPYVYSFz4yImsXy1KA2LHAkqglJvyev+BZGmjyNYFFm2eOjpr2O++7qr0GM43/Bvhz86VzQ/Kv0pNSoSAQCMAbHxla+F4eFFQZdj6/xCxIVZh3ChvEZeIH/soD8KwkWx/yd0toWGl94kNUNGx4oX8AMMjqdSJd0pp7pHRvHo+WFtxYskanjTWhOnirjQ5gtnm5uBg2m40kThc2HrBLlLeeZ3n/5gkCReTYLC9MH+zRu+tvLO25eLLW/JIg3ZVNXEa9ufyB7vPrh0W+eJk82wH2l82Zn2SuHj91Sd8rtYhLPSS2m4FjWtT7Mkb8nwO1QlNBO/iALWooGU0RTUBcnCKBZmg9honhlZXlP4SKs58lrtUd5qD/LWZD+ZmOvmkzsLPwwVBTIYFXV8FeQB3pCXeH1TWtTreRB1FSRye1LU71pJpw6rKicHWevIyWD7CzPR2fltjaNnIz/hvutLtIg1bR3b7bM/Mf+3KxuylWO6k49rDZ4FfdH0iKOz6qmaWtdo5fH+29JjUd6PTj9b2/mcvCt2S0CajrQo9mOTtJj3zEfTo0+373vhzvjI8Z3pWVIWpRIdiBPx/TmlnjrhvVAseiuSbSHId6ipk/nQm8GIOgyN7NDS9Vth5nE+Yhh0fckduXwu2prBjgxBPIJ9mtlYAvvZJq8rE+2RMgpRlOdLGW2CR0Q5YkuT7kLksq9xQPyFhIPiczq3XN0LJZOSPpPFD3uDYtX4YeD7gb9EU/WQ5IBMYeoyEU7o+dY0UW+bNTAxOqlJgOmobNA5Wzo6DWraR+sQmMxY4Vxlxw9N+iqeoYgfWqdUWj1FgCxJ4hsojVVHN0gqYaMXlOm1BLm8NDKlq0pkch6rr8ond1/n4rlqn8Fl2jW1XcKFJfbZVowLGFWKo5u0/p0qEPN8/0DkE/X2VyoPq/CMvuRSiRkv6Vz/Sjv9tspvqkDsgz0+bvzdZ3vqcqdin4MqEP+YeO9R+YDKf6mCXwb1w8j7n6gg4LMPERqvNv2SNVhnnN+i8r+p8FuA7y8WIigeVVGss/ftKkwKIgIE0ZwFcQOB4v9RIcWVjQCpNrsXh4BDwCHgEHAIXHsEnGBx7TF3V3QIOAQcAq83ApZE40cVYfD84PldiQHPSSC4kh9WL1cffj7zw8susY2gGE/ZpHWGXNE6m46F/SEvETr40cSs47VF+3PePSo/oDKvwnHPqXxa57iiCAZml973wDvf/bef/E+E2F/15e633s8PVi+JR27W81VH211gnSLA347/P3tvAm5HVpb717DHM5+TeU466aQzpyfoBrRBbFAvIMJFeUBRbETlwXsVvYLD9TrbXhFBRblcFP8CKhekGQSZoaEZekx3p9Np0klnnnPms+ca/u9vVa2TnZOT5GTqga46Wdl71161aq2v1lq1633X970AVFbrwYaDsoQFRAXgDkQlIApzEHkY3xCrACqE2GBeABhjP8eQ364Gndp0G66JvNZTYzrSwqxGV2Il69SwTuS3niD2969lDnhlrrIEC+ez3hWsgt2blgdYaD0ueAXEZN4jP3MYbSWPCXEyNF53dx8eLYm0aE3UWg2F6KklMeUnq54AjhhBwgQCeTnXXUqPKsfRSmWsfmQ/U6I54Jwri2052eslWMAKs5zqhwYUTUvkdXrS4hTphV5xKA+LeiX2h7SKHOC24EZxseCEi4XHS+NA/FSifyGE2ZfIQU7Ly3M9w25uad31i9KzaBZYxg6onBBo9CkA1woEBWSF3pt+o/ftxJyp61vWGhKD+9Px0r+9TxxIscMpdTSdDh0yrluwG6l4Nz8SzBqdm2hDUBbHAo/bMch4RAgalwPuxcYzUtXqkUYGpGSH67k9nu+VRVqAjocCnK2ehyUCTaFQF2NBf/9Y2D+7EnXNakbFrlrYuaAWlBeZ1fxeTuGhtLA/bhGuSO8lZ+G24mKu6eS84Y56UJor8mWp6gyxeVLkxdBQMPdI4OTvL3jNR+YVDtkV9ID4RhHiw7NfzKlPPLf62IlrK7t25uPgcS+Mf1yVeYH2L9arD2nR6dWvvr6xc9XiyvGRu7rWjx0vKlqR7/c3alBL/pyaV7xpV8eiJ46WZ3/upaP3PzovGOY6YBsIipq3UCHfBpyvxCMiCRrOBoWLWityYI1CHS3yC7KfrrK5QCIQ8LyQjeZHUll348iX98VBlTKisFE1zaTSXDfg/+mj3H5OrjLXqd+QIMlvKUPUKBEuypK72IC24z3RgFxQ+KpAnyJXS0YKPyG6ZEQlBGLJatordRGd34lRhZf+hl7n6t0adcur1ROWqdRZ6VTF3LZShMKAOy6yRH4aak9eXhZFkQ0tJfpoQcfR30VJmHqhwVHUpfXV7nEFOsN27PVF/ckXwzksk6BvgUB3FNadQ25VvzMDhYtq6dvIkDJ4BeDJZsOv0Wbr6WuIZhEYxvMoJS6wA6HR0EJCR4Jjv57a6ct6HZ/OO8LU68yNciE7CBP1WiUWBBFiijF52m/ZqYdO8ZCgnHERIHhc4PXzT0p4WXAf5PMtSoQwe73SN5T+VXmpM+eyJL0NQXWWqhoPj1DHfVAZ8AaBhOB54FVK3FMgRiAq6Le2rxDyyixuUvqq0t1KtBfvDHv/M+e7SI+Ps9Y1+yKzQGaBzAKZBTILzNQCGWExU0tl+TILZBbILPA0tQAEgcB/HoZ4UOOhnpVbv6b0Se3/kr63MbEvtgU8Nk+KY+v9gilERTtw2P6eB2uAQ9zjeSiKU6LDAi6sAvsdJTw2WIVGKBTc43mIm9G2cvXa9R2dnV3btt7Hw9YV365eu4EHYWf7Qw+wAi3bMgs8ayyQelcAdgBqtmtUMJ5tyDer6cCKXxLEBeCODd/C/LRZyZIb2A8wlLnCgqVWkJQ8lM1nVo9TBmAoJAFAFuDL1I3vJwHTti8t8Ew9LaFg620JGDt3WcFR6s1xfMajjHIBggFwma8A4ADSmNsgKKynhgXX4u17h/I7D454Y5WmL7ICEGm9Up/ICVs1QvokQtthMCYgm7lyWOF8hpuN+tihXduDseHj7QTwNE3Odl0mC+BPIDhPDgSnPCzoE6T2te8Cg6WgDfFkxLi57nhZoG1BCbE8LNx6y3WrBb0qbk9ejgYtrSwf1/uiJ5RfOhemyrwm7jXxfLk5jAa5fNz0tQA/dhe4rea4Op9Ww7uQCif0WhJBwXtLlnNf5731GDKeHimJYYp3mlX6+j4naB5UcLK6/Bck6BzL8cMpKuxS1zv33+79j6Vvp4xA+2rqf5aIpGz6NGOyrv1UWHosJgScynH26313FMSz1VcVzUrEQ6ygSIgqe25R4uBSIM/l6nFnx3jU13+iNWt5NeiQhkaxO3RynXJy6IxzeemRqzhCSZktL7uoCWIn4nzRw8cFJLskR5PYRwfEnR/EpX43Dhqy4FWRV5w7HM5ZHjX97T3+8Lau3DhjlDpTDwMS391xTbCnOP/kC8cf+u6s1lhNIhq7pJ5xvSzzHLUM8hSnDmcgHJ+1obbXfcjNVU64fQqB5ZaliS1ayV9c7Cn9VLVZmvXR8Pmffl5tx103NHYzF2EX0ycU4KslePhBzQLH5XmwQ9d6rltzFkUtZ4UIgHW6hgvk3AJ9QVsRt54tYH6TPDGWC/AfcQu6tmWF8+pyjsn3Aq+D0zdLlyXhmphTJV5uiFXaikcFHhq2Pswx/ObCywJCdUR2FAVg6IuCzrVYtGwffdftNaA+ehsj0r9Apr1PPXiZ8uHptkBkxjzVlXMxu891mzpSV0xXmcBY6uWT3EqRa8XVx3FMXh54bPRMzsJqj0iLHpWBLgZ/ngkPpVBTKhlpFzx8PK/gzFf95shmgyoGCsbVd6uVd1Cky7DCbw1r70mdBo8Z7gG0n75rQhaJuHBO3Hl74eQP/HqHCLAndGUJ7WT7MdcKHYYLJX3p95AeCHVjWxuWbcpFOv/HFPTn+AOp9waEAQuMFitBiLDhiQxB8qdKv630eSXuN7R3JhskzR8osSCANnNfxUbcLyEu6D+QFNxn0EiCHGcx0XHV7zTv55mcLMuTWSCzQGaBzAKZBa60BTLC4kpbOCs/s0BmgcwCT4IFRCAMiQz4W50Kl3MeVngg4WFlvfbv0PeX4hFgQ1PYlkwlQEz4iCneHDx283DGA1T7KlX2s7IaQcJrlFYoGXFaJdzVWQk2Y6+Q9VuuZ2Wa88iD9z4phMXqdRs3Hzqwb4/kMgADsi2zwPe9BYhYpEbaUE78brQhoGycfWsDVh4DuACm2dBQeFBYsoJ9xBRnBajdGOuWMLBAo1klrdS+st2SC+1hok5BeafKm+pVYfNYoMmSHO3gjA27Qx7mIQCdvUoQKbTFxD1P68PcB3hEPr7nsyUs2sGw6JvbDrsPPH7CkWcFtQMoApiCsOiNE8DaeJPIvpK1CAGFmfsIPTUk4HZibPhE44nt98UPfpsoIdl2pS1Qf7WRQjKbQH/rHGDh4+TaJqC8AGJFcwLE50ISuT/xmLBha6KG6zbqjjehuEklRRAqaon7RNN1jgpbLip+Dn0hlxZIqcJz4wEh2fOE0UqYWfrckdvhBk3xHr4Aaa1pj6MenceI3072N0I30RcTEgHoPQlRhqaG9ZgodISCgoecVmO37tCHnFxuhUgCX6GvusTKLBxszdv9q5s/aVawv/P+l7cUDYn20Q57Tzb1lBEgMkbVR/modfki60RwSDuD9fsA6YSAIg/jfaDaKs0eaQ30j4b9cyai3oXVoGuFPCMksuyKvCGQVBLjCL8iCXA0/EjmQtBbUYt8N6yHcbkchrky+hkSQ5A3hCfPCzFJcV62k7S0E3YHfkexGkazW63CotGgt39WeGL73OLRoZRYrag+EI2V435f+P/6bhl5yfj9313ZOLwf0kIweUWkwgsEiuNRkM/nQmepc3Kg0iy78nCZGPa7dYn9cqHoFXNFf3WtGpRDP9e8u2vd491O4/CaxkHmDztHBQLaj4syqEnjAm8PPxpyctFeERJ154W6GptbgbNcqHyP/A0KIkiw32x5WMxGy0G9Z1Cg/GxZfHbcod9tBTndIM5NuCird53MwAkZm3QcwkMxlzGnUhOuWRIiKjL7uX4QqkP6jG5FUd90691K5RkwFFdkxKVn6/1hldmSlQG156vksi5FSSUWTLCzxGeN8zkiLZj9IUi4KyQ+IclIUdywtOcpv76L1FMIEUX0u0STgzIgNKgvvh05Z46RHdc3RmpeIaa8nLQxSiIoKEv9TGUwx1ZVswm/5ByXh8cB9be9susRhZjStTYLaSK81kZvfGNcW3hdh9esjsR+3nNb9VFdREUi66PWo2fTrTD2m2ab4lWA9wIhkqbSSWc7/Hz7qRMaFrjPEQ6KBTC3mmuYeEYwjv5eiTBReHb8vs6Ph0gLT4pz1DlSPn5zf1yJexb9gomNezMExVYlS3KaEGcXQeKcr23Z95kFMgtkFsgskFngslkgIywumymzgjILZBbILPDUWkCEQV3kBKGReAiyK7d4+PmE9kMGXKyuBY+sAPQAAKxKnPS2SMM6pZjGJMCIIdg36c6eWoYHbrw/cIFnlTUP5DwA8uC0T+lr6TEzNuQGERaNeq22c8d2QMYrugnn8a++Zt3GO7/0n5+5oifKCs8s8BRbwEbGSckKK6LNb0ZLWLTrUwCcMtYBRiAjAL6AxCA2bHgoPC/Yj24FWxrv3oBwlkRgH+VY8Jd8CUCaHGcBPOvdMVMr2VW4lG1XkLMi2WpN8GoBWjwnCI+xKy2cNgEEM/+Rz3pv0BaAIxs6w9bdfh8/tHswL7KCtjDHWb0O5uXiKU1n4Y9xBChH7PCvKxFX/ECjXh372N/9bquj3H25ALKZ2irLl1jA3tNOQbaT+0Ra+IXI8aWv3RQbBeia9IsENBYHJQajJXR/tC5iQ5guLhs6IATczYmYWKhO0WdwZ7MkHSw3LkssoLcc1HtrlXBMFEYsjD6ncElaLS7vgrA1V3lRIqgrv9UwgGggWS8k+igi4CbWv+m3iq0kNw7qtl/grQBSbynwvLwYAEQZq4xPynB+4/rPUKUQAWu9Wm8m258tiYHXEWOC0EQCpU2AIfbVWDrP/mrYtXqwNWfBwcZVS0eD/mXNuDiv4Af9nhfnXAkXuEapG74nDnNRNFHyqkc7cmNHpO4RKDJSPe81a6HcLyph99yK17M0iHKdcQghpAMivyuS1ofEFnKtuDzPjYuzc1FjSdGtDOSd1vyBwuBeX2WoHtgCMJ/V6UYT4Ivd11fWFObtvKpx+MjC5tBw0WkdlVbIy3RRlsnSYkcazlXRkV5JkkePOkvjCa8vlJaFP3pcsgxRvFAEyA8Ebu47X+ve8nURFoRIst43NJw50M5LLa9X5MVVzt7osLM/GnbWCvi/Pgzcm8RMLRJV1SlTAfsjSl3UdwtENS1QCRujqsD4grNPlMwR1X5IREhFnQNtidOXfWDpRDuCedV41igf1wWPNn6j4SXBUfxmK+k7SIo+nZN5r6T33ZPKGXiaJLLxSamiJow/TcP0pGT+aZlzcD71J9kURRcJaOPpodBSgfaKoyOKGaLtpjYT+qxgUMrjGR0PehRnkC+OCcdl/sx5kr14VJSinBazxM5CkTxNtDBEgkDNFLVfwcdEUNSdg7pMT6jkHep1e/QZMrkVlPqDwZt/JVaorVl+bWhYPJhEz1udc+68/XDP9jvMHC0PDPd8gt2mrWfZUgLjQj00zlUk39H6vUrvVvqAEr+LEfp+dXrgy9JXfnMihP1PIiQgMZ44h3A4dRxSPquxZkO+hRdK2pyv8tn3mQUyC2QWyCyQWeBKWyAjLK60hbPyMwtkFsgs8CRagPBPKTkBYAExAOCAFwKeFx/Qd99Tngt96OKhCg8G0p70wcm0irKsnkV7M9OQUe3fcb/ZoHSbEg/ZPOAbzwwlHqp5CJuRbkX7eTZdd+NNO7Y99EAYBJMxVq6Uua9atWZtsVQuP/rw1vuu1DmycjMLPFUWSMkJC74S4sUSFAAeNuwM+wiNgbcAKz8B223ICoAygHm8EgBE2QALIS7wvAAgRSeCzYJ97c1lrrKC2u2eEjavBV5mAuJbwJm8gFoAmNTdCoJTR+ZIviNWOHMQn224KLMqV8mSMTZuuvU0sR4WU0lZs974Tz5yH6+cA4AQ260U+rdJK8uxG7Y14XZ86ftKD2dE4N63ZBLqYbw3oihoHt77WDxn3tILnavb7Zm9vzQLtNs+WdUca423eRXSmoT1SoS5jeeBWTlPjCctHFeEL8cLG57XaEZRPYoV50j3OnldaAV+XCi7Th/LykPFhGJ1uK/V8oUomt3hhYr55J8QRE44qVwtjioiP+SgYXgveRYoABHniMIunReyQSvkcyLPlCcKjhpSI/G0YFziZZmET9OpDNEBY1BUKKao1CkhJglAB4zN07Zf3XyHk5IWtJmQSchuGC8pfWipHegOQFIwtiyJ6B9qrOh+bGLDPHlSDEiruWuwOXtpw+teKseIrh532O/yxp2SJ4eROKwUnMZIKexHyiIAACAASURBVFcfLLj14S5/7Hi3P3Iyr5Hge/KrkLa3xLW1NL7jaDXq2lePSl3SvehU6q46XYsbccfsKFcS4C++RAGFWm6hX54bW0bVlvHgeNRfGh3W0v8OMUXyFJCIvetCyDCWY4lrN5WK1zQOPL6+sW94fjC0zY+jm/Qr5Fr9KlrRE1UHVjpHvL5gQqzBwsbBcF5Yi4p5Ldj33UawtiOq/2JXUMMWn0iNhg2sjgj2SjQkxJq4fRKnlni0yj4Q1XK7dNkOqL6b9Hm1ciwVWC8SR7/PRCuls2tBs8JiXakOiZjPVSCwcXkbHHG7nYMSxrYECfMJXgmQHlx/NsSzO1ULPHeYgxea71GT8LVABP+KhKhQQKd03rU0MN2KZGfWRM6aa9o0hIIrjy9CS3kiEeoSGG85B5XY36d+2yGyAp2MstoiElY5m4rrBXWCJoW0NuT7U5QNQnlcINSOpodCkskC6o+ioMpGIyOn34NJvYzvEr9YVX5J+UqGyFBrDXHhq6+Xda6ibNMnT72ms8sddR5Tveb6zcaxWd99b9fQjW/eEuc7KtJvP54fPbhDZAXXinnfeNGJtEjInVOaF6kJn9yXaTQh8Iyg7+g+4PD7EgIDbbfXKXHPYIPM+Ks0/azyf1fv96isaUO+tnlOZKGentzLm50ts0BmgcwCmQUuowUywuIyGjMrKrNAZoHMAk8HC6SaFrh//28lhPxeqMSD2x8r/XcRDIcvkLTgcfF+pZ9Ky5lKDgDidatcEycYG9jyIS60n4dlYtezkpo85AdEQMMCkO59Sg9NEes+rynRrkDD4iP/+PfvOW/my5Dhmo2br6OYjLC4DMbMinhaWSAlKyx8xXglsULZEgdAWoxfAH+IChKx0gHrICkA9lco4UFAHusRgcdCAqwmRIfdpiMd2Heu36XTkRxT7QjklsBuSQJYJXY3AC71Ari04aFoG3HvCcdBeA7ODbFCW8kLEQPRkQB4SbIgNuWa2P9psvWw32NLCAtsxnk2eH5urQDlbtm6SRgolJcF5hJKB4B5t/YRckQrld3G7W95qYkZdeIY0T2y7cm2gMSt209prqnCRAH6J/0qbAGlQlQQDioNBaU153EEIJtosSivMgRaHt+QcnXAkRLjnpDidRX+IO0oxj9DmKyvYEw9cqVYJKR2X82JJ+R9UGhGzYYhLIiZ4+s0hHMCfNUKcr1CNgjs9ToUFIcqCsSOtSLfoz81dQIRExFAt0I2GUJFHhqIRLBBfigKkuQb1C4TIEhtniRoIC3SzY6j6F1bfwJRbK2il8qAxpUqrtBOjhdEfuGhiZuWH2osX3e4sXRpyysvkzfFcqHUy4O43CMwO8pFtaAUjzTzhVq16FVPlNzKoe7c2GGRFWOdUnjp8CuMT9NMs0Jfr13+uH5LHDsuoqIgse6uStjTO9LqHx+P4mW12F0kvqJsjCzRkTBX6K/FwbLRYGBvt1tvFpyq1drpVhvxPBhWmV1oiegMnTuKiyceKy058KLRh3asbh7c48XRYRn1ZlFNq7uD2vzuYq1YjFr6F0oteomulvgRzyu3/PxNuXwj/IqzZdbsYHTXvNbIwfnN4WGN8HGVz28fO0dF6WKOVmPBtVUJig8WHn7kmGaLXeoUmwT6b9JVXaX3C7WvLA+CgqgoRxoYHXLPKeqEffLjaelvVnJy6TyU9QlvBdd4NjCXDqRno88x19Af+ownBRs9hJ5og4EmYaBOycYnYt2B6SnMc7EJ88V8xrVAkhs9jbuUDuq4pUrbokF56vjqc2XN7y2nEB2TeTinwk0Z29a0ryHChToqvJO+KwbylYCA8PNOZ4THBSLdkZKnubHozPNKznwRG534duChYWgWaAv9qZycUYlJfjX6+rZHZaGPsdgQGOhu5J3Fjc5V1fHVL7k6KvcudJuV7aWjD31qwWd/jZZbvSWswTxsveJaIi9OhdzCeB+44IU8doxclteUxOAK1URG3KVXNDj+r9J/VbpZiXvr9enJ/pte/07pr5T3z7jK5woVdVkqmBWSWSCzQGaBzAKZBZ4CC2SExVNg9OyUmQUyC2QWuNIWSAmD4yILQB42KvEQCwj3CqVPz5S0aBPX5qHWgArtW+pdwYMfq8PMMtB24kHfs4+VYayuJh/eFbwHyCPe81eUcHW/YGHZ9Zuvv5EwTY88SYLb6zZee71AxViEBeRNtmUWeEZbAJIijUlPOwBzAHcAvawXAqAmAI8V7QTMX6oEGcHvRwB8gDPGM0AdgAqfLeAPcEriGFb+JtHQr+zGPATwT70BayEdmIOYd5hz+I7wSwjn0h5C0ZGYg/ieeY6wKoR8oo0QFrSBDTvQZuYxu1J3Knlrg7dYwgeyBntuyueLi5oNRc5J7EOy9Af7KGdc12RU+hXTrphN65C9PHUW4Dqlq+kFwycwKv2Ba8l++gvvGUMQBIRnasqtQXGjvGroxnUtPe+Sew0r4k0WdRYkpwn/r2Xrfq4YhQtKbjhQVKglQ1G4Xq6pxf3cd0RSIPmQtD7RlUlWzYsS0Wewe+7xANfajAwyQL0RcddnZJIHnUgOEqJA5F0hAeRoo7KxaIDFDU0RFy2RFmfchyEQ5HFheyuVUB6to091bb5x8ofn7Gxcu6kWd7686XbNk1r2omK+NVDM11yvWa83G/ptkA+bBbd5stsdOtmXHz5WdicOdeYnjnZ4E5J2EMmjtkJWTLcpRFSrzxsa7s0Nj8zOHz1yvLno2NHmwo0TTs+q0Ct1KE6UjvbA+TvGwr7547Xhk/35KmPWlKtkQ9GtSq8TPg3MDd63etdX6tXCI0tax8e7ovqRYtx6gedFz9HMePWc1qgTNHLO4eJsZ1iouMJDuaFf7DiZL/3wiajzeTr+kd6w+m3NaIDLj+oSHnBvdSrxF3UNPNMvDFUw2PdGp9jc7cxadeCIH4wOy0fnAYWJWqpfP9dGFef5suYmeQ0sFh9VpAfJDtLqMAB+LGKjIx4zJMR8pboosaL2z4F8Mdc/p7YlYZtQEqFfSZ9E/+OxYGduO0MlcH3D9FQ8HSJdl8DMg5CvhMEjrCY6ExDV/NZjMckB1QUyQ91YfFtBTkH71Qs5T13hrAKnK2yaPgdtNyRSpY7iSDxifm/O1bFzVJdZGi2z1NE7uVSIbENG6ILhrbNdNelQa+forAt0dvKXTZQ02UFlDSh/p3qz0Ukx44b6q20qe77OV45z/tKJNS9x64uuWyTCqdH/0Ifu6dr5pXJu/Cj3JeZ75lMbZpBS7Li1GkSmz0NgQFog3q1XI+LNxvunaKMPEZrwnUrcR9B8+w0lBqMlLn5X72/g+om4+BT5nw5hn1QXazL6KffVsUzU+ynqRdlpMwtkFsgs8Ay3QEZYPMMvYFb9zAKZBTILnMcCgHG/r/SbSoRkYqUWIAax0nlov6StjdCwa/dMeSmRAXgDWUG6RQkw04rUsrL5s0rfVrool/WNCgfFubZtfXIEt9du3HL9vid27axMjE8+jV2S8bKDMws8iRZIvSjsGQFuCE2UiAgnYCvAAkATgD2JzzYUFO8B+CEleG/DzhArHW8LABWIDEBCS3AADAF+WRJjcgX3FWw2bWGlM4KjbJzbamnw+Qkl3BbIg7cFhAZtoZ7UFxKV8W2/B9RKxIxPeWZYDw2tHDYr7tu3+I8/fC+2tUApmj1rlBYaqC7ddJx5F7aaiARDoOyPwvBoq1kf2/fYgxdM3k6pQ/bxSllArgOGHFAkJ50iIeA8A96n/QCpYdOP5HEU57WzIK+KfN3xJxQzZ0Thh1p51x+RJPC4Bp+AdK0tN5IThnNQr3B9xQNaEHpuo+blRpQn6TNanm5OAVeQ5jecBMGB+GwC5wjelVK04Q7NiztXzgddOkbC2JJ9lpK3yWNIj7ioPNdo34v1AVAXjasJkRZ2UUJovUySrjrpcWGq+u6HXtH6o71/OyuOcqsiL7fKCxovEPVyXdzR3ZmLmuWY4FGqshtXB8te9f7+3MkTc/OHhublD1S6cuOtsldv5LxWi8obqgXlhGTjPULNxszphmEMfl/yavU5hcMHFUqqeqI5/8RoNPuqStyxTB4mni5JsR53zq2F5c4+wHNamwiBm2ddXThFZHNj8T8tz/e6gkbU3XRy+W+V15xcWJh3clXz8HcXuSd3lePmPQpJdXO50VzX50xcvSp3qLwzLwaiZ0AEhhxrFMur5hY7j/p9W/rylaWz/bHndjVq9+iq74u/YH5TTaBPod9AnLcy58R7x/T5iOs3K4RAEjmxQFelFPc6gXxejihSFtoQx6OS06va9qmcbv1K6pLfDD4FkBjz1fg+Q4Ghe5F4HyR+CLxPAvchtp3Qxsx2TaM1ge8EuinMRQ2VO6z3De2hfonnWGxChh3UPsIQ7UzzM48bkXWVXtE+RTKTLeWr4inJ4cT3VHp81KlGO/VdTUSrwkCJiKlFEyZsmPRXpOHhOsMaJXjYden4lXLNWaFL2iV98wiWDuoaAiOsab6VBob8goZF5XVCaKiXFkSAyErOQr32Gw8MPDJckST0Fd8IdRNiaiAqdnU15lyjIkNFFJtwew7d0Z+rHlmh3t4UUdKjYwZ1OhPeTKkgMxpPX32g30PWMJ8z/zdFUmCPRkpWmFrqvRnrkBnVNyX9tOMDF/eb1Xbo871OCRlF/dCkIATUG5R+SekdStyj2X4kTXhU/4Xy/aFeK08DMW360DpsrcQzB7/5sy2zQGaBzAKZBTILXJAFMsLigsyVZc4skFkgs8AzywKpp8V+PTz/D9X8VemDDQ9n87VvWN+nSzZPtSsV0rYiovYVEJK8ZoVpG1FxLoOwuoowSoAghIThQZHwLAB0H1MCPLzo1cToVwyePH7syMEDkDLTbtff9IJbatVK5VLDOOHJcc2Gzdd+5T8/bWNXP7M6QlbbzAIJYMNmYS0bLsPG+bahm9q1KFg9SwJ8gMxgHFtvK8buMiVibOPBgEcG3xEeilXNzB3MNSR73it1HSy6CVxHog7UG8LCrjGGGCUUHaAiwBSfISYgJAD1AK8sqMJ3FsziePKkq+uTwCrTkBW2bZSFLURSOJuUblTqDVpNW0eAVKQP4jAM9guYZWXz4UatMjw2eLS284G7ngxi50pdh+/bctvDRJU+OZYQF4mGBa8kQkbZde0JUK5QOIhua6AUJWLBVe/U4ENzYq48CxYBOye4PP0BFQCB8k4kge0g9ORE0YidwXocBYHYLGXDa8LEEEviJoFgp+a2sZQMu6CdOOkUynlJfPcqf6+0KtRn0b/watK60Cp91sH7UlmIblZZElF20XKhNPouW2RCYCX356A9XJTa7r1jd9QplY6NKuMHnVxpkxbfXyvubo6rU0itQ7RMtSEFnFrRdx/uzVW+sqB48NCq8raJntxYHm0cz/OsN1dBVea3BfbSkQaQ7hEX43oG1TaUhjFxok8uYQSvWisXq4cURmp8b92NamFpnkwkvQo334hLAyItusNYN2xVMOUFzbxHEYbE8NxCLu8VRD4QWomx2H0kNzByND/Q0KjdvaJx9NDi5omTS1on9nfH9UOL64NXjea6Fx2plzsbTd9FkIFtKN9TPOzXFvS2KguWNlpLC15wXNaDFDiunoCnggTTC9VivPeg4Pz9btgc1L7ZatIypYKuymy3y5kdz9J1TYTb4aCKIiUkN+3UJb5dFFif6FtIj4Mc8nBIZtWkt0E/oAcBJSFN9zTUHT4WCWlSVV7eU35VVxKAHk8JvCoOa5/ktU1JeFAwpyUedYRzgoCGEFC/FQVHfsrhdUJ1iFRvV3B57EshI3xCxIV+1cUnZV8Fkkq4Jaely4YQ97BOkOMS6o+az9LEWvICJy/XGl0ziXTjZRQ4dZEdkClDGEIy8b6InW5pd4yqlr2El1IP6VMJ3WqrSDjzWorzfq7Zu0KS6ZLnCCtO18lvhPni6Gq3rLk20O/NmvHyqKhxTZWLlbFgj9rU0GWETElCpyW/TfmdOqY6T+gYQ1Tzqs94u3TVb3PUd0WmED7tTY7Cuk0S2+RtitAIEfbmMnIt9fmyEs+p58SECIl3qXhCRRFm9a1KkBh243f+WqX/rXz36ZgzvKLb8l7pt/xWwCuERQGEuTJzzDT6HVe6Hln5mQUyC2QWyCzwDLZARlg8gy9eVvXMApkFMgvM1AIiGGoiIvBo4GH0RUqEiXqv9h2yehN6b8PCsJKaBzs8I16oRGgJVt0B8hHr/VOId+sVsG8SXJuGxCD/Y0qAdqzg48HwTqWvKwEAXhIwt+HaG577yNb7ifM77fbK177htv/1F3/7gZGhwZMv2ryC+l/0huC29LY7HnnwvrOe71yFc+zc+QsX7d+z+/GLrkR2YGaBC7BAm4i2JSoYb7znt58NEceYtIAh+wD4eQW8gojAgwIygnwQD5CQVqKV8mwYKOYOGyqJ7y3RmYaouYCKX3xWACLmN+Yv62GBtwSC2lZallfawX6IC15ZbZyGzkmjpZ+KRW/hwQQitITtmZ4V7bVm7gSsWa8EYUvYnaL0lTk+AYSTmY/PewSZ7tQq+EplbLh5YNcjQa3KtJltT2sLTIotTF5HS1rQBxlPFviXNEXc0odaPo7G++Ogu1excApx1Cs0faDl+iI0tJ2KhyQ5g7irHIdzfYW3CZ384UbsNSSQMKo89Fv6N+PLjukpZoLESImMpsKPkUz0f+Gsbk6gc3xc35flXSG5DMPj4QF0i/Z9VeVzP2e8Wk8gxrMVnrdKCHh5MD9s0TEv1eutTiG/Oi4UynG1GjkTtYZcJuSH0DEUhc0HJJnxRdeP75xdODYisoJx0ZlqthjdKyW8s2gXdoMgZP4R2B9L84BF9BLNUOAgreBPxkxbq3vyI+N9wdDRkWD2cCMs5iM/n5NeSF896uyrRZ0d0sdgIFnPT0M24gkQhHEubGq9f3KNmN+wKW03K9n3FOePHSzM2T2W2/eEyIvPCtgudzcqr22EJ14S5nrnV/yiol6p+qJEDgWSUVBR3U51/pzc6Dwvr9yomxBCKTTjGy8A1VvGjjTHJMQAHgd9Jp8IBXlVQBzk0pp6xicEC6MgwZ9VX7B+XUDrqdKE1ETEyxjqgpBQVUOYuPISSwKWyRxalFLQ/JY3tsWC/O6y2g0QBGyQK4uV+J2HZDZ0REI4sz/53YdGh+YqEz5vRD0c3QxEsSNvqciA+U4j3KOesd2EevJFvHB9E/YMvQpAa9d4cHTpomKXnAg8+h7zJOdClDshO/TqiX6R7vmo6LUxUWueiJuSesmAztqrtvTrdRGeKnGxo+f46t9yqv3XO8WJ3Urbim6hucrrEdkRiFKRqoY0NKRprzrIG0WvJaW80oiGyQGdjd+FEPVYFDKbulEf7LVXdeX3K6GlVij16jj2Yz/IHMhtQjax8OaQyArreWvIN30eEWkxNWSgMfilbClxMSoCgNCkv6CEQPdLlG5Py32ZXkl/rjz/R68HdMxlr8d52sB15NpiC+7HDz8NPD4uxezZsZkFMgtkFsgs8BRZICMsniLDZ6fNLJBZILPAk20BEQojIhr+TefdooQ7uXWTj1NhbPa/UQmX87NteGkQN5cYER9U2qpEGJUzPDW0j4ek7yjxIMjDMMAhq9pqM/TQOGsl5i9avHTW7Lnztj94dsJiYPYcVoo7e3bv5KHzkrb1m69jlbSz/aEHEOi94O3tf/gXf730qlWrb3v1j/zgBR+cHZBZ4AIs0EZUABoZuCw9HLAMAAEygvEPUMh3kBD8HuSVcQqQaD0jgMcsZMaxgDvAaQA2bOSzvyXtuSwYeBZQ9QIaM/OsgHF4VQAasaKTOjEv4dG1VwkQijaz4hRwkrx4UUBaQG7w2YZ+svW34bAmw0Gdw6vCUSgoasuxVqPCgteNRC8ElDPlaA3grbXeChskGFUrkCNnfORk9PC3vxDu2bn1sq7MnbkJs5wztUD9x8/g4fBIsIRdsqo96Qu+lqwP1hy/JjHtkeVRbWlXHC7TBS4oTJRfUw5waVDdhGeIFcXGkTeFx8pvFvPTR0qKGdQUwEu5EAeIaLeNrRTmba988i2xonRf1nryKMrrdIT30YIDQlGhK6NMhaLvNOsrdPL/ov14YHB/5l6usWBoAuaDvNrGuFKdRHaEIfHzXy1YmfCSVzmtoFOeHBAZnOcJteHRyPUfbUW5h123uK0jV923srwDDw/GJKv0raYA45D31gMrEQtPxmoxRJaZ1flh3JMreHhlqKrIgiTiOwpKpNBS1aGyN3FMwt89oZfvjiK/WIm6540Es4525iYqkj23hIVW2Bt/BYHwqiG1IaySPGDkycE479a+UEX3aGdVRFLwcHnF2GPFxRU3jIavah79dH9rfLwcNm89UJi1otHTK0FuuRHkis6JsM95ZNaK3Jr4oLMoOCmJdV1IX6vxteo/KmlxfqyISoF0OnwB9JbWsvQpVwmrUEvr52bfM8Ma/xbjeQDMnzN0gvV3kBKHK/hcBEHOTCeUEjm9ugqUSGimlpraI3n1llKiw6PPKkmBpYyWBUGl6AaRLKP+YeyOx4YoApO4GuhxlFQiBEuv/IcWqYyjygOJgQfHuM7bGG84je45Iga2iLAQxSWdi0AdmVIctyIT4EXjGfIL8kKa8hJtd52jOn2/6jlX+xZQN7Q71Pw+9C7yktjmMol4oI2RUl1nbKquFZEwpbjTK1T71vm13i2d+dpBp3//Pzndx7+ky1ovqzWLRG0M6PxBTjZSULRQdeeyw4LR7kAMySbZCk0QUWNmRDXxbkGfQ12NsFVVPEQCvFtUL7EeJbVBfUQjQL4a6lkn9X0SUtA19xW8a/arLejP4F2SkycG43hEiXvRIZ0Z4oZQVaZfXorQd0pcMF62ipggpBtaKiS7vV1vIC7u1PeQGYcvRZhbZdjwkc4MvCT4jUAIWrwMIXVof7ZlFsgskFkgs0BmgQu2QEZYXLDJsgMyC2QWyCzwzLWAiIJxkRN/oRYgQDmCQLY+Axhcq/SvSgIyZrQh/GeUOLX9jtJ7VE7Vemu0ERI8cm8jzJT9bkalnycTgttkOZfHwwff+67b7/zi5z59Obwa1m+57sYwCILvbd/Gg+EFbYVCsXjry37iNZ/52L/8fxd0YJY5s8AFWiDVpLBEBbCYJRHsaxLu45SoNGdg/LP6me8g+QAbICqAzGwYJD5DaJAXjwtLWLTXkPNaoPZKkhXWM8ueg88AuYScgBQF0gPIwQuMVah4T9BmVnqyf5KoTfMCxnK8bWv7K+3jsxbEn6FX0d523luygt/WVtgVGBJ81cSet7H5kR+AsCAslDZFhgqisaETsciKqWVmn58hFiBsUhpGif5ixwLvK1XXr/bFrYn5UaPbkA+gpJIEyLMUXahpGmZIwK7rgU6jKawOFwVC6RV7rIw4hWLyjxvljOm2U3oP7d4ayg3/AQ8ieDUQcu7EewTYz1NPVCAiXyoJRLiROoHvvVC5EOJGfB4ST+GDYkg8xrnGEzC0EXVert58i7mb+/nlIkF8p1YTNF0XAB5xzDdV/bvUtbeFTulQze8a+eYPvzz8ZlLnyVXeEvG24Cf14xx8tiGcVA+3oNBSSdXjuD9oikjwQvIxxhhf6IPU8259TKGhTtairqWRK4UFN/LrYXnuqNu3YE54+FDRa1CmgeX1X3JNbEQtIH52emqXLkeYGBcAm/mNj3MaXqHmFVwRF8sOX109eEdvWBkrR62XN5qtNVHkFuAcq37J2VtcHBbrYaOrVvX7WhXKcCK/HCr6VpBrVSRVLXge4Doy4Lan2aZbrRAkr734QcgrwcwYhCIKRZ4GepX4NMC+jhkUWD+hI+dJJ2KRW9dREt9Q1C+pcegKJL5sXEgTvk8MGUUR+qmppuLZkdNx/SY8lMB37KHAYngKJGSO8og2bYq2kTa8agaZkTOAexKuU+SBoWBELEi6fblorCHEulWnQeU/qjKPdJ/U78oRI59tgmGJUMBjBNFs6lbVcV36Zra6ab/KOql0RIQAIZaasnNFdT+plMfmOmKJzj1b35cIJcXwMO0QYSHyIlZZ5agqz5ig0NeKF4tZkD9SXly0VCn8qqZytFpEwIhay6mdhNFyffVe2c0YxsjRpx3JBm0ycjCW90vILB2UdFpiVplwZOmdTSo2phyFrZoHbabdJa6BBjX13Ck7neCqqt7YDeJjWH1st47ao8BsEIKE5mI8jcoL41hKLNmRHV6MyDfeCyIU0IODIHitEmGj2LiXvyVNv6E8H9X7IxdCXKQC2tYrk3oOsm860qItL7/P8b7kfnu30pPt4ZE2P3vJLJBZILNAZoFnugUywuKZfgWz+mcWyCyQWeDCLbBPh+xPyQruAzcofWOaYv679gH08RDECinAzB9TumpK3j9JP+OazoPwGdvlJCsoHI8HkL5zeTzw/e6dO7ZfuHnOPAKCREU93GzUk5WKF7ARuqqzq7vngXu+neI2F3BwljWzwAwtkJIViQTrqVX+AAxWUBvCAVAL4I8VoSTem7jeSoAbhOkgTArHMJYB+8jDmAfIA4A423YlSYr2c04lLPgO0mGHkiUrmK8IQ4c+BPWirdarwhIWJnSHEuXZVwukQlAYwC5d0H02qHiqLSB0KBc7WR2LpUTObxMRThAwhQpSzY5InuBArTI+MXhkf9jbO9sdHQUvzrZnogVSnYt24oJmGI8LVnePuPmJ7jg4IOR/dykO1xXcuMsX8mti8xgkGQA93ylcFqWEUXlnFBTqKK8YO/kgDA2on2QEETfrzxMzWcLCfGzn8QzMCkif9mutd09C2Ei/IV6vwDWCc7Vm3cut1tryJVq+8DwdLlLeVbgb1u9TWEzoG40f90V6L90Nr9/J5+c7pQ5kIgQ5NwSwB0+o4nhTSpvK5Z4Lclyv/ziY7embyAq7w2rDMFaStf4JwYrHE+OI8TeeEoVdWv0OmE2YGbw+GFtVzw29olcfFR0YKMk6ioMU5QcqQdc8hYXqLHhNeVZITeOUJtjJ3gAAIABJREFUF9jpc5RqR2QsMzYBpeUZYewFjcC8KPKiUPbntRQC6fH8woO5QvgtiY54bjNUiCR/YxhHPdI3j8NS2dsfzB/t9CrNDfG+hTmh+pHbMahZQPoQ4QKV2KMr92WVCXk6R+Vu1OeiAPOKviMkUxKKq6U5zBXx6hkvMMIwTeg9E8Lj0aDaPOasj2rOGol1LxX9tDjXKT0M+bcEefUx0S5cSbwFZETmdFIc1p0NCh21Am8IP3L6ZACIAOmKy7aIaifEBARQrAMrmvmHVLMTSiPoQKgpXaofQZ6IL6YATybEJwRGRXn26/s9Mt+g6tMb1wzxMKr8aEf0q41N1Wu7Xjdp3006GrFrPF75DcqiGa4pxMmjyg9R8Tx1VMJQzVHP4n4lvk7eGGkoJh0Lqa7QTF6+1r/JPXHdO0RjSdqiOeHkhoZit66m2IBp9HpKUJKXhCGGIBtS5RnDD6UyKYl3k5ycUmbLNXnULxhiViDcdGTIoITncnIIgzMMtS9QXrgvERer9WaVceJRF9BZ8dxwcznnxRIYhzAi/OCjyrPTvErsXnnpE/a+yn2MMXrBWxpy6YhIg/fo4C8o8Xv81raC3qn3/KZ/m/J8Tvmn/a1+lhPTfH4jUM9JT4tp8mIafj/gXcG12qPEQoJsyyyQWSCzQGaBzAIXZYGMsLgos2UHZRbILJBZ4JlrgZQ8sEACYVJ+ZkprEMT+F6W9SjxM4fZuV0L+ud7zGPjLSv+t7ThIiyXypPhjlW+Fa6+YkdZvuvYGPCfGRkcIN3XGls8XCtds3Hzdtgfu/e5MKlEolkpnIyPwkFi9bsPmT/7rP//DTMqammfVmnU8vJ3TG+Riys2OySzQFv4JY9hAI3hDkACsGLcAB5ARJOAcSDfGTRoaxhARJAs0EFcePMcCDXgmWK8MyIuz/Xa8UoSFQfeVbPxw6xFiOwDnpZ18T7sIV7JXiXkIAgNbYBvKsCFijNeEEp4VRjQ1/c6UJZSJ7802A8+K9npwLuxKHZfo+izWInnisxtQFPTK97X4OApZtf6Q9u1UGpYgd7UyNqSQJCYMT7Y9wy1giQuaYb0u5F1RF7Z9QumI0kGhflvDoLm2LJ0A3G+IV0MHCfRGsXxKgsV76pGnKEj+IJ1Si/DroSt4HAIxFtmV9GVFmtI6ck9oPZkm6QHe2DXh+sbwH2bTinr3iDnGiRAvXuIUCtIioAxP9/X8Cnlb9KiDTqhCzBMNlSkAVce7/hod26HvWH/eYeIzOa7CA7l4ZeDJdK/eP6IOfrL+yp7J8TP1Uv7q5jsckRbWi4lz2LrZMYoDisTJjUcTY1P8jVMRBqxV/yImTCAkEwYpKHm1PmlVHJQHwWAzdGd7ofD6nGgFr9zTdDolej0uABix+1SnPF1bn/A8cDGnTAbKT5C2CG+HZNPI1UQghFrhn+aKwSwo+lKg4FRDXhztEJjdpZXzVylcVXdLphj1Ojvv71w1MuGV/n1V0Bwr56/yy42dj8t0kCv8ZnpQpzyuRPkLZft+nZ/5GIAa8gaAG6KCsEHMY1xj5qeqvAQGlXx5FjwSjmrhSOAsVU9YLr0LwhotVvt7lLNHJfdGUntQWwhFhJh1t0B0PGP6CLekFuNNQgXyAtTzsjBEidy8jKMPJglU7jyVtVx+Ctie65RXOKWSbBZqX4Lzq0y6rGbcTequQ8pVdXsUyqmlubPpVIOCzt+UgLiO9UJnRMf1q+x5AvmZAq9V/rGWhE5kbmwI1XSDAP1O1WGRzo+tOrj6EAdiOKTdbkgTvEE4rx8WO5yR637Wacy6WvIgTaf30U86HbvulmeFDmD2bQ9kyNWX7Lx6cD0aUz+qiWhI7gd4d7RULu9pn7goeZvo/qhzcwMoKl+n9o2o1YSHoj39qnMBQXHV13ip6Ps+ha8ihBa+M8if0x6naAMppr2bnSKJ0AfpVhmrVdZNKuOw+tEelX1InyeUZb+8LgD5IakqOG7kJead9scZvRAqSoQE5P0rlNCh+0ul56cHYxl+39+rPD+pV+7xrXPpS6SeFKHyc4/kdwB1O2PhTupdgS2Xm56UlE2Iqgte5DOjhmaZMgtkFsgskFngWWGBjLB4VlzmrJGZBTILZBY40wIiF3i4YEU12hVsPCC/X+kBJVa+8RDNKrAkNEACCNpV17+p9x9Sep3Sr6Xfo33xSyp3oUiLKxazlvgq6zZfd8OdX/rPz5ztur7259781rf93p/+5Wt/5AXXfm/7w9OGcfJzudwbf/nX3v7aN775rbPmzJv/2CMPbf3l17/yJYh0t5e7Zv3GLblcPr9t6324tpsN/YzXvOG2X563YNHir37+M3d88ytfQNB8cnvlT/3Mz9/68lf9ZKvZbC6TdgXeHr/+P/+UB0fhPVE0NHji+F//2f96R7VSAaDItswCF2SBlKiwoZ8sVAn4BUnBK8AEoDljnFfIClYn85k+xzjGY2qNEoAaq5YhLEiMfRvShnpBatqwLU/V70ZAG8JoUG/qk8BrFtBMSFXaRR6rS2HnqlSidvIYQDi7uhtQDlCwnWw5K9iKMc6xYTNrS+q4XGSFwqCYsDaTsgOad5ywESj+ufs51WgHYGyjNtEcPLY/GBsfvNhzn6dq2ddPlQUsebH2w/cGWuQ9KjbspFZ6HxKA+iVpMTeE/i7Wwnihkrr02hkI3ZVDRK4jCgWORsI4FWxH9+DQL40MxXnGN+NTq+8FDZuxHTN25TGRwu8mfo0JcJMEv2kPF5UYgXGxX4REpyB5BSWS10TYEhyuaSMv4QU3mi8CxNyozPjiNQpZUc8afuYPMSrNIX0WWeE9ouO/oXIExrsArWPKnxNJYz2W4rT9p5kf0kIbY3gSjE1JDDsuATmZaxKSEZ0Fx8UOnJ9V6BxXLHitVm9ueJeMs6baKswXi9GtnYVQOgYTofwavUK+w1ewnnSpuyUurLeTMRPCIcmreMTJkHaiKoTOC76WQDd1RSzcen0U3bw/EjejvaJHAPy7AkWeyhe9ngmv3Lm1c9XBQ1H+vs3OvL0Fz9nZr4hVHWFDIHlc1xL/Uc0ElWLc4pIPqGXd+nUF4D+qK0kXoDzmI0hXtkR4m+X7S2TlJc6YVNx3B3c7D4msWCRlkh06ZrnbULioquZ4XyRpXmRIzqnrspdFGizRpexWXoSwJekhgB1tCW0CzcWbJeSM8SxIk/YRvknsiPEmEEFkwh7hbZLsS/QxiGaWVtB4d9SVSr5CVVGiSIoGFJj4gySffkG2ZABDq7kKO6pCpNKCy5CvHsjJV+XxXkh93yDvjAMRFxwiQOenHPapM4T1+Vui4S0/rQ6r4iR20rHrq2PR0Fiku15eTINMpFqUTfsYWI4oo5x6LiGiair7qLxUICpQG2nKDoTT6hIJ4at82lZRPWH4yjoduhonVd6E9pe1H8+RLn1X1/FjcFmqW29DobZkG+mhOB0iISAxQhXqQXzoe4UbM94Y4rpMr4a8gay6ylfXUiVOqA779c2I6rNfxz6u93hgHNbXJ2pvcg6/7lVO9Q58m2e4pQQEY+huEQl4WaBl8ddKzB1shGxivEJe/K7y7J5BmCgGgl3MQB2nu1dBNjG/8HuY+zEeJdmWWSCzQGaBzAKZBS7aAk/Vg+dFVzg7MLNAZoHMApkFLpsFWDmNxwQPL7jp85AEIMJDCeFUCPEwXQgYQAQeqllVyUouSI3/21arHSItAEIJ7WC2SxXZbm/x0hUrr1aEpd5z6VccP3bUrA5fvHT5VdMRFnhNvPuDH/30TT/wolshHEaHhwZf9bqf+4U3vPlXfv2vb//932o/3/ot1z+Hz5aw2HLjTc//qw/86yf7BmYBRsav+MmffuMvvvblL77vO9/8uj1u0/XPuVl8SL46MT4+Z96ChWMjw0PzFy1Zmpfrh7R3vY7OLh7ssi2zwAVbICUrAJoYq3YdJ+CB3WfXWUMyAIDx2a5kZoUkxAVhNwaUliixj/eQGgBllMMcQB4AF3uOC67rZTqA+gOWWFFtyBjAEIBLPMB4D5jJmAcg4T2gCe1gvS3fM49BTrRL3FKmDQ9FVY0jxCXUmeuBpwp2I4zeAj9X8APFk2nffGHCTqMOwfJ1XcvRMGw1R04ekf7xmeFzLqEu2aFPPwsYhXX9o28eCmL3XsWeKWtV/8tKAjJbxK0xHEOgJfLqplHYVXQV10gBh+i7kgc4cK/fi7Q1hAR9nL5O/12vgxjHvLf9WX3RiFaf2hJQ3m7qlO5jOofkhcUFMA8YMgL1gyS+jcgIKsP4AXZtCL3nfp54QbjuTh23TeQGXhUKASVPi2SOgbBjLrLeAYHIC3PW6YiLKZfIAqDkZ6y3h3KiLYxhCElqRzshECJ5WYS1sHPbeNg7J++11vjBuAgLpzAaD/T2eYNehy9daERk8kn7hW8bffDTdMuT+YWBCrBcmOR4Ug8MQ/8AQPMdJ2/FVV23J/R5rkiOJQpHlQ+QkwYg972bh/3yyL1O+UDLXxi0ci+YWNAarBcVmCjwCsHu4oLg6sah1o+N3XPQtAVPBbFS7g+pZ3z5jN9b7XNS8l4r+HM3iktQ+CXVmnBLh+SX1a0ZTzSB0YhYYjQk0LyoOxv1eaWSdErMdeyW10WXSAw8AeQyYWoAKZEzvjts8GYpz6UeYAS9sRtkARVAe8Kwu2l4JPLIswIPiORQSZvnekRwJ4LhhGMyMap0kAk+RQglzitvC+OJYLqcqJq8gk5JEcVptpwJ+rjKLSlDjvBVIgbs3N2KCl2VwS0/W5LqdW8sF5j+bR99ovvg3Y9FQVhWr+kxShwiCNTCRXFBIbDS8+pzQV4gA6rrY9L/eFz56jo/5D7hsEz/Ml4jeJ8kfdmIw5MH9gLyRom83FfxvuB745lnvDMIYxUZWzNe1STdS3WtTGgs3RNEVvSY4GTKII8VQ84QXkqEzCylPogzAqxJ5wLvmu+pzN165Xf5Nz/8CWeHBtaFhHBKL6bE6Zb01ERI/Lt23KP0i0rtv29fo88/qPQq5XlcedHXcKZqVKTeE9xvsRe/DRjvjMX2jctJmC/ug3zHXDD5DDAlb/Yxs0BmgcwCmQUyC8zIAhlhMSMzZZkyC2QWyCzw/WUBPRjzgHaN0gvSlvHgtUuJBzY8Er6lNLn63xIOOq59s8DCP2snDyt4Z7AB2uFN8PNK54p5f1FGRb+CA7c/eD8PYNNuCrFizrv78ccgU87Yfuf2d78PsuK3f+W213/+Ux9HbNzBE+L1b3rLr77vr27/g/bwUJuvf+7NE+Njo3t373zs6mvWb3zvh+74/IG9u3fd9l9/9BY5XuQ/+oVvPfian7ntl9sJiz/8zV/5BcrEi+Pbjx0e/8S/fPD97/qj3/mNi2pwdlBmgdMtYBaeKlmhbKvFYAEUxiWgCWMccIW8/N6DmABMx4uCjXL4HuISEgNwMondnrwCOFgY60pdA4P/pXVpP5eFVm2oJuoE+QJowupOwBsAW94DspiVrkq0GfDRho/iM2VZ29iwMzYkDe1ihfWlEBXOH3/43mTtbHJ+wOMfUpovUW2DySUruEGqhNk1G4S1McSKFq8PS3A7rowOhzsevPOS6nClLlBW7mWzgO2HAJL75dqgoPtG42DUDeNuFtGz/D3BpBmbUq+I43WdTjiiCP3fPiFYW0h6JL0LGADKoA/pozugvkW/YxwJLk49rGKRDZ5fkN6EigI5Np4CyWhI+rtA4Ph78rTQmHKXO0FrwJQVhWgsaCF7lMarl5ZLbLw89qTnUOii+IAIDdVB0saxdBTiUHOLSBRXa/0T7RfAf44B+DVEREpcmPfn8Lrg6yj1tqA9aaXNPGQ/pxB60l5VVVhwcFQa2CN1r6NYEuETh0FpLOiZ350buW9W4bhs7HRHxNqSnfy8V8hpWb8J9ZQKe6vu+KckcbMIeNV2yY0IAeYyrIWxjKmjPo7rY7LIw3VXiwTp8nOem8+VunJRz83V1nDYiCe82Cvu31NaiC3Q4wB4rz9eXFR/z5yfmPQuSU53Bws7zjUHQGgkFIPsIn8PK5yteui6z8JnwCkrPNQRtaEotZJ+eRQcEJmxWp/nyIIlHYknTpdOQqijbpWm8GLA6s6oepAUJpxZOn5AVoc9pS52/s3jiWCIjCRUFDoPgPe+ZriKviN0GCGnijpnHBUFVOeNJkePLlApaIrvKDlDKpsO3K8emWvJw0Iofw0xbZU5ok5zQBf5qMrEm4PgTr7ICggi6f8YLxvpbbjjleU/2Dm+5kd/FLJCeutjpYP3fttp1faqTrSlW8HSPIXOKujTuOq10iuIVKIlIkREGHSp1UvlATIcn3S+l9rS6GjDSRhyRufVZ3NtksnbGAJdk+TKE/gpNuMMAoh8yTWhLa4zpjbwHb46LZE8CSESO/fpfUFtnaX3i5Xmq9P249Rk1EGgrNTT1eiC7NWlt32q+xrlI1TW83SG+6u3iXBwnW1lwoP93Tn7SdKd2jbCROnjPhEPv6fXv1d6vdKfpVm4//N7H6ICwW7cn6b73W76rhLeg13KO56Wa8/EggcWKkEk8mxxp5IZv9MJdJ9RyWxHZoHMApkFMgtkFpjGAhlhkXWLzAKZBTILPDstwPz/yramE+/9uBIAJiv/ziaebQ6ZQlzwcPNBJR7e/iEtkweiP1LiodDkv1xeFus2XXdDELRa33v0EWJnT7ut3bjl+opYhn27Hzfnb99e/KOveNUrXvP6n/vge991uyUr+B7PCpETz5uqZbHxuhtvekTkiGQuyu98/4f//fiRQwff/FMv+yGrn1Gv1aoLFi9dNl1FVq5eux59jO0PbcVjJdsyC8zIAqcJNKfrnXWgxdFsuCYrpg2xwAaYwLgFf2EfBAQbYB9kBSsjr1ZargSAAeDJSma8KwAhIAXY2kGzduxuRnWfpoz246aWRz0AN4Fu2gkL5hJWadoV1XgsWBKG+QmSgsT4JgQU89ZaJcBS2mTjr1Mm9rK6FJMgYeqpciEaFWdtP4LnLOJWBuvZsVzvO4gxYzexIgnSKMZCefFk0eplt6GPzYmRwSng5YWYOsv7TLDA7/70jRBb9E/6NGOMleriKERcOGGHL887UGDTWUUwRLEb59xwTi72ehVUf1QsV6Rl5XHg5oYk8kAZqfaBe8zAwNx/FRJJ0wRjn/GkVe8K+xS0BOQS1ceML1QEJskzoc8aO7FWQcdHhfLP06ywQN8vTTQuBC9TT2BwCBLX3adXAdMGvB918iXg6wVOqyGCIzespfeDqnhF3zMPTSiPBdd5tURiUs/zbGnIKI6DvCC3JSuwH8PIziOGJMy5wXE5p4y03FKhEvU6laBcrDndS8vNRmtFeeeBnBMMiKBQqJ7YC8Ow28/5ZUHuzHeA4TQTiWZCA5nPhs6Bn5icrRKNkXR3QifJK0AX74Auk2QW3A4/5y6TQ1VHXubXUvl5Lad6kxblDwpX364yWZF+FL0ajXkbkg9bWC8v09bz2aVNfyzSbyprExv6ztcsWHeLiaeI7gAn3LkKMVSVnk9D83tLQHJR9wEJieus/fpMSKoutdV3SyIYBLDLa2O+yINF6iWELPL1vkWUMuXJC3Avm8h2vhEDxxjYixBQI5FCLak8KUWY8kOd+wl6I+SHRM3nqfyqyjmhfXVRNj3NuvEomJANK6K3htVTjqjsB2WMHaK8erWPUE4teRugs0GoJfrucG3ehvjkLW9/jUKpHfQaY51es3LIrQx+JwqCY0yvKkPknUiTmtpEmCr5kejKllRLtCPQzxaV4yzVKGmEDWdMthmSLSTMbsiH5ManwXjquidXhMvdxmLx/jRAPz10QuefgPWStwgjsKA2FBrS9dCJh1V2Q14VIgWdMdnyiEiU2ZoA+lISqdwKHEUQS/yalPCC6VZdlohNuT5wnetULgTGp+oNZ5t0LvDQM4RV8QI0LkQcBCIauH/+jRK/+f+JMdDW7/5N7/HAeJ8SJFv7hnnw+ICUoO+xQMBoyKlMegS/gSl7pRL3Zt6fi4CbUnz2MbNAZoHMApkFMgucaYGMsMh6RWaBzAKZBZ6dFmD+v7at6cv1Ho8FHjL26MH4nA/P05APgR6gEep+odLPpOXiZfB2pfMCFBdyCfCweHzHo9vOJpJNWYZk2HrfPYRsai+bUFC/8fu3v/uYSIf3v+fPIVQmt4fvv+c7pPZ9A7PnzF20ZNmKz93x0Y+89Tf/158outPi1/3YLTe0i30T5gkPjOnasMGGk3rgnhmJf1+IHbK83/cWAASwQKN9tRAar3aMAtZDSNiY74w3K/wMsEE+YlcDJKxTYkWlDRFFORAWJDZbJue7WLLCXhjrxWDbMd0Fo67U5fTwNQmJoVAzJqSEJV4Yyza+EmCtDYkDQAuZgfcF7WUOI18SHf0sXiKX6lXR3hg1lGgmnIvz4/WBZ9ciaRF02IW5bfmtyHcJPYt8odjMlwB/s+373QIiLWKRFjY8mfVgAngkOowJtZNECOJ/guG7+7Skf5sQ5u8tCesTDUGZu/xOP3B9QG/Ae4gJ6UkYAoPPjHOARIutQ1b0iERgH3NEt4oQpGxvyUhkpOSlK5LB8w4oLx6WWi1tNBvwwqBcSwTaAwXz1pMI/dLbcHKFWTq232nWiLekleYQIQbUtSHYeGWcM0YtmTijyz2FvLDeWHa+YI6peV68J27FR4JWGI563bmWNJvrbvdAvd5dmu89cWhj91bCxSF/ZY4XdbFcr3hCmWugXwnongOKX5ivFWC+I8LIcR5RKkkTfUXcVPAnp6LF8s35IlFeqIs5IND9EREe2heXlJ+5C9vYsHZmPhAxQ924bpHafN75ICUvzAp2/fayJI4NbYW9IWRKkkevanbcb/woJHytfXP1vgeJDkgJ7YNkKCq13C7NubHTq5MTYqpbziqEepLbiDQcqJEAeHlslBSxrKEjGylQn9wnEr2IxPMgp2tccGoG+K+pvNCEUNL/mh/l5+Ip6hm0hgiNqtJRP6f6FUSslOQdEklnYlReF3t0/LD2iB7A+yMszM4ffdm7n1dfsPmVblDf7QWNw4XhJz7Wsf/bd+v6YUPSLJ1ntmzdrzKQ3BANpdqUnI167cC/RYRLp/yCVntznXI47Dwg36G96hWGgJgkpGbUM6fNZH5wNqE0GiJCJOqNCeRNkWhLIVGje4MShPWowmXN1/dX6T2hlJZoP4RZINuUsb3s1wGJofBZy9WmWbq4CkPqfE3l3Kv8kAIjIi/GRVrMOFxUqm9REcnwYR2PNwUaFyw4Yo5gw/Pibfoewe5jeFFYDwnt45zMMfQjyI+xVPuC9uGtTahTQmDRPqt9d/HWzI7MLJBZILNAZoFnvQUywuJZ3wUyA2QWyCzwLLUAD/x2ZTYm4GEdkOFrehAGVLjgTcfV9eD8Vh14sxIPYL+uhLbFGV4OF1x4eoCCHPvXbNh87Wc/8W88bE27kWfDlhue85EP/O1fTc3wyte+4bb5Cxcv+b23/dLP4RlxvnpsvPaG55KnOjEx/vNveds73vOnv/f2J9rCTFEWYZ/279kFSHnGdt1zn/+DJ48fPXL44P695ztX9v2z2wJt3JoFn5IV0afCPwEKQE5YUApshO8ZxxAOAIyA+9ZbAkAMEIc8gAzsJ2wDoAIAPxsgBaGWLADYTohcygUxuI0SY4w6UzfbLlsueTgv3wG82g1gE+AfYI9XAEHysp/3gI+0zbbfhsSCqGhbeW7sRB14vVTyZbJy1jODHZAe7/74Vnes2kSQGNvb0FBwpaeBjklYKCFZrlaiJ3OtOb7c3Rvlita5pc0K2dvvVwsAslvgX6Cue0SfIbdKsZBd0y+SJeyxF0dane1GBXlIlMPQ64tbQcX1x3f7nZa4S8pKloRzsCVBCM2ETwCEBCul6ZtzlVaKYFB8f3XT5Fzqt0b2mPOJITGeGiTGGuNKOuEG5DdAelI1O5Ta4V3Oo2Ri3Aga5n0cMUa7ld+GFbIaFxWFhwLQZHybTSGizgvQky8F8mOB++QnAYrWy351dy0of3ci7HpO4JbWB35ndxi6Y4HTHe5wrm1s7Nk63FZxhTaKmQOxlTgGt1PJs+Gh7FJ720wzio3bhRmvtsqpGcxn7LVfK+Z7naYvr6pgbuw3iDFVVPalOqYuV4yGiqi6saB/zYkqTXNiLCFno/1xwNg1macNOaT28QpxMXm+c72xnhf6/cVxXC/mIerF/C8iSoA5ngbJ1tSZWL3PdTeeCzo7ob0CQkPp82LVUmv8RRhUFCoKSZOimUdN8ChpYBR0dQORMXL0MR44p5PbSS+BHlHf0fu8vChC05cIVlZP7GgUNyZEhQHOq0vrvOqVsgtA+FDc5zSiBRLEbjoNTyLh8oTwDq9450Bj/vrrdHA5zpc3OEHjb0oH7v+yVxnD48PG9IPETrxVRBbI02JEZxpU/Vs6z2qVPxc2UP5DHZ48LXL9IkdkgdaQs8eXRwcuI9bVxVz3KXeN9o9nfE27IMOwcNqb9SLXO9PeJKAYXynwloYfThiEfkKvY6e+QA8FaRUCe+EJOZBqX8xXXq6HLxv25ULnZjGb8xQm6nrl2aUS9+sce6tvch7u+EByT5nplhIXEyIdPq1jCGHI66L0eH4v3Kn0Dn3/KSvIzas+08euU6L/0C/47ctxEBb0N+7RD6TXYabVyfJlFsgskFkgs0BmgWktkBEWWcfILJBZILPAs9MCPHQYgb10A+zbp8TrpWwAlGhC/M+0kBfp9fF2j41Sudzxk2/4hbfIcWGlOIPKiWNHj4yPjgyPy0sB7YleqVmvXLN2Pd4JH3r/377r61/87KdshVZefc06jn/04bOHWFq1Zt2Gjs7Orgfvu/vbUxvy2p9781sR2P7Cp/4d1/fzbhtEWAA83nLrj71i984d2z/yj3//nvaDrl67fhOfd54lPNV1z3neD2y95zt3nfdEWYbMAqcAfetNYUW1sQ1gE6Aj5IIlAoBF2G+1E3glDxoVAHJJaJAElFqmBAhBfkuCQGCwGrLiygRyAAAgAElEQVT9t+DlAvYpB6IAYNLWf6oXBfupi/WgYE4C5ATwAMhjLqGtEKh4WxCyju9oFyQH9eYcgCSAnwA2lIFd7H5AUt7PCBBN63q+l8RGQpQOHB93PvZ14UauZG4TQmiepouN+gxQKQA6OS2vivijd+C6MaE49iiZ+P6/9zPPOd/5su+/jyyQelkAKtO36dMAfuvFs/cFipGT9BnTb/AIUMz7+Gq921xwon0Lo/rhlzZPDP5duZM+bXUr7HtL6tE/Uy8GA5MypoBDqyqnT94VCkvjof+dxuQ3KDzERjr2zbkTzRfLuSV+B6fPDRa8J+wZEsNJqCiNSjmKhKFC8LiLtU+hf4zIOElgtUufZ/zy2wMbGA0AERjWG+u0cXo2oe6UuJj09nj3Q86Jzx//iYeDOLfVLRaWaDhKy6BKe8tHvGVd9ah8QOLctMuE0SMsE+GZ9B5SQWC6CQ8VCDEmtBsOLpNzFWLUcaJuYS5Lcn0SSqnNIhJYdp+I43xP4FbFLTVEhqDmIMYkjJYJBScMnNosOypQko7W/OxCYjCPSdvC2Ie5mVfmMgP7p1oe8QUSF2GqdWGJbeZYSGPbsbA/ID+EDe3Gjqz+55wVo2vR0rwMyaCQSsYa1E26EtpjiIjJjkCJaF/Yq5bQLvaT0QXRcZR0usduoklRU6ioxO/ChC+TB0RiUVMn0WrUxEiINGYt86oLb/qhKNfxO8mF0GmDymeKg48cU+5I1FxJvZlyGgq3NJpG3xtSj8vFh509CquELHigaF2dkBX4gYiv64jzzlX63BQJMxSOOsdVDvWEOEkub9rrLf+g62Uj+51mgvauMKVfmAIZHmzWMIr9hCaIxqA6nepGyCh9fVKvgzoHY48QVx1KC0VQeBIKZ2FBUdditiqHl8U61XCPznVIRezR53n125yHtA/yq1b6wKT2izXXWV9TEmKrMhDqCdLhA0poXRE+ErHuV4uk+KzyWZIUgpXfIZBQa/TdXr2yQInvubfh/cGr2TL9ivNegixDZoHMApkFMgucwwIZYZF1j8wCmQUyCzyDLUAoAFbX6dWEM1BKHiGThwk+m9WNyjM1LBMgIeCB3QA4bZiJS7EIz2fteg1nAB3/5VWv/elf+90//otznaQij4bvfvOrX3pM4g/t+dCm4PO5CItN1z/nZkiGqeGd8JZYcfWatR96/9/8ZbPZsA9f52zrxi0JYbH5huc+700S2Y4UALv9gKvXbkgJi21n6GnMnb9w0YLFS5b98/v/GgHybMssMK0FUlB7augnwBdLLgA8MZ75DMBlyQsAJ8abFZjmM2OaBNiwUYlwD2zsY+WmJQfYZ4mLK3VlmH+mhnCZei4L/NAOQEzADkhT65mBXQCwAGKsXgWrcCkXYAdiA48FiBHsZNtkV4qblcGXM/yTbQAB8fcdG3Pe9pPXxn/0oXuoIyDPjyndogSAk4/bNCw8kE8qHrR26eVhJUCq6cRNr9T1yMp9+ljAEnFPqEr3K92ay0uTV0rEyZZAm8LOr5LXBaGc0HD5nNLEQNw6LCDfgP0C+q02hJ0/uIe3ayNYABhPCQpnZf8qeVdArjEnSIkh5FgRDFpz7otsiDSshPqe8qRIqnJe01kCI9DxZj25J7Ii0kr+iPOMap8NB2XHqA3jYz04rCeG/R1jSYzznhoCo/TxD6BD0SHSwHOlNe7mmnPUtrWVsGvlydb87YuLcISTniLML8wZ3QDdSjZMF/Nsh3xOSgK0zfnFv8j/Ag5G4gZNIdZGyGFac5zIeZ27mtFolzQslshihFbCFAOaK1brmL36ZcZ5uD7QIuiDI2R9Qnm4bsz52Ah7WC0cQ0pBXMyUtDAXq028O9W6SDwkkvmG6wEpwr2AewbntfcQeeto5T6LVxIPjE7aoVeI7VmaXdFlSAJJWbr4dCqi/VphpDMNNcnHpS1NgHsIdUu4UQYhujin8PlcPNz7ugWh3/8rtnA/GHt55+g3HuzuvCvIKdBhdNJpKLRToD8cGqxnHdQJIaqK0QnnLqmWSJddQHvBWSeioiytDAXo0ueGs1xc8qAu7wGVwZwMsZ83l1g14gKkHZH6WQ0V9CbOHTe13RLpe2uMFoxIajdf7Vfqk3cF41zciTOuPjGUEkVDygYJs0j7uL/MK/gapdLkUBHrVJ7E3p3nq+636vu71FbmiAcVJsqERVSoqLNfnbb6tYWJ+qJ2EwqKBUe/mmbhd8SjIiYeTz0t6KM7TH9IFgncoPS69Ppxj2ZOm9Hv62lMlO3KLJBZILNAZoHMAqdZICMssg6RWSCzQGaBZ4gF9OBpwzhZsGGpqt6h/axmAsR7XvogARDw00qshII8OKI8DxCyqa2pPBQDgtiNZ6md59OumKGpQAY+qYSoN8uH/wHR7QfXTEaaev8LNy77eKRt2VWrVnf39BKmxmm1Ws3KxNjY4IkTx04cO3J4akgV8oiwuE7Zmrsee5SY0dNum6698Sa8IabqSrzoR15u1Du/+JlP/L+ZtIPlreu3XH+jVkZ7X/qPOz72wD3f/ubU46SpvYl27JIC+NTv0NFg30P3ffdbMzlflufZZYE0tJAFdSwwDxlhE+BZsuo1AbHsylu+B9wgDAMACmEwAJwoA3CJxByBpwVx2gEImRMsAWINfX4Q8uIviQVKqQfnte20cFX7Z9pA2Jq9Sqw255V2A9BABDBxQGawj5WdlEGbOQayArAPII4ybfgnEwpKQ3hGgM1Mm4lor/KS4mojcB47MOxJk6Cg/YTkghDaJGJipc5bZAG7pgYDbvoK0i6yc1j7IDbRyaGNgDqnrSifaT2yfM94C3DdGdP0X+4dX5T4uvpufA2eOGm/4RYkYXZP9/YYvSnAQLRRjqjPjchToyXiwvTvNg8F5gjTP9NkvTAgLBhnR4S4J8C4644k4tqp5xZhkqKgQ/u75CWBqrQ6rh4T8SiAwGCbxtFiCrGR5E+8LTzjVgS87YkCiAV+R6EFzhPPr0SAuj3ZuPfUK1a7GM8mSs95w0a5ruZAhVgKg2oc4jTh+UHsr1KoqGv+48RPfemXFt9uxc6xjbwaVD+0Q2LCIAnC1kJ+7evUcO3V0GUBB9enHiiwkBxMujXG+5U3nzOKyolJDHkh7wsTF8mVPLqTHxGt8YhcDqqajFZod7/ne7nYlY6I66wVmt7QEZAB4nMUayv2ejw3ulrlqO5GK6Sg75oS827g6mEUmJNrCWmB7Zoz0bdILlZ6yZIFLdaOnIN7Ac//9BXmUDunYXMxPYbAqOus0iIxtuda8Rttke42hBUrGb8JkQN4Regz9AVGSGqaOp+Ysyd3mPPdZyA/6B8crz4jXQd5psj6BvSOvG6/mV92vReNydElx2/dfR2172ybO/HOemHecd+dpV60UOZXj1ZrIvnNhNGYPFpUP66X8rf0d1z7vuP2KyyX6zxf5W/QGReppR3KMaCesFJGeEgB0Y4aIe6EpMEOVMu0SlSeJ6LBeqQoKtNk2+xFap/LT6O0pvJbZohYw8DtqWyRFokAvJI0L+QUYnRtJrT/gMiMUaXDqle/RDDmKf9ciDDV21efKspm3fq+rAMW6fjd2n+XyvqaiAt734xnQl6kxMWQyIl3qCaEdXqVEouGIHHGtf8wefS6W5/xyKD/8ArxxX2NvnUgLSexULZlFsgskFkgs0BmgUuwQEZYXILxskMzC2QWyCzwZFgAsF8bD4Y8GJjVX0rXKL1eCVCPsBI83K1Q4iHLCi4SPgVgk/zjKueRtpV3PKwCpLM6io0HtPNqOsygvZwbkNLqY0zqZExxDQdwdB558H6Evme8rV6/ccuux3Y8EgStswr64Q1xz7fu/OrUQp/7ghe+WFGnRs7lndF+zPKVq6/pEpsSBkHwN3/+B789XSVXr924ef+e3Y9Pp4exSYRFrVqtiMs4w/tixg3OMn5fWiD1qrArje3qaMYu4xywzIpoW48JE9tcKQnfkeQDRKIM8jL+AcwR1uYzK1ZnK9myKfPJ3gB3rDgD+E6yojsNy5K+h4xgngJYwYuCVc8kwDm8SchvyQmID+sJxj7mPfJaUgJgzICbHHelyApIC5UdHh+tuWOVZl6gEmGgVmjfVTrvImnolORFkYaOSUzuCwBuNmqDApm0AtbFuwKgJyMrnuwe+fQ5n732AHyshv6yvCtmC6G+JsHRky4dhkJdBWWqf3HfZ0zTx+g7oUiLYcJLkS8F8wGlSWYT2M94YH4w4yF9HRE6yjhjzCHWzRhLdG2iiDBF/VIlTgSC6Z/JHxVSWSkRYU8ACmtDRrHPorJ2P54atAXSws9rfXukBAZrdDEYy/K+MOGiIG3wlKIMS7xSBztnWGLv3OPF9SAktot0eZETNFfGYUAgtoVRXFx9sLFi7r8f//nhV8/9RxsizobkYjW7bCDdDSgOz4UQHYOwUOsIWzQuJynNTTFjfLnGONoC5DXa6EnEIwQKUOwueK1ofCKMWiP6WE/n+A75d4l0EpsROat00mNRnDvUinJ+s1UoBnFB84c7S0i1hMPD0YLX7Mw7tZznxkW5hdUFrFMH7M/cz2+2MYiLiyEt0j5gPUQb+j2ILWIWqeg9baIv8HstITBccz5syjHsH1Nz0bvoNYGhkt+aEBh4YaCRcYomM9fyrEQFRrN4ffLO0szqKapJl85IMnN5Kz+/O3aLK7y43uWGJ4940cT9A2Mf6Sw5j0uuxJwjRD1IPReKvinCIlDwrVCvLd0dpEyRzLPywhiVr8/3ctc4u70O56U6z4t18BLRLyWddZku5lWyyKFojwmNSp/rERcFcWAIF4Vu0ryfnE9Jvjamd9NPjRZKehOC0TZtmmxgStdMEhRkbqNwYD7sRSEPLiJ4XYiAyLNfGhaj8vZBwBxvBs6zSJZhHlimA2fre1/5Mf8iHbNAZ5dXsMNiJgiQrarIIVV0QuSFMxPSgram7f8XvUKQ8tzBwofVSp9R4r7LeOWV8/C7g8URNyqx4MCGgUyLyl4yC2QWyCyQWSCzwMVbICMsLt522ZGZBTILZBZ4sizAwyGrqW9RItTIg0o8HwF0AGLw+AP5wArM5Up2hTYPDuuVvqC0v72yhIjSQ2p7uCUeRqwo46W0izKoAw9UPH9dqibGZF1YcLhm3cbNX/rsJz9+tgpK/mL20hUrr37/e/78j9rz5HL5/Op1GzZ/62tf/jweETNp4IZrrzfB5T97x0c/fGDvE4RJOG0rFIpFPES++B93TOuxgYfFjm1b758aRmom587yzNwCWu3nPgNX9DGmLbFodSjSIBSm7cAvkBKMYcB5q09B32U1P4n8vK5TgrgEVICkYANEaRfTnrlBr0xOADdWx4LBQI4CcABOEloCzyXalYCYCeGJsDbfAc4CrNkwWMwp2AMgzRIg6brUBOAi/FPqvXLZWpKWlwK3CQC2/+i42wrjki7Ccu3Yol2kHisN0H5yj5XqCQmD15sJpq8Nm8xoLrpsDckKejpZgOufLNdPQPshwoadGW3IdDfGOvdUQiImIZYSz6NJgmJqwyAxRFqY0FHp8ZRB3wNo5D2grA3DpNX08rhgTJowToYYFB4fUkcbni6l2IBqz7do3laZHq7Tk4wOBJCv9DNct0dlcw6YPYS5T2kpJHMd56Suk2NcbTHkyzk8LbAJv2kOy8siqaM8JtSK+UHsrrh39PmHRFgQ8gd7YDfKFpkwGUaO81IGwDD14dpgH47BI4P3K0U8UGYyH3OsauVLrdmPSr5CQbEw3ohw4x+heYNrhtcG7E5nK8r3jQazF4wE/X3NKK/jfb8ZFQT4i6Hwm2P9+cEDXe7JAx3eBL+bmAOZIxOSJ6kT88WESAsb/s4QURdKYOgYwkZZnJz3gX4Pci7K51yGwFGCuLLXg3tRooeS3Ju415Af795eWSuJeUfN2qmlM7uKJda4xqd/e3pv9WK34I933LJwvPOHnqOQUP25cOjo/JO/ta934jMiiHVvxAvEeAuJpKCm9Cx8hOYIrB93WtERpUHVqK58unqiw+L4oPNdBUXLiaKarV7WK5qmpJYX1VM2eAudw/FJ5+54wlxz7kXcd6gnNaP9nIV22jHVpwYsg2OQIdIObqxgDGN2TDFH8u30mzUGIaPYeJH+hVydnDodiM7FbrW9qQ8V7dsgOnCOGVo6oZx/PJEWXfLCuFl5uI9+XV99Tcfdr9dRkRZpzqRaIjDORQJyLsbTTiWIKcJMztHvrZOp7gX38+cqvTS1Cf3zbivQfa52Zt9lFsgskFkgs0BmgZlaICMsZmqpLF9mgcwCmQWeWgsATLKqiVVvrEb+T6WvKeFlwYPmR5QA8gA6ycvDNg8QPPiSmu1xjdOmAJK0b4SIAlC7qC3V0WA11quVeFDHs+DzSpMPxhdVcHrQwsVLl3fK5WHXY9u3na0cvBr47qF7Tw/DtHDJ0uWQFocP7Nsz0zqgeUHej3/oH9433TEr11yzXqup/R3bHsR1/ozt6mvWb/zkv33oH2d6vizfxVng6UpWWMFltcriEGgp2EbyBvAD0M6GarKAOGQDgBDAPt8BygCS2DBPvDLGAREAVVghzXhjvwVXrKbNxRn18h4F+LNXCQKCNkJW0Cb2QwRCpjJX0V7qzRzH3ARgB0iErbAJ+wG7EmD1FNgKNoRtJ8H/y6lZMYWswHPCaGIExLQPUbKIFe9cAGzi/aZQUAmgy3Jcs9hWCGfQahxRHrQKEA+n/mw2TEv6MXt5tlhAnhGOPCQsPEs/2KP+8UAUBY8K514ugktaDFHah4xV6EyMczvGDeCoMlzrZTGd7drAfcgLS+y166bYOQdBbIoA0mUOQTQbiJS6SaQbCDin0DN6bIy0C0KADV0Wk09Dz+petHtdkGcSEk3XpFuXBE+Bb6IIjQGt5pd+Rhho5b4C9yTC3NSL91QKEsGGkgrS8Fe2ZNsmvExa+m6/jjkugoSQRgr40+Up1uQsJ2wt1b5OAfv8RuKYSKA/ZbeIuoQrht7zTGzm2nQlvZlD9R5XEcghfn91anyznr+gg2cZ8WyRF1EQN7lCYVxTUUaXuYUOgVwJhrSCXnO8X2oKEx8NehYPtuaVxqLZpSDyFFopdkMnV8YbIReF1UZcntPpd8/rzQ3P7nJHOsrOxHFVAHFuQ5CoYOthZ4kmEyZK6azE1XT94iz7TAistCzOZ30mLObOlUvuK0k9kt+imgb1OiHAHCKnSzkkld12dDuBkZSUeP3ZW+HkLXFKrRQzq1lY1jHYd9vNkBV8OzD6obv6Kv8heihcrnK4B0CgyGtIr/JqUcqr9BpJBAaWDzUrt0RO5PTOdYcULuqIg+vRw9q3RLVYq9e5uqJ4RSzV/uv8G5198Qlna7RLHn81c48+5e2ThMhiUx1ETjPfy/4ySpkduiXg1kPT/KJ6tbwyuB2IQ0jaa4aGXid/EKRjYyr/l95CzInS4SS3PsNJEDqqqj6Fh9SEDh+VqtoS9eEFyten1KF8noiLfn23UWdlvvj/2XsPcDuys0y3qnbtdLKy1GpJrU7uHG233ThnM06ACQ/BwPWMBxgGmwEGmGHuPHO5PNwxyQy+dxiDiWYIDuAANo44x253zq2WWt3K8aSdKtzvXVX/OaXTR7HVsqSz6mhp711xrX+Fqvq+9X//Tequ9+r3J3QdPCboT9TKQARGshhpUfGGprzO61FEBe8dJu9I1rjfvV4JzxxIjT9Wguzzi7eAt4C3gLeAt8Bps4AnLE6bKf2JvAW8BbwFnjEL8EKIjAgvGwZy8JIKoAcAxguggV8AffOoqNz9j5ErALTqgkv3wnUnUyhm2nEOwFReZreW+TvWLK4TPv/Fl1/BTPLg0Qfvp8yLLtfffMut+/ft2f3E41u3VHdYtmIlL1fB3j27TpiQueaGZz93n/Y/mmzVZVcUAbcfvv8e6uaIhYDbyEltefgB6swvS8wCJVlRINZFcjOpK+sBBSEb6Cs2m9dIBgusDZkBUANIwD4QisziB7hkH4B/m6FtUnFc5kw9282BhZVyVmuasYdxCjADrzAjCwFRAP/YBvDiJpIqQWAAmDFzk+2AH8z2xS4mAWfSKCZx48DH00lQVAuwmGdFeS0na5KkhbeWVG8AttouxgWVrEjJyhj7OHkVyf0w4xoCl/I6KRalFODaL0vWAtaGaUOQWCLvcpEW6UpJiLXzLBfe6RqKU4lRs2qoDTFuWJ/Pj0VWLLSqyUaVUlGu2SqZpwG/yc9sSRIUwCQkYJaxDnJhueatE+uh0EBiMXJCwPvc9apoKyuPQGMhNjiu9ICA8Kg5IoRyrVAYB4HOTtoJlwxJECkscmEbPEAsr/QfxguTyHNmgshQGSdbHzyoCRqKZRGFGxWLQ3PvB8t0nkt0POMmclhuKb0S7NkEAoOcGfDP+iKmw/x4CkCuANluLj/rExkiUXmailkxPQhnYuHVIjLCYZ1IM+7jpJ8196ZpvCIJm61u2goO9idWHk5XTHTDsVhaT4LUE9VvTYGl0RhKk27SWN6rN8eyoN7UoBZpNGm3o85+xblwUoHleDStPPB8BVjv4hop73OTQk7F28JV0yucWfC8NQ8UI7O4n2AXymySo2QZT5L9jiyAYM8kRZi7e5TILWrEkQAsyEvNL05mSYHMGSZdW3L7EQmEI1xW+C+JVtafWPXOF3Ybz8KrOBjufPXby6ff91gYJZIWc/dESYs50oJ6PaxzkGgTso/aTBx0ooa+j8pG7An/pxYWbRapMNDEnLpiWoQC9fvBMpEWy/V7RJm4ViJpkbwtmuHy4AvJ7QrEzVmLcZyM2dg9omORA+yqricpZqkdNaPfkAsNrcOzRpy2a/FNiATH7XGikrigY8/9ZnVJZliXcYYoiY7SYyMU+5EpzejYGR3LtfdKOuxyfW7Q+hW6I7VqNRc0fEi99lIdf6kUCl+k36tk4c/qE09s7rG8K8yUXhdWQ9nRvC5EYkyKtHAeP/qkD0DS0/44F8/V92of7zFYaer+q7eAt4C3gLfA07fAmXqpffo59WfwFvAW8BZYohYoXyRNRmShFRaL5XCiBAEzpvDMwEuD5af0svpHVamAY5m8jK1hu5hs1U9pxbXlSsB6F6vidCxrLrgQyZtg22OPAIAuuiDDdNdt3yD43xELclKsaLfbvPgfsVx0yWXPmpqcPLx/7+5CR1sLck+XKaD2P3/4g3/DFOrFLnbZlQVh8ciD9z8l4DYeHWyrnhMPkVSi5Lt3PnnaZLJOh139OU6PBSrNpJDGKBaHZSgB9Bj4ZXEnICsgLYywYH8AEbbjUYDHAaSFeVIg+0SbQ4rDZsByDG27es3TU6Djn4WyAVhwffrVwrmyjFl4VXxFCQKRPALY41WxVcl5JCgBfEBO0C8gLQBSAC1NnoTzGOnDNU1KyXk6HD+bT2sPrruQmHHX/bvPP8Q2gBtIJUCzQj4ld8FzKU/q5G6KegTUY9moBLhDOZ/pvD+tgvuDz4gFDBhH8pHxgNnMSab4C/pEuok+YMSleWTR/+lvjCsnDRBWvC5SgfzV2flcE2DaJKMwgMBmJ4WkNi2hnGSgtpwzNgEYC2aW1pML4yDIV96Gc8G5OXLhtPGqOW0bnhl9nT7i9NqhVhN5UV/pPDZSRzRAbk7pXIDolJexgfwxjkBkzEc/wI1BpIU8KR4M4sa9Iis2Bok293tITt0oIgSC96jemaUtzZ6MVY5ULK9rYL0jCCidEuAt4xS2mMlyTbQPFbhcmv69rLWyk4+NzGTjncnBeDidjgaxhoVu2mh285FmHms+/hydDUoNXB/FApuHRFqsOJyP9pM4rPWjxvDycN+TQ/F0IsZomUgs6h7ShPJjB8pv3hYOVDfiRcTFSbcNV20iLkrSwkiQqicQ9ydybsQZnifmzYunCIvagb6ljqggiLeCuMNRObE+FTGsDeK4oYjjYuRqcaZo5XUFY6/nSU8aWtkgrNXTqF6bHnnl2qnhlzuP2Vp6aHLjzp/6VGOwXfcCHBbcVfGmKOTLMo2/uRtjaY0zSvuUaB+FB0hN91VyQ9Bs7pyxozDu17o/1OcW7fFmrbtMrXhc32/S/sv1tyK+Lvhf/S8H+1SsqseJxa0gH5MqvI3nztNE+zL+t9WDIW+KqykRVFvxJsRgzLsci05zjcn19hNYqruVnAdSUXskAcU1D+r7hSIykKlarbKNocTm7pB4ngTBq5Q2K31Tq76mfb6l73g3FnVW1KvzunB2LH4jGzW3iJBwhJ4IC+ShrlGySVRMdKI9+sVbwFvAW8BbwFvgtFrAExan1Zz+ZN4C3gLeAueUBXhXAkw0wuJ6fb9WL6t3EYjxWCWpkBW81ABg8GJJ3AheqB9VercSsR2c/ERJujwt44zIZYETHNy/D6LlKUu93mhce+NzblkYv4Idt299jDwFN93yXS+qHsjv/+99H/rEe37/nb/+J+/+nd+0bcS7QELqW1/94r8cLdPs01O07b27d+LpcsRSq8Xu/toeGnHBjpGH+uMPfPzzf//Xf/7H7/qN//Ifn5Yh/MFnjQUWyD4ZBFV9tuLFH4CDdkACvAbEpi3jJWGgfzGLuNgHkA4AHACTgJaAmfQxEuQFx53JxUgCA+jt2gA0AHYGulpcDpsBDlm5VQmQEZvggQXA5WZ2lt+xB2MNAD/9iGNMloT1XMNIWSNECKh9ghDPqZvJeUvMz2Y38E6BeZlLK9blicPMeIesIFFnq0IFIRAkB6EBoMx+AHtMSKfOqHdbv1Dp/dQz6o88Jy1QkYWifZdkRMjMbUkSAWA7YiAXyCuJHdDO2rDaFv3fxgbGCpMXOyUbiLyAtKje62mzAPG2QFgUpJ0j4jL1d8kg0ZaLuBMsfW1ruKDdBLCOEMdxp+SYBaGXyynkdnabCwAG7S4juDUM0ZnSv6gtSwjwjnRehHWQ8s81XqgvFQSG9UnrS4w/SvkWbWcW+WvKy0AoQBRit6MuAvjntpWgf5WoxCZGXrCfeae42BLKdHcqHYsn02VhmkXxbMUDkt0AACAASURBVDa0oZcPXzSZjK/s5+1GKiS8LpWoTDJH2hyE0uhxoXaK+k01omhMyxIF3u5HedZXrIuhqWRsYyrvEwXgjhtxf0c77vV0AiebpwMLuSruLYWHA94O5IXEM1evjHORqlwnLclZfV4ryQsbi7kOFWWyXc5fRknRI9z9yXnMiauoTUZDjZlac0xuJFIoEtlSC8d6YV0xf5zrRTxo1MayqNag/K2gf1CERYda7YaN0UHjmrHp5e+Ycz+rd76yYybojfejuiSYGlFD+zbDQUfnUdQGXVFEjyMwikWBzmWXPBhTRhVEXvfMUB57indR2kvx0fG3kFNLFGzRNT+tbRPaZ0Kj9SaVbFhnuky+M7eGa4NvNl4SfKn/efUzbF7cdawdcL8mjgTkMzJYbMW7g/gSbf3oa9u4fmOXhCDauqo8a5y3BR4QEBU97UfM7Jgu4E6/oIu4VeWdz256cx4Yxb4DnZP7Zl/nPeCuKW9MVcIm8X7LJBfVbtSCSC5/Kym/zrFKnzeIOfq6vn9MJ+C+SxBx13Zkzh7nLOs1E4Ex53VBvDCt5z7+75RuUtpa1vmn9Enb8Iu3gLeAt4C3gLfAabWAJyxOqzn9ybwFvAW8Bc4dC0BK6GX0I8rxTysxW4rlzUqbtf7T+mS257EW7iEvUXq70usqO/6Jvn9ICWASkI4X6lOa7Ve9+KGDB1zMjbf827f/4u1f//IXvvt7fuBHXvzK737Da5939aZ+r9tdv3HT5pY8KKTENPG//+mLt/3h7/7Gf/3Cpz/xMY7B0+Ern//MP9/64pe/+lf+799+9xc+9fGPXnndjTf/m5/7pV+bnp6a/Mjf/dWfVa911XU3PZvf999z56LxKdgGCSG+ogruzJ3i8ccefRjPjB/51z/zDgJz/9BPvO1nZ6amJv/8D3//t45jU7/5HLHAAtknk88ASCo0uotkAUsBmkgAjhAQgCsWABfQ34JLQ/ixHe8D9t2khMcS+wPMAb6dyQWMxDwdKJeBQuSBbZTBwDwnfVGWkz5vHhOA9RbjwbyYAFg41iTsICFJ5okAMGIyd3Njx5kgKlzBCokbh6CW5XSgbfX6Cl8hyY8Qr5f12n+diAyBYyBILjlwVASG0DuH6Zl3jQMTlQwQOpN16a919lmAxkF7INGfXDwbxbCI5Ix3BMAuLqyVpOlqtTlmbuNtuF0xLKZEfJw0IF01g3lciLhgtZvwXW4viIqCXES9R/JHufoyCYBXYjuFPJL6saIAiKfT94ZyH5eeFgTULgkIB+fqu03ctiuUSKxliNgYJKD8Qi5KQa1rkgBSEUlB2HL9K8+LPBXjDeA5slWcRb8VqSDLNXM8Ub4k7sPkgSzVDPx8ucpYJ9bF8ZqByUWVxIWNf1zTxnfKXdhKBNP+werwjqnnrTiQrFrTjjuX1oLkqiwLN0+nYyNRlLXasbIoIqcWKWJF1hfkTpiFRECzwkAH4UyYZ504TDu1MOnmCsQ9yOLhXtpanuUiLKQbNdyfmoyzngBpDFgQWUqMTcs19ujkYUfFdwC6s0WRnHSWysB6N96cilxUSV5wPdcuyskqjGPhtsaacHd9eTieTKWKOE7b7SVh3OmEjeGd9WWjnah54XDaWTeRzq5s5INlU7X2Shmw2wz6A2kbrRd/0xIh023k/d2K4eG8C5P68EQ69NxlWeNZTsZTrhl5MvuPtYO1xsVROA6wHtXzdKad9Q6Opp0D8spIRQOlNcJek0s8OwrbjKluMlmMvI7rO/dZ6q0lW1F3h/X/DoH6j6nlfFZH3KDf65xXSNNNMniW7t6vi9YFs81/FXxt8IVgMpW/hrgn4pV0dCmRLSKP3H1hzuOkWxIWdTVh9lutWwCEdluEBAGxIZhGdT1IFVSxIDuK+2MYKKiLu+cUxS7Ziaqj0tzG8ovdGLUPdQPzeEjXiHXsfu1yWGmTvq/Wp4K5KCZ3FIzrtKTLRFgQswMnD55xdyIzpc9ZbYN04T5sBFgi0iJ98nv/uDHVn7lFXNqb1Neeq+08m5D/v1R6/GyNJWb29J/eAt4C3gLeAuemBTxhcW7Wm8+1t4C3gLfA6bIAM+L+TOlXlSAXIB5+Tgkpl99R+qySybNwTV7kkFYAVH210q8tyAjngwRh1hazwy9Ruk8vubyMzhEXp+Jx8cmPfvBvf/itP/32n/6F//TfuGaSDAbv/4v3/k/ICn4rdMWufr/X+8mf+flfhpz49je++qVq3t75f/7Sz73nbz/22R/88bf9OxLb7r79m1/7tXe87S3Eqqjuu/nSy6+AcDiwb++ibu5ITLGIQ1k0yCBeF+/7o3f/7o+97d//AsG777/7ztv/40+/5QeO5h1yuirTn+eMWsBICuADIygM4Ob5ykgKk1ABmAC8oP+Y9jP9jH0hKpilf7XSxeU6ZjKy3nTDq2TBmSxoMYO2AqaUF3dxG5ToIw8rMU5gC8YR85IAxALYAFBxwTuVDFADpDXPEtYBrNlMXvOscCil0pmQf1rMpjapdbFtAMroq99IGYv50uXuLowF6vRqFsJL02QAMYP8BuOFlfNM1qG/1tlpAQOC8TziHkSMhUQxLGgzR+Q4Q0um8MDCExLd+G1KkIJPi7CwiwjI56uDfEvywvBRzk+bJWwx93+8hOjPrKN/29hQeB1kib1b0tc5B3km9kV5+hOoiNKpQ7JQRZDvUgXIxaRIE8ZTni0YexhHGWuwG9fTXHJhyFkyqWgMO7XvZkdYpC5PjLvrVLbtFVmsY2am9LpgTCJOBPsamQMIjl36WzpXDH1r6gXLn+huuiINmy9vp/2X1eNkIko6ddETCm4ziLLBYUVn3pMPtRV6W3jwSHRQRpxU3INBR3EuHlVxdzRr/emaMipPjeWHkhWb+llr+SBvjM+kI+smk2W7m1Fndqg24+TxFJvA3VMEthPcW2JLc+Ay27EDhDDPW+STcZl1HZVhcCoeF1UjVQiM/F133jokDTwRSsmoHERWt/Nks9wQLpb7woZ+HF+kxrRxKmytnolajUaehoeidj1s1vNWLctHpw/FjUjDuqb/h0m6Ju53e019kVPGUNC+pekaXzYdpJO/qZjmj2zs1FprpDzWEQWcpGFtLM6zw8NZd0sr6x8Yzjq7J9KZ3dKiMiK4NRfWO3V1BrG8tvQCKeJfFN4gkAp7lc9t8rS4U8ds0t3r0rKWl6uFfY9a+Rr59FzQeG3wN+GrgumZ1wWpfH6IagFZRcuGlkOayWQZ5S2Dx4y7L1If9G28JU3CbWFcFCScLhBbsUqEQmiSUQtDwRyzoR65UbFVgt26Pm3gITXSderVl6qMm1VG56WMPBX20D6v1b5r9ONRSA6tO6iycI8iWYyUzuTV3xfPbrjlFXlU+0GtZwIF7Y9+hyTUY0rWL04im35XbwFvAW8BbwFvgeNbYMHUluMf4PfwFvAW8BbwFjh/LCAigfvAs5ReoHSlEjIKfLIerXkICV7MASQBHl5bJtzBFy7/Qyv+Quk+vdR2dG4AAt7yASYBYj+n9HmlaW0/FhB4VAMj03TZlVddy+eWhx+8f0beEdWdiSsh2YzskQfve0pcCfZrDw0N3/KCl75ieHR0bMtD998LkbDYxU4kaPb6DZs298WQLCYJZeck8LayWj90FGLj/GlJS68kAqRNn9o8D/hNv4FgANQDHDApJ77Tf0zOCaANQAGQAPDtCiX6HdIlHAOQz77mccE5z9Qzm/XNKmBJBfObshooxG/KQV9DEuJeJY6lDCzYg3KTOAZAFqkWQFaAHPZlvQFrVY8KBxKW+3AuCIvytM/8xyLBtsmrI000q72AqQqy4iVK/0YScFdrRrxm1TIRvchnyAzxPDuodZBSEL9fVEJDn1mpvZMJmPzMl9hf4TthAbUlLks/Yby4SImZyy+Xh8VNimNx+VNA/jBSfGehuEHw10ofUOL+dfjpelksVvYKaWH9nk/yahr+5Bnwt+jnRbwJgFkkrHhmmJKnhWJSyPOIMS0SJOu8JCrEnusoR+vX7FfJGfvRpzK5LOV5R2lWv1Ef0u90m4IDHHQwMuMGQbbz4C1BvXGL0vKg1+lq3T9o2/t0vY+LsHhaHp8rP/x4fbR2eFkz7Ax10pGNhwbjL5a3xI21KL+q1Qqf1WwlQSyHgQzFoqSTtfPD06sbO9P17e3x+qEnR9viEFq1Tl6vpZ0kCZ9QbIoHoiB9WJ4Cs1Pp8old/fUX7+uvvaGfN5bH4WByZX33HWsaTzy0or5X9wuNMURwFuqcKngBwlsqk8oMR4psV4jHy4zGIYgK7jEA5xAWjLWAzDyPubgXpxLn4rdve31DROxKXWuthjuN9fmlutY6VY+kn/JV8nhYr+ytDuJwhdaPtxSovZl1A8WpCPpN+VYQa1z6REPdGWkjKbw4glqa7t9I+kEri4NW8wVBY+RXiopXNWeT/ylIu99UU1K4lDTL8FkLxQOl/SytB8l+kRSzcqGZqmfJwaG0t2tE5MV4NntIzaIg8grBMFxa6E5qj/oj8krubMIz7qTWt7Vuk1ryDWrdL1QL2qzvyExhrUOy3Cf07b+LkrhfLbnvnoif7zwr3LJPFOLQ9dIzi8QFKIMuaZuKxX2b+/6EftvzgX2Ss564uOWy10ZVJ55TQ3hIyJAmq+j0noyvM7moI7pFkYVFF7efTK3jmGDEc/4mZWu5JMhqIiYyfe8qrgbeFVtVlxBnT+iY/eph3KOmsubwdHfdTcHBZ//k5Z2Nt74obY2tkIfFDWqA9POeHFt+L57a8XuXvevqw0cL1n2M7PlN3gLeAt4C3gLeAse1gPewOK6J/A7eAt4C3gLntQV4MdqqxAxFJGgA1PCc+CElSApmR79e6S4l9v0JpYWyNO/TuvcrEQ/jQCX+BRIvgHXITQFaIjeFx8Vfi8xg2xGkxYl4XeBVcTSSgVp6+P57yOdRl87s7My/fPIfP3y8Gt2za8eTpGPt9+T2bcwsO+YiPgXQwC/nmQVKQBvQ2oKPLgyobeSESSQBRtAHAIy2KAF5AOQJlHTAN2QFpB77ACjhoQTABCQCsMG1LBAs1nym0Xs307q8joEnXBOgDzKFPFJmEvnbpkTf47sF4mZ/k4Miz/R5JKHwpmA/kkkkWfBfR1KcSXKCjNlS1qsjJljIS5mf6liFPfAiMfJpRDPi6yIs5sgKzicSIxj0uwTI/Wf9vFOJ8QTbDDxZUbX60v1eiWNBf4K8fAhryLsiVru5XDJjDqhlKTx2JDCU5ZADNh7gxQX5RzqtS8XjgraflQSGxUigv9KPzetrvxo/IOcaF89CMj2u74ShxrNczwsh42AxF91GLqG6c48A5plECQrJp6IsC8kM5KLwL4iiYUeGQFDUG4pG0IEkEfDshir1sQzpnR36PS0Pp+VyckCm6llK12i/T5fBxtnXERwn6nFR2mBoOg1WS+7p4jhPVqV5eIUK+oPK9UYVO+4OBFMzdKqq0iwcBGlzv8J7bJ+JRg6ORgdGV0VbbxRiPlQTtB1F4ZCcaS5PiXoQ5PuRExqKpqZGa4f2HI6WHR6k8WgW1JqddGhZJx0eDSAsZELMAOhPcUVeYFHiWrCo3ThZrDHiKJRSQUUw6mIxySje/5MyzkUCcVF6kATVWB7/7VMvC8aWj0mWi5gLoeLz5LpOPq50o37frOZ5pcDuG1SpFyov0wr708zCbEi5iGPxU2Ssq+gNA3G5scgbVUo26Gfd2V7Q7QXNQStLhuIkladIrd9uDOfL25c3xoZ+Ze75Mut+PEs696SJFKRkT7V+fBCySC4X3AEj0UKrUkV8GQh1nxF5M1trPdFL6w8pwPdDo+nsfklHEVybsheEP1kqqCraIQG7N+hTnkMuMPi0tt2pOzTUQlPbLnGURlvyZ1lwndJzteek/nZqjyT/nKrgU2qpk0Fe+15HUGSzb9ZREi2jpTf/NMhnf0KeF+rCOouLdVIm4lfYuoG+Iw3Vojr1Oao8tlWUYRWJIOxSznIxLtwdvyQgjuwWC3g9IzXKQziOfsr92TUy8qDWOSpfJdr+kFiLSwZpsEKkSZN1TrZKBGPSWtafufK7R2c2v+SCZHzDuvrBx/aHYxc8ORjfsMHdoPN8e/3Ao+9f//6fwMungWwUfUnExdMiA8t26j+8BbwFvAW8BbwFnAU8YeEbgreAt4C3wBK1gEgDwIY3KBGvAfAdsoIXG+Sh0KUFlLtKCbDVyR9U7hvM2vuWEvJPzPQErMirnhP6nuoaXyjPyQyvFyrdoARAS4wMCA5cz0/J22KJVpsv9hm0wIKg2qZf7gAiJUgJCzxrs+6ZdQyQbeAEOit4HEBIsNDeAScBZdChZ9YjfQPygmcy+gLHQx7y4g+oYFITHL/Q++GZsIYRE/Rprk8ZLA/knVmpbAMsxQYQEZAPzLoEEENqA1IDkAZ7UC6OnwNpym2QNyT2k6yJZgmfJYsRF2RnkbgZlIf6oo741KTiRbJegK2Mm9gEezii55mYDX+WmM1n49QsQJ/m3ko7oV9BcjuZw6cs87JjeGGh8c/+k/LU6D7TJFhJYLg2LeDeZunzmzGC8Q5glDbOmGD9nm3Kq7zRsoHWaXp9ngsA16OHCD2FcdAmdZGjERRHswHrpQ/kNvdlqixTDAAJ9TA3nUAZ6YBp/AolISg2JWsE8naSe8jsQQpjN/McySuBxx1hegwCg7GZ5xc8TG9O8+gyTae/SGXZlCtAdqrJ/3mqSfNZPjmIwn3KwG5hwA+IO7g9jpKHl9f3LIvy9CU69s0aV1alAt4dORsyyz68VOOOYln09y6L9++aSiceY2MvbS7r583x2WxYbiFwHIqOYXapOKtUJIQE7SvIcuLuI+bpxyHmzcZ36ohPRzwhFaVP83Cbs/rQ2BDBtPEAvEwJcB8yRJEc8ufLoi+pt2qXijwYTvoKrB1DSiGUScx4IfLKEPJGChTeUVyL/iCv9dNBdlD826wq58BYNvtgK0gugDQYhPFj9WBDZ6T+o3j6bi7q9Z5OffIvnwwH+3VjEHGT5yNqKi25kkS6BIyD42pcPPbC0yRI4vraw+HIsPw5lq8OottXJlNPQPmVZZ2fAlAYkP+Xl61AvhGy10D2UEwLWeIRjdw893KfZj/G+hcrcf/GTsS/wE8jUySXJPusnnUflQwUfj2V51lFF8kkJ4VtcZLolV4WVeyF/gEtIr7C9X/ntakML9MtRWV29bRKqlnumF5RTPFBxVUck1jWFt+PMYuBet6GR4U+u7roTeqFwwXF4E4gYiy4qp8FI7Lrg8no2m1Tl75yfLD6WbTX4XhqZxx1DjaSsQskV+kI00fErtw2dvcHDjR33TOkayOB5SY5iLjgWq7M5FIEhl+8BbwFvAW8BbwFTtkCnrA4ZdP5A70FvAW8Bc5dC5RSUGjl/7LSc5QAHfGqACwhMSuYF14IBwJXW8BgvBN4zWE2NfIuvGy5F92FHhJlcEZeWrYq/b7St5V+VImXaKSlflzp15XuUPKkxbnbnM67nJeANeUCAyCZ/FM1kDaEHr8tPovFJmB/ZnRa/AY8jPCkQJ6DBcAMTe1NSkg+mUSE4Q0lyHcEOWExHYw0eSZtbl4SkJKAD4CQ5JO+jsfUo0oAEoD15PlxJcoOMmiyI+Y9YSBYlWjhu2130iRleibLdELnrpATxxqPqAPqfoXaCSSNk4KypZSFEqrmFurNNOQBeb3W9wnVxNLZCS8LLUiNmdfCpNoNwZiLWdWlzJib1FwOCVo3qt/0Se7bJhd3Ju+heCW4ShLYb7Anfb+QagoV7LqQhgJWpb8kWk/7L+LxZCklU7iDlH0Ex5aOGg5b1iGQGSy4ErCYp8VC7wtH4DjEtS4sH68GXA6K34HkkQh83O8ilsQM/eX6vFb4NbJbX9dvPA/MQ4QyzMXLKQmMuTKW5eR56GId/0qd5xWqm4tEN6xxXiSNtsogHaB+fyAXgscGWe1BRYJ+SDEanqyF6UPyTXho49DW3StqewCgscMGAf3P1TlWU78iOEY0YAggD3eqlvc2o+5eeWFI7iiZ0HT8vB72Z9HTUlyLhmJZCPhWgVzbALAvTFQaqopaN7SN8Qn7D2t/xm/aGL9d0HCaVlnucX2hbpLf/dYbO5xWklMCpoON2ulq7flsUSWbtK4pYuKQiAeR7eHFtXo0UmNaPspccRglQtRFwiAFtkflOkRcBB3ziOKxg7UrVoXkqvJ8qqGyjUu6qZ0NlmVhuCKP18+sHP2lH67FGwqyQsvQ4T/7anv2wR39UHE9wiF51ATr5aSxJo2iMfFCoQzQVPZbukYsMSZ4EqizOM1ryzq1Zm1vOJH2wvrQsmz6ieGsN7PQUu4i+I7Mo/zYpa3fyqMIi0yEYKh4MWKJtJ579vOVtmrbk3hYuN5ZeErMal2Pp9ycp2U6qVq2LJ+Hmu5zeEyU2WtkEelXKaAJYk+FOFVB9FEP9JueqpHA6XJ00P1E5IXKpfIFQ/rdER8jeS15zDg2TjwQRIm776jVKRfOBcO1B1VghcSqeluU12Eygfw2nEKXPIIKCTcdT8hyZKvUjhuxRLzEieT9oNZox/2prL3zjj3h7MHp7gU3NfNl9Q1qsKvbj3/lQyu+/j8J6E0ckEO6bL8YsVyZaOOOtKh4XljV+k9vAW8BbwFvAW+BE7aAJyxO2FR+R28BbwFvgfPKArycvkIJGRoWXmaRoeGFpot3hD55oSftLAmO6gSuI2aSLWaZCoHBvrt0jr/XJ7MciZPBqx2kxXuV/qvSp8vA3O71+0Tkoc6r2vCFOSssUBIVBiYYsGAkhX1CRNgsYtqrzTYGDOI3+4HmQfIxM5UglcxSNS8DwA9iVtAX2J84LAbmWR8zbwvXHZQgRTi/zfg8GXtVIa2FfdjOXz2feQUAtENWQFzwHTmnryuxHVCCfJPYzuxQm8lK3stAu3PBt23WpU0EZd9CXRzPrIXSLydTujO4bxm/wgGAStJtDy/SZ1thc+ZyUZYll0QU5cM+jKHmSXLWeJGcQbP5S52YBehXjAP0JbWbfFpA9pDa05yevRFjWqUZ3zltj3u2Iyxom8+0l4UVo+JtYatKpkFjQxQZuUq+9N2Rdr2SxHDuDgI8hcWLrGCcDKO2fJRikRSMTUK8pdov9F7fBfsKOnfDXzmEOW+EcggzcsPMg3RWT10O1DaqJdLPUr+TTNWgN63fI/LqGAmS5Fod/ybXH/OcmDuMVQQTx+700RL6BXbOstYHUOnSHPnQeYbgnfEcfX9lkZAnKhklSVWKfxFRE2wXiP5VZftrWRbfoxgWeybqB/b+4sZfLT1mwJuDe5XFfxYRwDlfJpeJus4EGcL5L9Ip98mH4rC8KnpJFncFzXfq0WBaxEfSTZvNWGpKcaSWUZiE4aY6pjv+JtXU/GI2f8h9iAkiEKwiEFzcJbUvZ0T8H6gb2td6nY/7URDG4aQ2ptpXQaCjKwVmXyfTSkorWBE34ZZCF3hBYkvZoCvsPFeYhTRPAvFCkiuDlH9MSd664VaVbZt0sbDzQNltqXqiep5NrQ4mJzf3d0fXdLdmg3h966H173zVIN7wIlciLfXB499aNfPVTy7rPXFQ6PqhA/FYJPLhql5Qv6IfxGsGEpjSqSaE2q8Wn9BGiirIIoHwIsFw1VNQ7umoffWgHo8Nkri1Jjj0iAJ0qx3YFfSJ/apUOfB6oVKGqBPlgJi/RHepca2n3V6kdKu2SZYr+LK+A9CrXRf1oHPVXe/lvobMlEK+55/VntRyTy26iNvmxv/Oj4h4wHelCM5tLQnSn3uLono4UoHGT331RVCovap+RDRof2zZVxpWog/BV6hJKJeu2udyVBQWAsOKrWO1fYcyIQIxOKzvz9I2SAcxbiJL4mA8y/px/fCT6fgDH36we+CRXUl7Rd7afdfBwaorRpWldpj0uo19D9297iM/Ox33Dj9LV53UORpqEod1cSPE7NmJKzvvHREXNkYEPt5FpR36r94C3gLeAt4Cx7SAJyx8A/EW8BbwFlhiFijJB9zdeXFH3oVZVn+jhMY6sg5VgNNZB6knHcd6gErSnGb2SZALvLj8kdJtSoC4AHm8pP8HpRuV8N7g5dbPQl5ibfIsK64RE6YTbx4QNgvXaT8rsZ5+QHuFhAC6YJ0RGhfpO4TFJiUAKSMlAI9Mp5tjAPcBwKsv+ZikCkSRJwtwewRA9QzYzoEmSjb7GNAdbX1ITdYDbAGqsg4ig+2MG5QPUMJksrCXxd0wELOqYGFlrCCSz0BpTv8pjZAR6RS+QvjYkAIkV65SFEd8BZ4njK9GzjD++cVb4GgWMNlFtiNZdJekxq4Wmjku7Lw4xgIV1BtXJ4Me4wVxpgoS4Du0WKwLeSXYc4MBsxafhrGBxJjJeMB6wbUhhK7GkVyxBBT3IEvZTh/RDH3JORVeGoV0UUXv6MhiLlJsh8U7PSLGq8dEoCguQIQkHxsYu/6Vu4YbkxWBIFDsiyJ+iD3TFOOsYjWU+yO9hTfLeq17lmagXxw0WwKHVcyBipJIkyrpPq45918T5CuZy/wRXe8Rbd8j4iE50F9JvRpRC3GxR1n8Z4H7o+JaLq01apcQ76HXSYYFUV8jgF95zDcpAk4yyBvjSVZfl2W1sVo4SIeyyQPtqDYtFxXyyrmwGeP0YvXv7kcEgtbF26ImFCQ7n9V4BfjNIhmtQJ4V4QqxHyu180qtXkHYFK3viBGYjerhBXGjtlockkgBmbQvhS0VWV4UPR3XSQeO8LhH53uIIU/rHtex3Be2KEFwK66FJsBQfnkPpAqZLUYra4RpKrKC/NUeX/sHzbR5DbJh1MVYmPceXnH4L9852n/QeQPI0J2JdFqxyWsHkzTaIgmuCZEXcSdsbOo34sv69Vg2iseStDY2CGqr1W7wLAHGbyZRY9P+oLayGQw6Q1nvYZiyI9vPAsuVJJCjHyAtMudN0XRyUUS6qAXPU0lWaz0SUcQl2qZksVxsQgL3RmwMbZFBwcmHaJB/Vd9Wqob1gT1PfwAAIABJREFURND+qyA/rKDd9cvU3nU3KT1dyBoElMkp0a9pi9xjsRXX4TnC7qWSb3IL4UxGiGOuvVrKxDAOSpTUeVtoB+uY1kj0SXvnOuT1ZqULlcea6pzMtKNgcHneHUy0H/+avKjDe7prrq7vfeEv3po1htutPfc9Mnr3B+6LD21frjgbSGplEl5DDAtbQaBC9hj5Yu8L5JnF5V3khSujl4sqreI/vAW8BbwFvAWOagFPWPjG4S3gLeAtsIQsUJIVzPYmlgSkASDjJ5X+gZeXSsDsxawCQIJ+MyDsfUrMQIPIOBmPCF6JvqlEvAyAi19UukQJcIJlrdJnlDxpsYTa5dlQ1HL2Mu/0FjfCgmoDRDjZBiUABEAiA4r4RBrJcAFABkA2YlPcoiTpDDcLknNBDNLO+W6gPkWvxqg4milsHwP3DQA7FlDJPgaSH01Kin0AvsgP+wAoAGbsLMvEOsA9frMNoIZzouUNIA+Iwm9LBqZgK0ALk4ZwoN0i8SCeQo4ezQBnyXrqGxtsJNXqdcmTCJVyM5ptqq2T7pFoS9bXOuxCm7H6O9fKe5aYfUllw82apv9oTJKy0DzgaPJQClIAcMmkg4uUiIFDn8Ub6jt236x4XRCgm3ZOXmj/5l1Fns2jweTjeIJQLADNQc+ycgwJBdBK/AdpHZGBEryBvGD4KFDYIzWQjmwYc55a7OvAaQXeDiXOo4DbuaD4Wsz11+r3C/U5pPn+j2nHA3IXmC6lrGZ0GWSqNmreu4jlfKW+X6x1I9ouYsV5WegZRbeIPOX8j2vdffp+r2STvqIy3KEg34eCkdHJ7msac+D4O4pc5mWQa0DiHcrdZzU+tHTuF4sAuEIlXFNrhEODXnCxfE1GhhudQ/uSbLSfNRXDoD8cNeq9OK4dkvpRT+0AW5UgMOpIDtB2Y4y+y+uhsJe+05aW6XMkjHLJJ4UEI9fYpENyEUZRiAzQuCJ1i3QVUB0J7FbABCjWPHLSXgQHx5tCcSLkQ5Hm+2XZ7Tr7IY1wIpbU5nJJeuaSBw1FTIThAX3u0+fht1/3Ier9WEv+7e2TulguAin8A9sxTvf+9tjMZ74ZZzgRFPekWEWKXawTRwQMaap/YzZqTnb6zYO9vD6c5LXlkuG6YCoeSvpBfV3cjJqyLwJLDfkkNCbz4UubquOV2SSTcoqlgt7Prasi+5I50vp7db2GWnJxH69rLO9rAkKkeBbKg9Y1ZAMS9AR/3Es5Dpko5Ka4/8062qIIfR26iT8K4hG8yAXqrpJ8wX6pw41IhAqVMO1t/YbA4dxLIS6KOi4yDOHkJlNo/1kdUJP/TiSvkyEF/RjXLWlC6+viwpxSGq2VQBokbEo+aSvkU82lI3tt0v60AfpeW/tpfFFLqcXd6ctfFWZxq97e/g3FrpB+2favHJCPS5Pzkhk90LTluhHr1EiL8byAnRmT6AP2TGDyjxzl+oaICxb37OTJi6JS/eIt4C3gLeAtcKQFPGHhW4S3gLeAt8DSsgCAKe/PL1MCeGM21F8qffs4ZIVZCSkbgFikBgAteTk7oaUqEaWXNl7A/orrKr1OiRccznWrUl/bP6/Pp8TFqF5IL7vMaod4efjGDWMAqn7xFjhpC1RkoMABjLAwQsDAQ87LC7fNuqX9W5wKgDiACl7MISsuUrpeCa10wGoDrozoYL9jEQ3VMhigUYhVFMnOt9AjY2HZ2Y88G5hlx7Ie4IP1AF8AC5Ao9CdAEYhIAXkuqC/9lNnelM9mkDKLEs8B+izHm92qwAT7W8yGhXEsFubzrP9dSkHxzEy9E38EsHg4FTwmVGyOrHCAcllTZfyKORmMs76QPoNnkwUc0FcQfMVQYWQF31MQ5GKhj9IemY3eUzudPlOyUMcyViVoNQG6DbQ0YpR+ZGOCAHRJRmWZCIO0iAEURfpUuZEvCsNl+kp8ZaI4Y4SSFawMn1UCY46w0Ha3i0D1XLbJdf5I41sN+FbnGKQilCX1VIux36RcBriGyJFQYKuLuXEZM/VFljDzXxMq3HUHkpbSGK58dGe60kZiHPy8zv1ZrX9QvgxbVG7G0qMu77j+7xmDUxEXHWXlNmalS+dpi4rwehEAL06SbCyu1+pxI1gzVuutqffSoNtv5c2oJw8UeUGEWQd3E2WmrZEG4sPFstBCuQSgi5bInW1l6zCWY448Q3LI1eUKxC1vi0iz8vMmJlPSvSpv1+qK0K0hLBE/IO+OXN4UeU1T56M4aqdJOpidTIDaJ3XV/SJL5KUgWUDJIkkGj3vFDrXL7br6nl+44SMnRZYVZAX3yPA9FYPtzcKRb8bpnl0lGG/xWSil2oOTW4IoGB3Ke7Nid7apVoD3V0zWh69RsdLp+pBm/DcuVNnjUJpc2EjkxuaDtZHp0bxzoJkPaIfFfbVKH9tdjPWFTwz7PaTrOc8FpfXu6ng5RMGVuhvOOGElR3A5jwyOgvDiGQCbQVjwTMs+EoUqny0gKfra9zNiYQqv5dxNY6BFMqXhm3Ip+dGgn8nFRvXiCA+RltQ15aYvkQfu11yDazXVBhSjw93rFTdb8kxZcIHql+s3lalYvUkeQxJeK/Jg/5EvvIvuhvDQcRL70n1NklgiN0I1gbq8NtalLfEe9eG98cze6cHEhuXj3/7LOxp77sM7OuiWw5ALHyLii8R3BSxZpvNs1y6HqTNW6TvXoo3Yc4TdG934UJGM8uQFxvWLt4C3gLeAt4CzgCcsfEPwFvAW8BZYIhbQyxEvCswsfLESL3IQDn+s9E2RCSfyssmLBZ4VEAyAsduUIBaCk/SyMItzvnuUkBCAPPkBJSKQ4vmBpADnX3TRyy4vXnh68JLY0O+mSItCQdgv3gInYIFKYG3zqDCvBwsITRuDcAA0gWwATkBSxCRCeIayF3GAB/aD0HiBEkQaREZVNdtytdi64+XYyIrj7VfdbkSFERv0N0AmwAb6G+UFCNmqBHHJNcx7grgUSHpgC8YJjmMBVGRfCEI+S232Oekn9jeigutZmgP1T6YAZ9G+2BJCh/pH0ouyY5enLCFT4hVJVu2L8QvZEGR7ADKPN+P4LCquz8p3wALcywAh8VyirTHeXBnF9RWZvHiOXBzuSN8zTyjaJTOb6X9zco3fgTI85ZIleTEog3MzNjBuWrBhCkaMCMZO+hWfLPQVvmumOhEACNLtxpi2JJksdoT6Ga4AZdyKo8bByQGNAZ6vDOrymui6bggRcaHEaUoPMsWogLwIIwV3TjShX+dURGmREvo+KO4LoUImN5WlzuxA6/Cq+JBWfkXr6d+HVIa+yugk8FTmp0oPVSwj4iITacE+u+Wd9UkdS71hi8s1Cl8soHosSrua+q6Y4Vkz2NtfE7fi2RVra4licaSrFeB6t8YZxboIJBfm4lIA2xNPYlhpXKbYVoLTPCMNK/B1Q8WpJ/0Meaiw3lCgkUQ+FMy4FyoNQVHERxeVk+SH5TUmJlaEDeNWzrNYyHMfYx4kDbKdeFHQzjDmzH+44cMn8vw4Z4Hy+Q2i7d9WzMLXf53WJu5pDB437xw+7f5FezevR+rUgG9Y42VDWXf2gjyZnMx72/bG49dKMup6lXpEZRarU1s2U2tt2heM712RTm5tZX36WXHHq3BfR+SlWM/1IfAhLS4o94WeGFXarESf2+eoAfaXYhbkib5jG85OX+Z+a88W7EV+rT0XoP20znTbfIyH9vtk+B8K8lYrUIzxOQ8Fe27g0+QauV9bnyG/to3YGHu5luo4kjTUiC60Qhcdbqqq7amkX3QdaBgmH9xOXtQcNsmnSZE3ZJpa3EgnLrxw/3f9/EVEYa/N7t+/cvLJr0SDjnZz3jxzMygoEO2p1D/jWuSx8DYpxirGM4hViAu8Uo20JN8cRluyWE9VKontfvEW8BbwFvAWWKIW8ITFEq14X2xvAW+BpWWBUgpqs0qNfjOSTLx48jL1aZEVgJYnugDC8dIBsQAoS/DBk3pZXeRCvKgAvADqAYwWs9OOvRQz3QqJnVcpEf8CkNUv3gInaoE5aYKyvfHizzoXJLJsW7xkM6sewMFICcgLpEHYFwAOoA1QApDxOiVAItYdbTkaRLJwfyMpeJnnWuZlwfGWqscsfMlnH9O35zt5fUKJfn9xWS76GmAF/boAcYqy0Bf5bedgnUlUMF6Y5nsxK3o+b3wfLCL9dAxznDObIK/MnqMiJDRbWVVSqU0mgivewEDb8EoxW2NfQJpUs9/PmcL6jJ5xC9B/AewAGumjpCeyJAHcG1bbOmLcUBtTAF4XB4I2ydjA/fB4980zXii7YAniIxfFeGaAdOF1URAW3PspC++m6Blp/jpeA24WuYHTQyILNKNdrCDbmG3faBehCQi6TVrocRG68exBJ+mUJBfhVRDUBdtm6ZgIDwJ7d+VioPgE8Zg+BdTqUmjd4CrlziWzp4OO8nNQIygeGKqf/C6t+5Jy+ZBIDcbJpvYlj4yReJVQxjnvqkWClAciLTDNQMTFTnkrfFGOJIwRl6ten9/vZs+Lkt76ethXiWJFcBirt/rd+pr6rvpQNNms5/22rr1KXhe0i5q8J1JJNnFNPAFGlP0RPHJkltUylWJn03oootwAhF6LpOiL6Ej1qZAQYinYN5e9w3BavMUeHSvPFFd2PeuFAPZ4ViAHxXPa4/re4bqUkaDwKkNN5VnIqh2rrQFmM0Hlxyo78QynGCC6f7zCTYIpse+5ex0Zop1zzyniSxU9wkkNSTJqJM7ShiJv7zoctndO1tsjeVq7TA1pKBbWLh2t1QfCkauaeX+ylfY7TvjIon9YbVVzPN/baJfbtPcjytEGHTfkvCVSB8Cv07d1Wuc8Ccozxvpd+H240NmuPUuaTM/ZhUQUVzaJxmKdkz8L6qKuCJ2d6YkjDZ99hPnmiH95IpAzI8Q4n8k5ck68JKAk+O76mPOmEamkxO9RRexu1uTHJIelBpJhiqPOCWcU6v7xohkEe9XoNmjlqqDeau590a/URVboUDW4L7zzrvaTtzvGzwiLai4LJyhHZDTVo5AiU+wTF6O9eHZwMVOcx6bFYCH/rs+UdetOqzKSV767cnq5qCPagv/hLeAt4C2wpCzgCYslVd2+sN4C3gJL2AK81CDlhPcCM6fvUvqq0qKzhI9hJ14uAOIgPiSV4MDZ+0/WrosE6sY9HmmqTymRV8CaYy3cv56nhNwBgISBrSebFb//eW4BgS82M9HFUCg9K9zLvZJJGvGbNmWzfzmGWctoV0NE8PIMUG/7AyICsrE/QCH9CPDw+UoW08Ise6IExcKasBd2Xt65joGRi5EVHFv1wlh4TV786SMQlTZblvJxDNIN9GkAMxb2ozwQgJSRuDKUne30taoXhYGPBqJg44XlOB9+UyjaBGPTuNrQFSrnhiLuCShPEcNC0KDAwBQtd0A+iF1mmAJ49c4GqZ7zoSLO1zKUZFYiWSdmbQPqkbalyeACtSeAaeHrQkDdpyIAF0Gpr1Lb26Xv9GsDQc9qE5UeF4lAfcYRI1JtRjp5Z6xj3FG8AhcGmIDXDZEIfCdQtmIGpAS9ljQPHhHpsIwh4gFweFHJKJ5ZHpfRxgV/KnpAtjYI06aOFbAbjYh4IOC3/BMGgpkd5Ko7Q1O/hewnXQyOsXfquIeCrMez0y5JQD0ic9O/7T4Bic0Y6fp6WQYGBxdcGFmsxUgLClsSF46gEvC/Ull5JE/SQ7r+i8WnjPTyZms6HRtPO/VwSJzGymW766ONg6sZepIEwkHZbSgkN4ESpOUD96KSrcMpJRVjod/iUGXIjvgIDU9a1UkySJegV8rXCed3A1lPFpwUNr1H+xyWLQV2h5NqW7THus7B/VLUhyszJJLJHTrZImSu9OmA5hcv//OntEF5wAbyrGA9dc7xP1XZiXP8X0p4cbilfEZ0gDUevKzSOic7qN92TyQvdg8C/N9RD5LBqnTynifrKwTOS2CrFlyRRDJTXd4Wg2jzcDT04Hg4u6OeJ8VEm3mppiM9Lubpf2iH3TLvHdpb7VDPnE4HEJJKoL48YlTLW/VJ/A7xS/qT/FZJV+FFwvMD8Sb2aB/6NGU1cpF6OKizsc7krxLdNXqOsCkpr/DV85YSeJ9334pc3FyMKHtusWcYIwOYNEF9YW8ko1jfLiWj6njiqJ0QaN3kog5r3aT23qY4GFeIpLh+dv0t6ztrrnXPHfH0nnz0/o+sDQfdVdrPTVRQbys7XJE/06uC7pM0VF1NsS4ihLp2hIvyQLu1mFg0BgWBd+eyGGElQzhHuBhpdUyPpXnr+G/eAt4C3gLeAuebBTxhcb7VqC+Pt4C3gLfA4hYAdOQFk5cEwEhkDLaWL4AnYzNeHD6h9CYlCJDHOI/S05ahKGNoALycyGIzSrmPISll0jQncqzfZ4lYoCQr5oD+MrA2oDPgSyGlMT8T1gA0+gmkA8HpiVXAb5O/YH/OBxhwkRKzLAEfLPFybnINvGwDFjydWc8cTz6NdDmZmqOvAphzPGU2Uo/1Xyz7jHmVsM0kngAUSC6gZ3kOtjF2mP43ZTtCvuE8JSrM3tQhZYYghax9nsiJVUXc3fklrtWDfupWmqeYBR32Ehcn03KX8L4iLlKRFhbE3oF6EVPjAdKRQNKS40lQjEE3KzH2MOa4OE7EWzkXyDEA/DI4t3m0GRFrhKhmZDupJEhSCAHGYRb272obY5YEc+SBEkriLssZs+U9od3wkJDLgRB9jAXUrRnvGc8qHKN90xX6vdIF0Y4iyT5BWCggTVwXkaGuniSTuErpOMY4CIqHFNTh8SAl0ENmnqCM9YyrEEdI7AFG08/ZbqQL1wOMxuuC8hkJvSiBQdBq3aM+rxDTD+7sb/zElu4V372/v/bVs+HEeEcxyfcmh4O0MeqcPQaSOqo3ayEkVnd2IHpC0cmlliXlniDppyIfFNF7pN7ozSZZloj4oQVBRAQhpAteX3iKAMZDtJNH4i/MqmkRc8C1PxEaNDTIIMjtIYHLRvJTDuqjIDrmnyuxV/L5Az9OPaVIX/HFlpK0AMBXxAbn5WfLG/QF+bxFgemSvKiOoSahZSQdeQD8Z9ztDmfdTjsfvF+xK+JOVF+ZRTUFTyeoRz9tZ/3aeDRTW5FN7VPpILMA7CdEF8SudOTARA3nuXfInO3ab5kjvSLFs4h0ROrIfOST8GzhmXqPoxnmfU2gLhTcXO0yceQG92OILXtOYFIAZBWf5kXJ0XYGRQt5qgdz671zkxMyeSOYnJKR6tiEa5hsFvd4EusoHbarqS6dh4juVrRf6pI02gjVR1SWqTXXDT/x/X9xYdYsnEWX3fG/g3hmz2bFsj+sC3Ee2jt9c67OzFxUlOg+ItGQUaYwSHRMCmeytZL71DqeKbA07YF+wvgF0U/bK7ysymcnldEFmYescZnxi7eAt4C3gLfAkrGAJyyWTFX7gnoLeAssVQuUclDMUgR0fUDpa0pfOQWywkzIjGxeLl6k9KASmv6sO5MvE7zwMVOclyxecvwMrKXawCvlrsSlMHCIrdUXeSAJIxdM+5kXfvqGkRI8G9G+eJG2WYvIQpEAztYrAbZcVK7jnAamcT0AASM/ni5Zwfk4h2EBx3JfWLgP5dlW9g1AKfon4ARABePAViUABxAJi8cBCGHBMSkvABS/AT84X3XGIyDC+epRgd3dIgCY+qXeKe8KtbFbpIKyXsnF1WZuciSQE1UPBUPeqZWMiYBvjEuAlwMvBTVnTv/lxCwAuIjX031qTyNZmhBkYGOtFrfxroB4lYNAjSDK2ucqefWw798qOSJfbbarNnfW3xMrXgd5SV5UxzdkmBizADMhBso+KPko5HcKDwx0m5DYAY5X/wzH5Cmh2e2hQGgko+R5Eav7OqJHQaKJhxGEAKUCnkVYhOFefTImMv5hWHlvyMsizzQO5gJu5V2Q5/vlmrAjiOMZ577Qm0VGijGUQN3kD6+PMeVhXGsIfM35KAfjBv0f8hdg1uBwR2Ka14U+A7PD26/7kJHMh5Z9eMfOoWByXScfef6g1pYE4VBtV3dd59DsyKGVrbyRJVlbrh/71Ba68pBwHnh5P6srmHekJrJHk98HSS+lfYSKeZFquEJf6pB4GAH74V6hyMyoJ/+M7X39lmpSCZS7WqB4rrEyR59o5SMiMNbC/+iayP45gknHSBZqDoTn/kF9OTkieV2YjKB7NpTnBfnk/vnr7szF8r+UviAy44QlpfTsyvnyMmi1yUSZ9+NAgbUHz5+9/+73j73gkl7UfGEax+NxHDWztBvH4XLFY4gOSCNq61gys0+BPAjm3S8DaENeEJ+ipRZBuyqWwk70yS36xvPDat2VG/qOPBQeFVA7dZ1HbUz3SfMTIGd4Y8Q6X+KIDdpGT2t4XuC+Pqx1RewrvDMKySiuU0imYeFVcx4leTmpp2I6J5fkbFGuJHg1x2J37tfkgPNzPWwPGUUMDZZpHTSr+lMA96CtOqR/rRTRMB7Gre6B57w1FVkRKV5FvupffjNbcfdf1eJs0FJvu0SHx2oGj6inPKHjpxfGuneZ0X80ZmcCHVB2bD5Eq7kA3fSHRPuMaNe+s4Ocx7SDI2mV6KeUw6w5oGyetDii+v0PbwFvAW+B894CnrA476vYF9BbwFtgqVuAlzu92D0mO1iA3Tu07qQDVFdknHDJJw7GW5QgK5gtx4y9E37hfDp1IlkB3oGIFcBMQQDX6gvb0zm1P/YctkBF6sm8EUwHmfZhcj4ABiTICIB6vlugadqwk79QApRgH5t9yAxTgJbNSsymZTuAvnlTVC3HSzbXtngHx7PqQqKvSjwci6Contde6o2ooUy8+FMmXv6ZfQzIhh0oN2VgG0An4wJgBQAK4JV5VwB4cCx9zM0SVrK+JkkKB9ad14uAX+zlZp4qYVMhOLUNYHWS6mESswgbh8WgC5WkWfZtrfuSfiOTh+cXM2fPyLh4XlfE0iscfZJ7Ngt98KCA5u8O4tomfQf+czPrQYsbraGRfjqLJxj9l3EJgNJAy3PGciVo78aU0hsBvBPClEQfY1xibDWCQUCziIm52d5hIcmUpZAVRZ+t1dRviY+BeA39UPsUwaIZG3dpP4GkIX1bQZV1rozg3kQ4z7WP3Bi4pkwtl4VEiayh/ca4zgQQxv9Sjkf7hG6MEDEsTw+uBQAdhOSDmf/kjXphLKA+KSeByN05S7Jmrq6wRScdmuoF9cc1nuzLs3ijRI2GDg0mOo9PX/i1C+MHJLmTrUiS9F5t74i8Wg7ZoLgU9WSQ1vMs3KkCd8W90B5WKOC2ZtSH01GY9cTKmGSQcz0pbeog+Xk1v+K2U4QEochqXLEb8N09U6uQ8sEgzNSP9ZuxUffLXONdeLCU+bH7hyMwhmvrFdC5e2UtbP2efr+0LCyEzp8onZKHbElcOI8EPZOSB6SkCrz800FvMmo/nIT125T5tfVauC6Lsvah+tgN/bipsOrR3ZcGOx5bkU5RDrmu6D4H6RAEF+oMa3WnHClpANqO3et2qV6JH3KJrqYg7c7bQnFU9GzQdfcJgrsTr6IgCx1PRk27X8hIQSCNzE0/KKJoANTzHE3cCxoE7YXrGbGAbbj/8tztPA2sjKUNj/ioEBh4X1CR5oFhHpPmwaFwFngqFTKY2rGt74eU3dVJY3x1d+31rsyNfQ/tHr7/Y1E0vX+l/JDCOA5WyV+HtmwyTpSwU5Jfc4aqkBRzZnDkfkFe4DPmXDd6Ohr5KDEV9KsWBIg+kdfaov1oH5TfvEwjvC1UxrOejF2sbvw6bwFvAW8Bb4GTt4AnLE7eZv4IbwFvAW+Bc84CesE5oJcdXoaYpXU6gMZvlUZ4jT6/ofS5M2gU7l2XKwEGfl1ph2bnnY4yncEi+Es9AxawWa28+LLYTE/aBi+4AHoA84AGgE0EzjbPI7YjlWYBPdmHNgYxxgszx12kBLAACMS1juY9YXJTJ6Mpz/UL+Y1Tk5AywoJycx6kMQDcqt4TW8t1aK+zPzaAuAAANIkHC4LJeQAITfqJ/Y2wAKhn+1JY3IxQJcgr2oSCrD617JLJoN1A/hhRgQca9iugKr94C5ycBczrC8BuqxL3vEvkSUE7pN/Ojz3FnY+2aRI7TgrmXJGGOopZbLwxWT124zuzrosg1wX5CkjM+MWYzDjNGI5rAJ0U4mKTvCUgc0qvB6BSYbOZJJPyVEB1SXLMS+6VoG5ookDzZGMZTbi4rqMpOX/hhuACbrso3UVsJA0Ijugo7jGMBTyrMI4YkUz5LG6HEeuUEakoe5ZRYOSYbQLTE3mTBO1+3pi57fCt3xqKpr9w8+gXAXYpJ6kgqsRflcQD+eY+NKbsteWB0RTdUFOuxmWaBjEtihvGsUnn6lAHjVOOfNjdxbOo1IN4EBcEm/uNxV8x8pu8zaxrvqwWhfWf13cjK+AB3qo83IlU1NNdFj7X4o3w3m8G98n940/TQb5KIUleIbJ5NG3FwWQ/XjuTxlfXsvQhERbUDeaAVOKTOA593RGJP2H3+sJcCDzVRHQNJKmYBc/Wms1KhScGsk9pcJW+QVY5ebYFS0Ft25QCO2NNNsO7AQsWXjrYkOs6kqK0p8XPckSknuXdpIjFPC6q1yzJi0Qgv9EmlgMX+0M/rA2ZPKYCbMdhb9UVzf7yi4lPFyQjaw6kw8sfzQ49ep0a96ZBIq+MTMcpqLZOclk9DtqD1Mlamf1cFqoPJFZku3OyDcko1wjLRdvq+umIQH26BqF11l+srdHv+yqPs433tliklflV3gLeAt4C55kFPGFxnlWoL463gLeAt8DRLHC8l5uTtBwvDLzsAJT8iNJvlb9P8jSntDvg8TVKvBT+qZKbpuiXpWWBivwTBTfpJl70TW7BSSAo2csu2wCNeOnlxfhSJcA/AAu8DfjOdrwR8Bq6vkwAYZwfD4Wq9NPRDH684NgLj3s6ZBsv9ABf5gHBbwC9bWWZzEOE7QoU62ZtA+pRDmxjn8WsxuI85Mc09E3zGgWQp5PPo9nqrF0Fwv8cAAAgAElEQVQP4KvM2cxO2gVjziWgLA6MKdE8YvemaXpYv5ntDMBs+urOhl4O6qyt4rM5Y/Q789RyqvoEchcOvkqfN0jeZ04EBokoLQB8N5V9H7LSSQSVbfFsLueieVsQoNrGHeJAWNwc87qgXzL+GYGhWA2OKKDvttRX8XhwwYeVmE2eqrPqd4asEwSDQiRLoQauAQ+KKoJKzgyxP4KkZIq4+VUZ6lqu0wR0ESQEmSDPpFGds5AYLOSiDICm0vDycNitEr/dWFsGIzeiBlKFeBQSHsIBpFbfnWwIP7D7J/a974W/8MC77/3+KEkkF0ZMADwduH9JLUzfuZbFLhiX50VbRYNQIPjz6rhRW0uRCcnhlgqSrPtqVeavVH4qTFOMe674RsbjYcE2ZJVGpJilaOUC37NgVKehzIe072w9HJmSh8UFQvx/zCpcbiu/NZNs/9qWzt+kko7ifJliXpzWe8xbn/Op2d+5/Q3fDrP8U/KwuKA+1LxloCv1+tFy2fOGxyV2dEX/iQdGsi5tw0kclnWBVBNWQUqRT6sfArcTpeIxtajV2rJcaUK/8cKgLUIa8jzBPbaQdLLFSmYtw9ZDePDHUshLFfJnuSNNIKrk/eNIFO7rJCMGIheYu2g/c54llSvOfa16JAjs51ouN8qeeSrYhI7JmUtePrz3Zf/leZKD2sw+te6hv9N+u9WGDupCL0WNDnuoRYr8CoaTNIh0sr14RjRLVIm2Im8MdxHj+ZwpSns4I1dqGpUxNsvrwnks6TrEucCBDA9G2m6XHTTskU8mAjjZTZXFJLEWK7Zf5y3gLeAt4C1wHljAExbnQSX6IngLeAt4C3wHLAAg+v8ovUMJPfzFpHGeqWwBHLv3m/K67oXNL0vHAmUwbZstaB4NfEKgmSwKIJ6BzoA3Bh/wHXICiScLqA0wAVDAyzjyTwSUv1oJj4qTXUyS6kSPs3ydiEdGFe7gOMALABJmtULc2axWAoBCwgA6bFTi3JAV9yoBpmAbygtBwTEWQNNghDk5rRKYP61A0oka5ju1X4WsgPDBdpT/UrW7jWAmFWOECogs2Xvp4xcxdSB+sKsF6fZj03eqEs/h6xJ/ogy8TSmMNNuqvsh4dCMkmbwtXAnLmBYuloW2361PNjivKZ0jOxdiWZxoVYnImBPZEbDPOAupUwTfLvodYz99jnvBsJB1CwjNWKk+mksrPwWcJr5FIecURtovEtAvbwmWKjlxxBRwG6aVBYN55/bVChBYgn1zm4Ey4Hx5xgrNmndxLeQBkWv2veJszHvtmWedAc+A5iaD1VXlKt5B1HcCOkNDYdDpjSpGxzJ5XHC+4Gevfr/ZIxHoz1AtCiJEVgewfFI5wRaQXMj99NM0qylQ92bFuUDOKEpzYnVrjyNH98L9opwjX1IzR5hF6wz0zhWvXKFUYDG0SyS5LMUByUORFbK/rgtZNDNSuyiLw+EbqSeFvNie5f1v7O1/488enHkv9y+TKqIMTwnUfaJt42j7/cJNH+n91jff+C/N4XhTFuU3DKQRNQjjdljLLz0Yjl94e+vS+otm74FoxhJG8u1z5FZBKlHWgsBPRVLkeNm5vyeVCOZNzAuCGEHa4LG4Vt/xtuOc85atkEJHEBl2p2U7xEVN7TZSIqoDZBwSVCJ+9Iu8KJ7KHKniiAMlN1lB5MVxPS6wUUlezEkqlbJRzgMjbY1PHbrxLZsG4xt4ZlDus6m8Vt8bz+z9J/3aDnGgur9a1b1e2V2uz6Zivzf0+bjyNaUu0FOm5npHcQ77N9e1il5TIXO0SyavjbwvRkvyUJI7k0RUHqzS+YitsU6JiPXTuj73WZO7c9JWeI94T4un20v88d4C3gLeAmevBTxhcfbWjc+Zt4C3gLfA2WwBZmP/d6V/USq0ns/AovgVvObwUojMAy/FzHoGmPXLErBA6VVhr7p8GvlgAbT5xAPHZEIgJiAjbPYkL9O8+DMrlxgoSHYg/QB5wflM/od2hRfGmVqMfDne9QAxLLApxB3lQOLpLiU8jtgGWAKJAZhn4Bf2gJgwPWyTheLlH8DPZi5X87GkSIoFhje5GdoHbYfxDfsRiLfA+AzMZKryvFcLXizYHmDF4uscr079dm+BxSxgsXVMrm2tdnKznqvocUko0o8Z1+j/JkVkQKsLvnC+LUZelPEu6JKU203ELr9jCwBotmEDSAwS/dI80aYE/gtgzjdo3YqgIb7DnQkCQibNSr5xIcK6mDHnyAsQ2jK5uooUjDmUTBTxhF3eeG7hnsO9qQiuXCxs5zfjDKTypMgKfu8LEgnxoKGTKkZxnhE85ylEKN4J77rzjQg3udgS5fl4z+e3A7bFo0gFKT8o3mS35q5zX7T7pnmlFFJPROThBBVQeUGRjbCYVwcEdYa0KRzxYilvTahEI0FS18z50ZGReON/LgoZbeiku979ePdj/MQWNmPeySGKtMAeri5VpgWXPcWfebBFklCfTJL8wizNXtEajtekg2ykl7SuuL954cYr+09sX5U4R10rF3kyLyeeCUxSSR48ro42yEaPaC3226B14yXtEmnrGm2jfiEZino6uh2LAlXJDEpfUmdOZioWAZJp4oSkmLSFZ10MTJ3Oew4VfR+pKLY574MT9agG7C8Ddac7vuc9UeeCm5tpa+J5Rb7UYGYP3CUvC4xzl9oD97UXqXG8shYFF9HKpOO0Qr9fJoLhYlX/o8rAQ0oQUcTFcN6m2mZtyciMhXKaeFI4Uki7xjoPx7LwLFePayLdcAhKgknnzVPcfhVHa+6889JtxXF+8RbwFvAW8BY4TyzgCYvzpCJ9MbwFvAW8Bb4DFuDF6MtKBhCciSxwLeR6ABgAaJldNjdb7ExkwF/jO2oBk35yMhhKzKjlxd1koPgEyMdLAjABQISXXou/YLNv+Q0oBJAP+XVJeQ7OyXGcw2bJG5hjINDpNkAVrjjWuU3+aZt2gpRAuop15mEBmIGWNJ+sp+wQEZATlMGC1FvQVQOGsImBfQ6nIhNLKE7FYjbHBrStdUqJ0BEAostrcX1VBpDJNFcXjFbwW+SwF2uHBhACiva9HNTp7ipL6nz0SQtcDLjNODaqaeya0Dzf/lzw7SiS/FFwuSSjCAhP0F4AU/o3QON5SVhYSyhjPhC42khpG6d5NqAfmw6+7g0iDohEUMhDAb4qSHfSke3wfJDYzwDGgtgURUDvpn5CXkBc8FkMjCVKWpISDtVnHRtLjrdK9Tr5KG10DhzuP+4veMoUhEWeF/lUxZZeDRAtEAeScBL6n2X7tM9BKffrnsR5uDeF4/X3HwoH3z8X78JlrRF2sn7QEugbih0JI8SdaEOlR0QC/ixpnykVZaf0dhQ4O6RN0XYKoqcIfNwW2RAVAbfniVl3PziiXAvuE24mva5cUkZcS8JR8g1p1Te0Xv0Gq68kn92ytfMPu2aTXdx36+V9hvtx6Z7i2quLpYTHRWnUp0Ve/NJzP9z7ndveiCfwZ2TSK0WsrJYd4kGmGFVh476Pjj7n9jdOfWNyRXIYe5m3i13b4ljgtUJbYowfV1EVB8XZgHJc40iL4kmBiQ6Xay/67pPaZ3ru7ooRFpIX1d9mX86DNagRgnoXfh/kAxMTI4PvEE4sJucIoTHnoUPQcf3OTiRmHaSFJgNxLrxgfkcJcjQI0+R/jGz57D21zkECgNMuqRtufU3FrVgnQ2yQU9GQsr1SZRxTticIzK3f31b2eS5ZGUfyluBUaslGMpSlm9OYdL2n8NpBpAwfkpjoMBroGOya5rgkG7TUDGdK/kNxWQqZLBEu2DrxwbjLFuE/vAW8BbwFziMLeMLiPKpMXxRvAW8Bb4EzZQG9BFWXM0kY8EoHYQEYazOYl/JM8DNV5Wf0OnOz14ur2sxUvpvsB6APoA6/LS6FvcQDIJCqhAPbjFiDpLAglrzgQ3IggQB4U10ALNgOQm0z7o83V/JU7LSQLDAJoiqRwYs5iAJtnln8SL+QpwLYKkCWKkBJeQHEKBugJSAmAAIzR83LYnCUuBS+PxU2ZYyBGFXgWkmdBMHLa/XGpjQpcFGTykoTiWIUIBZtCBkQEvb2djyV3uCPMQvQfmhbtD0AbtqXZjNnfYHJillQuPZAoNXieExY+K0KprylbIu0XcaLHZKF6og4O+/bIh4XJWlh3geMn9iPsdNmyZtHHuMlIKeA2AiZHfatyYNhRHAs+7QkTqMYDIoDEUmgpogTwlKMyU6Yv/yc27Lg1mDuCXas4zXcPja2uDOUslUA0YKnnUyV7k8ueLfqV7/DkDFbgbcFr8cKcZxHFwR5sk4gbqP5wUNJ7/sm5jL3M9d9knpO33PXS7Ne3g5TDVsiJxiwiDVBDAs1n1zSOvlunZf4Etzzlmm94QHiMfKVSqMiG6Q7hipQUUBjsu3evJDQLgJfFHpFHDdAnCpoxhuHvu/Zo/Hma1k9yKf2Pzj9Z5/YP7hzdXltxSfIuYcZG6QY2e7+xH2O5LwFKJPIC/Zx+51SrIswPygptbtU1U/0Oul1LoZJGF6hfNw8GQ3/0/uWvWzy7Xv/3mI3GZlvzwx2j+U3zw6HHbkjGSR9J9ZES3fgm1wsi9hJRF3qZKL4C4JHHbnBcrSpCbZ+4acTPSrsXx7LJAXqCs8/iCZIFO7v3O/Nc9TiXDhPIqSisNsJEBeclyd7no+Y+KB8p//vqs/9hsVasWchpA8hFmKp0r1RomJX0hvqxN7Ig836PiImAvmmb+h7BxvICJHaIdxqQaGVPFjZi4hNYTErCnK1Yge8M3pEcilWY//1OkdTP5BWk7dQsE+/uef2RFy4PHqJqLLN+A9vAW8Bb4HzwAKesDgPKtEXwVvAW8BbYAlZADCB2V+85H5c6c4bN4yd92DMEqpfK2r11d4ICz4BWPCe4AXd9KYNZOAFFpCebQAbFpfCgA5AK4A8XvZZeBEnGeGx0My0K172C63zZ26xGaVcwWmTawGmqM4UZnYocSnYDhhOvgFOAEIoP+ew+AkWaJuXe7wq5uWM5vdntq3vN4vUaRm/gjYESHyFEvIYm5XWpf0Cd2IBLxb6pxACyR36CYiDxw6kEHJ5gKFnkshdpCR+1TluAcY7kyMzLyrGANrdzfLsWVMG3HZIoJPVj2qvyTOBsUV7xLNqqxIA5nntZWH1bN4W9rsM0m2eFqxmHGfcNEkaxlk89ExeZ0YdG1tPy8ijCsS9UiDsMhm4GFMdRwSET3LkAmOojaPgqUrGPx+V265scPBtKcvkKAH9zrkWnl1GuPB7NIgJaezOrcp21wa8nhFpQVyBpCy7K/rbrvtcNV/Z793xJvwlIEBYppUYq7gXVscoR4qrFa1Qc3IyiSJFmqHCZ4jkmI9HvkixMk2EPzhYuTwOkyQOB4N+2mxBV4zGq4ZXNm56DnlK80F/e/eLX9mT7EpmsvF1Y/XJg6HsKsLiAoHOeIFQF5AV28v6g2zn/kv9WXIRH0ReWPkI1H1C46yuw7kf04EHVEv9sBa14latPegmGxVZ5JI8zZ8UqO90oUqQ383aV+L+6eSqlHhWwALYn/zxyfaNagWrtHVjGfFCxJJkJnO1NTwimGQQ6dOiThj7Uxb0JD7IA22VNsHZCne/giQ3j1LKSZ7Iq8lCdlSmwXFkongu+mElvE2JdfWpPG4drHgtuHgRWo9s070QS6o3vCskdxZsklgZmmeKZh+sFNn1OgXjvgLSQm1pr9Y7z1bZXa3JdRjXZxbwN/zEpiU3caRVSpO5fepRsFa/J1KdW5/YhHESO7vyKp+zyvdTZNNOws5+V28BbwFvAW+Bs8QCz+QL+FlSRJ8NbwFvAW8Bb4HzyAK80CAFxQs3C27qfjkPLFDO3CyEEOZfWt0s4nIddQ9ZwYs1zy+8PNsLuYE7EBoQF7zU8wmow2ehzV0cBxjDyz3AlQWgtutULWnABMcs1Fw+VYsbKAOowDUhVaq62Rbk08pFHln3kBJST5SfdZQdgsLiWfA+bx4X5NdiV7AvyQB0J3chwOqEQJ5TLeQ5fhz1DiBEO7tY7fKaZmtoZTLoBalms9vM4pKwgLK4T+u+rn0BjXYoORkeLwd1jreC73z2DZSl/wKibyv7/T61yc0K9u4IC9qjGqFDABtqp4Nehxny9HG8gxj/aJdLgrBYWGULCQxtT0ViYAsb040UKoJzhyHAZzFmyoYujgWETy5wP4p0H8lJA21jP4J6c19hkTwQIjacV2QCGjZzElJsXgTlNy8NhG9YLO6FIyNElhTryACeHrqOCIc0qem8iuGVS/rLTdwgr4DTM6V3iZxswryfDaXB96PEUyw/f8M/OM8Lvr/rzjfpXhBCqnbdDHjdR5QBtnE/wevikPgJXTePsyxcputoJr/LUxgJbq7JyaOraBiDpEaO4ySvN2fS0fGDyaoN+t5ykcZDNLQa7TRcP96ujSOvKBePeuP2w/tGDyQrLq1FE4M0au8YrR08VMtmR8QDiXTRPUmeCDopTLDqIujJoD19ci8zabTCK2Ze4jErZaMI1n3MOAa/ePNH89+/63sn0yzbLYsfkNnX1wShD7oEss+vECXzbcrvaqvwIHb+DQL6bcIEzwDUN3VPe+F5hISnxReVd9VN8DJZjrpjnYKtOyID0uI+JcmPqS5zbaP12V1/zm+krKwS0Xe/FiD6JZSPpwzXAvY3AmPCeVu4Num2UA4jLCCiqNtJlcXGgSM8LiQHxXneogRZwUKdfYlyllJRgSYGEbDb2hHnvLvzkwEN67DayPPV3DfJrmvlaTEs/6DVarnYoaO2xL1xm/ajHpuQHOQTqSj5LrlY9SRKC6HBp4WHQkDNsRfQePwr9iOkfUOrGgrrwmbav3mB0D7cRBORFrny62NblBXqP7wFvAW8Bc5VC3jC4lytOZ9vbwFvAW+BpWkBXka+psSs51uV/lbJv5Sco22hJCnsFZ1XeAMF7DvEgs1HxHuCmafMfLe4C7yc850XcfblJRkgh8Ds5o2zSd95ATctc0gCgAfWIR1VndFX9TowGahTsW71PBxv0AP5xOsBQIH8AYwDLFAGQAVICcAk2jSfVW8KysrLuT272exTgAAjZGyWIUQG5+M3x/FppI7vL0ep0dK7gjZIvdCGJD8Rtntd8Bk3P3n+yGIyNUooW7USiS7qhlntS0KC5ygm9KtPkwWM8FKbZNwi3sJjZRsDVJ4sFaGKaflluxRZwdUhK2i7jJWMcXXa9VKQhToR00NiCNx3MkNKjPHY1sZW182VBDg7kB6DHtR3xmjIYpFADkTvC1SXaJILYMP+XUdQIFXj2IpCrqtYCrS1+FqZWr9QMsrtYLyzU+3XfcpxDuQllbcH8Sy41iad/mpd/359n9Y28m/EdT8K87RZm+kFHzw44Mrd71t2xHj/juv/YfD7d75uMstqs3kUTulCgO5gxl3tr7Ip/kUWNMS/NAUYIzm0XOuHKW8mSFnqR43D2Xh8qDeELM94mjfGOtnwqulkbEM3a6/Nw1qjEXb3jMfLxp8/8TzzGAzumtrae2B26EY5VPTrUfdgN2kMT8T1J5bVD+xr1nr1ek0hsdNsiGspL3iBOC9CPSPI+yI0wqKIO1IQBmYsdx8UccG99ZiSUTqXRmzJpoXRVu17YSa3AJ0Fyb8b1BK+9Lu3vfFJRd7IRPDM194r5kB6yAuu4UgepUI6zHneaOJDrok0PZFboeJXRKojvEHriu3Ql5deKI+FXHWUuXvEWEFs0R5cmr+p2JPQIvyW298oKNteCFaRjzUlUVFIZeaOuGAhPgt1QILoMCnMBC+SiscFJAKeWbZ8VV8etCtCViy2qPV/Xuvx5rpHWXuzmjQBuUcUEt6RClp/s66JbNMupQfUqnvqJoxJTBqBTG0qf3OlneNwyv5SDG7FlR13gaSZStylVRa/W7oN28QUizlCGd1zo0iLno9rsWjV+ZXeAt4C3gLnjAU8YXHOVJXPqLeAt4C3gLeALAAwC2Bt7vkLgWFvpHPLAkYWGPBj8kvzYMB8XTPjnbqHlADEg8DgpRcAgcQLMvFNmCW4XokXWYt1UYBQxTFVb4nFPCfcDL3SjBzzdJaF0AP5fKLMP2UxCILrAMJsVWKm55aynJSZbSDmgOG8lCPlgWQRoImVi5d0wBQLzL1wJqr1EwB232eOXaO0QQAeAMoL4np9aNA/coK6C7hd4CzUHwQU9cZO1IMnhJ5Oj/HHLrQA/ZW2BYFpgXVnjKSw4O92kIgMxrS1wmYZO2wMNDEab11ZoBKoG9va2GnSPzxjcN9AOd/iK9DZbWzFm8IIYIOYzWNDx2lwILwwsS9Y3HTxMlX4ikpFlPPLcZUp1zrFKSBaF3Z4VkTFYZ1nVt+H5EazMkgGV4rAuFJ7cy/hfgAJDwkOmO8krwhwrFEqrb//QC8La4P0zeNz4/7br/8Y3we/d+cbzUtRP0NyzbAmNzIn0WSxELj/KEdxOt2fiPZ1143u6F544WzSvqIdzVwWE6A7i2r9sD2heAZNcp1Go2suG95YW9/k9oyGUBp87tAjcS9XrJWokQ3C9mhv0F49nY5eOJku27Ys3v/kRL5vbzvqdHTthiJ1U54h+WmY1CFeCiy7yBtVSIaVyJvFmbB7NpJRbueFsS6Qj/rtb73h8/VmeGlzqPYCxWCAWiKTr1AWH0uTbOaXbv7onZW6OeJr6XmRlQGtrT3QRsjLpPKIJ9RrlaPXK2eXl2JFy0RPvEmt50ptv1t7PqS7hrx0XL7b+n+kDL8+L9hodNfx/CALm7A3/Zzaq5UEAAQENqQdK7C7e54ZhTzQJx5XPDtUfTsYM66vFPYD5X5HM4VbLzIgyN4W7FN0lS+7shTP569WeYebiuEh+45FcfBiNZ714oaG5W3xKbUr7HufvmuMCjaqCBv12xFbylBHv+lLjaM8pLg+pXNUKRvKCTlL27fnQDdmerLimNXnN3oLeAt4C5wTFvCExTlRTT6T3gLeAt4C3gJyTecl5Sql/4N3JaXbi3ccv5xrFqh4VlS9Kgz0YZ3FleDF2/SiIRt4MQegYWajeVsA9PNCzgszMxuZvQcZQBsxQMZiQhzvuYcX3YUiDadiXs7ByzNtFjCgKisF0AFwQJ4AxXlZt6DavHQDTJoGNWVjXzwvkBviWMqPHcxzgn3sZd3kMixoqIKYevmnk6hA6spkxGiHA4EqzFg36Rd3KiZWK3YFoNmjSoCGFmTbPFpO4pJ+V2+BY1rAgcvlmAAYTbt8dDDo3UBbLTwtGArmuFEjOFjJOMmMZsYXxhS/VCxQEhcusLO8LhhHLVYB/R3pJCdRo2SMZbG9iCExJRLB1it4t5T7g7BbkBkK3J1zP5o7XrXGocwPLx9ZiqnjBN2ex2bnWaiC6KjFgrVj1X0qMDwFZB5WCOO6Ilpz3wDodTI72ln3BK7vFuIEoF1XeuCFeSyRnfiDUnoSldJ/88Tc9X7++g872aM/uPNVcuEQ11DIUyVitWf0ZW8mFaqZbDSU5FNT5EJtR3fjyLbOJZd38+FL61Hv4uWNAxc0xSpEgSIWYBcOFzq9PB7KXzRx2Rw988Dsrnwq7St/Lv6HChy3ktpwayatt5J0aHgmWLZS539sXWP7YyON6Vk1adiemtwhWgTlllnwYnDPBDw7KKbGTq3D04V6ctfWb1dei2kh0iJSsokQ7r7OtsN7+lvWbI6/3u+mDys3G+N6xHPCqiTPXt0Yjg/omO2dw9mhX33Rh4/6bGnEBecs410AoXd0lz8gy5uc4CXqtWu0LlYu1yqXo04OKlSMjkzeGLlrUyKkVH9dJxU1pvU8w8T6pCySxirjWFXR++oUiPn19dLnwLx5aH/cx4prFAC/2qZ7tmjrF8TKjPKeTg2/VIE9Oj+ehW3iNbFsU7qLspW/j/kRvcdRSTtn3xp8WU26px97JAd1gy54saJtr1ZpVqXdYDlxSrQfwbg/p/rdLjbNyTdpP2wyAdElEqPwjgiDEY1qQ2pOYSkXtdDTgjxZ6QvvEe2vc6vDuHYyxfnkYeH6tpeGOpGa9Pt4C3gLeAucnRY43ov72ZlrnytvAW8BbwFvgSVnAYJri7QArGUGPeDL9spLy5KzxzleYAPyLe4CxATgmgOJy0/bBihBMjCJF1Q8KCAl+M6Lq8lBsQ6Ajt8AGQbcV4kIzluNWVGFA2w6rHl+nIyZ5+bH6iCAJIgGrkNeqvJP5PkRpa1KFtSb/QEV+QRoIFFeZDEIuE3cFl7mWWzmK/YCZAPI4tM8LNjHynGUiYonU6ylsa9kcygoYAcz01eW9t+fDPrrFhAWEnNHTn6wV+vR+YawQAZqaRjKl/KMWqCUcnLAMhdWO4Wc/LYIsyvU/m5V0mz6eRRTcS3Yb78DdAtyE9m7wzpu2stCHb3qRF4YUT0oyQuLM8R6xmHGWcbgZUJPGcNnRD7MRyNwKk5aHEEcYnfFFciU8iKmhQt6c8R9x+2tpDHaBbRgrOYkgmnL+iQUhJOByiFHCAiukV44b5oIoJbsV57j3QU2W9wLkDwKQ+6lIqrdvWSqCGbtbgP4E6SNDxxiW9b7Pldet/z76z+Zv+uO1wdxJF8Iha5QFIrpr0y+TKeLhnp5q97NhtfMZkPD+/prL9zXX/PKKMqXDdemgpr0p4aibtBUaqWH8Ppp1Gq1fG0cTw3VGpAqbrl78oG9WTrVqAfZQDmLRIS00jBupVGzNRMObxA7sqGfNCYaUb+noN3bmmmnJIIwBXJcsqF7BnBlmxCvMqH1BxU/CG8QgofIA6UAp4tyYlFJdukY7cexGCARGcHzgIb07G6t+aC+/1C9GW0a9OQ/0oxu1HkPD5L09rgZfAvbWf6P9Snywu61brf84/KiIFZFP7hMW75LNbrctZoGslpu3SXK8zYl7hsHlNu+IzMCbWOyhcB67QOYzzNPMWHDKAfLiN3VF5IXxlsiTVaQHYXXReF5gVcHclTFhI9c5dPx/fpFbTXLH7FTq7l8sT544omrtlxrsTxOxCMtgkMAACAASURBVAzB0HuDLb88Gmz5z98bfCauBa9RjIo3iz14rUrXkHcFVNat6gYQT2uU/c+pDW7VOp6ReI6nf4l0cpJR9VoUTIixulAH1d1oVlZgtbha5Z7RdC68eiiPpL1Uvtz5qxxQj2qWnhiHRVx0vbfFCVWj38lbwFvAW+Css4AnLM66KvEZ8hbwFvAW8BY4hgV44SQBABfC8n45JyxQelWQVyMDqnEqAOh5keZVnEDYvGybnBMvoGwzjWKLL8A+ti/Hu5l+5SezTzl/9TnHJCOqZEXVdtXtBXB0cgvHA3Iwi9Fialh8CqAEZk/adGhe1G9T+kclJA0Ad9jmAlIqsT/7VIkKygIIacCaAWgWhJv1c0SFl346ucqDcBCoS5uirV2m9vp8fV4sb4o2OCCLye/ok7ZB3eDltdeTFSdna7/307IAYwAk5r1KN2mUGjYFoeKsbqY9gbdvKLX/GR+QmPPLCVqgjHPBc0ZJKLgx17xcmJ0OQSAg2YHhdq/iO/thb7Y7STntg86+ZJMyPCGGRV4IXD2CRy7uh7buiLuO845zBJSOE0MAhu2GeF0rBOTmnlJ6F+aKXZBD1gN2E42d+4M8v+Y4eP0OY4G4LlRA4wMHBv2kPQh+SHi1lrdf/1E5VhTUydgHdurc6bXNOLmxEfWuqYe9zUneWNkP2isHtaGJRm0QZeJDZtNhuWyEh8Kov2ek1j80UpvJ1w2Nxd+76rvw/vn/2XvvaL+u677ztl95vaMRBECwk2YRqyolS7Jkx5IlW5bLzNijRJkVT+I1lp3JrGQcr1njP5J4Zcay4jVpE1vxKF5WLIuyLFmRZZuiOimRFCmSYidAgADRH17/lVvm+zn37vd+eEQnQDyQ5wLn3fu79dx9zj1lf/feX7fsaT/7XD167OEtzfmuOC6Gunl9UOsJeW5sLfJYhOJQdMdBO22MHw7XbR+Opw82IgMs3C2Qb1T1xlEUhYO1enS53EW6nSUnG4AZ2mIkNwCXhWSdqf5TXnheWFhHvhsnG30veMR9WRdszbq5U6KLRCPqdrJrdd2HBQFy/DF7hzNZhz8RLBZf0bVF8GldhyL9HUrwSlAUKNTfqi1CW+2o8i4+FMrLGTBQZox3KFf6oUj/VGd01OClXpOK42WM4yVIYeOcskbhoSIgQPcBOBkBFBGmkSbpob6wSMdEWUIGj/S1fvDxLft+BbnW8MDQ+hiC7pPJ4nc0+vmdPwoOL/y94B5loyagYqvW19bjQJ40QVNABjwZk92M/jX4G9W3h/WbUGZm2AHANq9XxVtiKCrkrKNjNjA7zrPdO1Y+SoAiQ/LqQObr2tmyQQvGIZBwdyvS8DMpTn+ul4CXgJeAl8AFloAHLC5wAfjHewl4CXgJeAmcngSqkFCm0P6GrvKx4k9PdBf8rErBWyoeysWm34xDUNIzOTceB1PIU76EPsLinUk8v/Gs2K6EJ4WFgrLrLfSShe8xL47e5x0PhDClkIWNMkDlTAAL7gGAhqKDfDH7553Mc8LAGANdUExgWfi0EgAF74OSgvfjXQE+uBfKMe5RqiHKhfk7+4wAlOcds3iwYrVETv1bYIV5wSDPcQEVN6neTlbWqe4GeFZgxSzrdkKSoAhB2ZLrWqcE9Bbsp5azP+PsJdBDCr+o+keIuCfkUHGt6upAySdMhCGpdEUUr3S5Kiqg5z1KDojT9Yuqo77fPI0iEGjBWYYsmIdLW94XABIl11IZjwvZWvx+fptnn/OUkKV4QzGaYoUc6ld4Gzy3pDiWDblDB9Rt5ICfOFj0dDe26ZBSBdgJw8NKBxSHbl6FzLPo8wiJOKFLOwIzVPj5iOzY+3UehOBUhtKu3/Uvbv+BiiWjAlnChUatvVh8drYrj4c8/ExcJP91Meq7OxzXfW7QNe9Ks/yWpSDfnsSFQvpkw0XSp/BGaiY7hwUI5DMKBnVIYXx2JsnSrrHGobmx+mxyRXPs0jhMbkV43XzuyLML//mL48m+ufEky2e7I8OdoL9f4Z/GQjlzLGTDWzpZNCaecKEI0YDIuzcu5MOjQ8HMfBykTk9dRsmSjCrvAZFiR3Et6ncNrvZlmS4mFFAmwEbGAngW4XXUU8SUh3kl8u4tfSFtfStPKX1V95iKkkh8Cji6BJNxEr1bHiR//S+/+f4n/tlbv3B238qS+u5a8HXCIel5w1q/0ZUEIaFyeVLkwduU6MMfVXpGoyKMHJxHjMu3I3V3fhUAX+WiSFhuj/mH9gIY5TXHLsbzQA3m3BLCkLePUurCMKV5PBC069s25dHAFVwc5UuPTk3/P3ua7ScMiAP0aQm46B1/4HlxUs/NgT8MXmp9NPimToKjQizuwY1yr+HJg/o6rlLhjOlbqKlUKbP7K08LF4ZNxX1YdYrQTpfgPVEPgyFDDVdEcezrWmb0ral2uO+x6YjjS5DxoK6n/GOBFo6Y3QMXq+qK/+kl4CXgJbCGJeABizVcOD5rXgJeAl4CXgIvkwCKXsIgfEQJK9OveRmtTQn0eFS4ubCSkZmaQod5JhNyFPYctzjrZdzlMqGU2aqEBwVKGsCKbUrcA4XGOiUDM5icAm44AsdqsbkuawvfsVpg5MOsaXuP9U7KTwVekB8URBBabqgSz4PjgHAH5AnrTsK5mGcE9yRcCwpyFBW8N3IApEAZiTzMa4J3JY/kifNJTgYenFhdnGf+W4pcyop6RP2hHJIoji8RNCGFGPrCsvhl3iudYQYvCIomypZyxdL5sBTBKJz84iVwPiXgYrVXdZX69oDq4oTq6mUiDK7qKbpqNbaNgaFOa5H6TDvCNbRLeyvQ4qQKx/P5Aq+BeyM7a49ds6BEe2z9GyA7oALnHXa02eLAqWH5rSKSolbrjPIolepODe3U76VoTDVsHBdlOz+r0FD0CS+qkLfqjuJDKLZoe6/OFyF1JuBU94iiMnwiJudZJs+BEB4NQJKy/4Rzo1Tm11Vv1BcV0woBtBSFWTsOO7Eu26BzbhRPhkIZJSKiTrdmYW0gj3EOaeVhR/QWCuikCD/79YSnakHnwcFk7rnN/bsO3Dj0PZEOrJu8su86Qhu5ZefS5+6Own2H5OxAExqN1qaPKpLT0dG8cUhhpBZfam8psiwZkAikvC5kkZ8MLqYDY0vJwOGheKYnJJPa36oHlkdEsKjE+IL2OKlHInfOp5Qp2uG92g9gwbYjotYCqAzAzBq5O2Jy/V7UNfdFieQZBD+adrNIWF8ticMr9S1dr1BR35a3xoHVxN32bidbhx9w/fYehYf6gkwXYv27RsVDfgAN8LbAy4LQpt/Vnq/oN2tK3rxB5vU70R7CQymMluOzKHktYu3njgZE2JdsIybL2GoGCnNTKM04BF9ESbtxxfCB8V//Rbuk2Xnyvv6lB8iDheGkjWHcwWLgHLwdmUAL1m6pOD2OEQkhn7TjU5IxZNvjokPZpDeI1Z1CsjIlsOJHlUVkQjlDxM243nkoqR6qllHXg6GOPMiUZRdwzV71ZQOzqm50CMam5CxjJD9t0qfjwcrYjHdhDMa3au90TJ79Dy8BLwEvAS+BtScBD1isvTLxOfIS8BLwEvASOL4EmJYwASmt1sqJiF/WrgRK00jMOstwFxaiqYpH7eaVFv6ASasp87kOYILwARBBXqqEwgVwg1BPeCGYF4YBETY9x0r+eODCyQAHA1M4pzdclD3DiDtPJmnj17B5tXlAEIoFTwl+oyxB6cQ0H+8KwnfwbgAahLbCGprzyhAg5drsKRGgeWe4MA1KyHa1WuJkefTHjiOBymod4AFwjPpGuRASyhkqH7OUmhLqCXWRNohkcVq8fL0EzrcErELSltD/VYSzL8cf5F1BXqifdyoBXOxRQmGHss7Ios93fl9z91/leRHI44IycdwIlVzZplwoo4Z063KxCFrwLKSlytUAckAN+rVxkWvHQeZ0qCo0DouhO4a6IRPtQw5KiheGgKdQvANRFtTUhXY6Cu1TAA5UlvryxHDtFac61EM27YlCLsm7AoCkyKkLixXPBX0w/Q6ef7LuD5d01VZd+j4973r9vjyoN6TIbzZF8C0fj674OkR1LdLmqNN9XJ4VO7th/elmvPTIluazh7f3PZkpdtHQRO2W/qFky2XuRYql3Xr203pvvAdG4yQcFDgQpNIqi2W6NVV/aW876B/KOvXhhaz/UhnV15T9uJsnDQEXtQrOOWH9sXFFioBX2mQMGFw4IyVCPQED1JWk/5biuxyKzGtNCKk9ikZ1OM+LF7S9MyrCS4XLSOguOtcbVQJPaf/nBVpQrhB2nzAvJzyQOZ6KL6i37pea/F3K2S36PaJ3A7S4RE97h2oN5Ny36pwv6tE7lCzkqXn1MDYiKJTzdtB1Q7rPlNbUsRU9jgFdJ8pM7whI50KnMtf3jg1pPAmg5ZZ1R//NfKP9/Jv0LITa0po2w4wpHNCFLJQ6xT3KD+edwAdFXgyEYWKc8ymlXWqOfkKF8AY9elO3zKv4XdwY78P6Oaky+bbS05I9zyWMGvUGEIP3nJD3RJjiZeIKqML1et6p9/XZBs/SmeSXbwwjEcrR5V/5wsvi7LxnTljY/oCXgJeAl4CXwPmQgAcszodU/T29BLwEvAS8BM6HBJiHoARg0sey/3w8xN/znEnA2fJh4ugmmeVEl0kioIKFtWCbiSTKehLnAkih9LipShYuiXNRJq+ESSizeiZT9eO9nIEeq6b0y6BIL4hxvOeRf/OKYJLNfZggAzqgDAGIMe4Kfj9TZQKFIwojLKCx+mNtii8Ui05zVd3PgT9VwsLfAxXHK8mz28dYmHqFtwtWr9eydgpfF2KnrBauGrNN3PrChR+hPLDcpKxOEmb77DLlr/ISOI4EqHO0FdQ71k6JqJBQalilr+6pr3kZUYf25Y1KKKtpSwBGaZs8YHGOqlcFYFh7nAnAMEWz45ZoypZ9OAnzRhx0diy4vhDZ09bTjxFyrhVkgA/LGcKdoS8oC5DQUQrjo2LOM67ZJ1tz9Y2RLO/FYxFGAlkLylP9jwi4c4VHsgWvDbwp5H6je1mbJSWzi/iPVp46URIwByKoDsPbRX/ykzJ/31Ra9otQHAVxns0oPaXfe3TN83m382g3jF6Mk76XNjVeeOnOkXvk7hA2+qKNi1ON22+IwyZtqSzcmxONcPR5ZYl+cCpLiwklFPXu+Y2w1R2MZvbNBKP7FovmhjCOaiL5rreCgSmFito/khyW94drdI+NltUTOov6LrYK98a4sfA+1XijzIK03oJZ+iXFCR0cJjSllq4u6we8UErlRAfPxyNRHApUiSbaiw4zuknn3aX1N/R4DA4SARc8yBkKnC54Eb7P9efPFn8VfMZ9dyKV1voG5WejRrL4Skyq9CdVIxjjADzdo2f+UOfhDVICFOX4AY4LtsG8CAPGd49vzqBU8MnySGX1qOBEZho6r9W8bmh6+BdvR1DisEjHFj79twOL3wbkuUL543mL+gvhN/XLwlIig0U9L1fuVLfcXzwtbGxS9HpbAFro/MfaHw2mRZ69oJPmJPu3KCDapcLcQsl+nUAMvE1Gsjy4VL+/p+1nCAulRH0HMKFOrxfIAe+GAwFVrLHuIWzNsLnKJbfC6lyNKKsN/TSAh4VsszLMKtBi5avjGr94CXgJeAl4Caw5CXjAYs0Vic+Ql4CXgJeAl8BJJICSdzUPghfYGpBAxVPRWzbGKcE+Jq5MPJmwW0gTFBso3gAqsPbkONZwVythOYqXhWJpO2Ubx5h0lhP1crFJsinzVwMLpysVrl8NVtgzDDCw373AAe/E+6BcIDwZ1oTs4zfn403B+3EPgAwANiwuLdwC+WM/1zExt5BP9qxeLxL3blKieKvA0y3V0z8PIAzLXKzQIcql/m0iHFQl8+W1PC5wu6CcKGPKkrBQhIPy5XL68vZnnqUE4EiRRxBtCm0GSk7q64JIhksdnaFr2q48LGhr8RqifaU9ApQ7pHvMeL6VsyyEU19GW2ChdBY3NqPkysEonu4W6cF2mM+nCstUtvW06bQjUkiHA5U1OMpV+kBFakrhqwCwgJhavBeJvBzS3epZrgm63XHHn5EkffKA2Kxt9aHhoq6iL9VS6WVTHqVtR+oskBtvC1FASMvPSRP6TZs3rsoyJY3/m+TpcXVQE0VyeykLFudLID0MdygfeAV+o4hieR0kqPSPHvngVOeL2vm+R34sahV9S5f3/w+1oWT7ryrmEfVSl6T3Hk2f+K4iGQEMCFAJBRiIW8DxFoSANeuiImsIUdiv7LSLKOzLw6RPHBZbZrOFg1NFfU89bHcc1UfV5YfQffT01FR3Iwp3r01wLWIkuq9BL60waYSNkqRGYPUAfoFWRAeRc0PnHdLtRD4dPCZujBs0hhlXaCiJNd6su9yq31cDFOi2FqbSjWN6wQuedEoAIw7gO/qSnk95izw9eJNU/pc4KKB0itmg9NPaGtZvdDMPubIsAQ7GC3zzlAf1RF43btzAmYSYKj2Ne8GK1aOZVcBFETWjhb43TmbRKGOroNF5+vnJw598IukcyVzIKjxAIgFZ/CrHXoDyZUhL6hI55jheH6VHBPJxnp+AF6s5Ltp58JJu9CV5SUCqnam1+qBkL54dQWRlfX+7Lr5Dv9+p9F39/qYSazxhAIx26hUu1XVbtT0mR50+3Y+QTyX65QRQghfut3a4jMttR6uafluYK5OUGYb4fruSnV95CXgJeAmsVQl4wGKtlozPl5eAl4CXgJfAMRJ4w6XDhYi3sRC15UThf7zkLowEmDdaCCNyYJ4LWHHahJd9xlvBRJxwA3gnsB/Ldiz+8KAhPA+TaRQwTDZ7gSp7u17g4kS2hGcjCZsD93o32PuwZj/KAzwlCBsB2EDMbJSH5JV9KBSZDBPyin3UW8IbYC1peUUJwWScd0QxcTKvCe9RcTYleYprqnBQAGHblKinlIUUXs6D4pil3ugLOu0lFCh/q/Q1pcerMqVu+8VL4FWRgIAGSN5pM4n7Tn2dE6/Kj8rL4i2QwmfpMeHZaavoJy2GOwo/6jBcFpkHLc59kVUeF3ha0Gant8hu/7rhOPnhbFY8P5/jDmEh/egHjIuoJPEuQVPWHDsozSsqbfEVFCq3fEKAAt4OgKQDQdIQ+KRHhJH6yQJgH6Xx0+665cV1NSLhcSAJSfwWWKoXAB5KUeXll+PhIbJtgRkKAaVnUF92uPsVxcO65nsy59+p7TmtFzt5Y9mj7Fdu+utc4zLlOb9NXSNeke6ZedD5t4vZ3kO4SCgX9Jf0fbwb70+9nGxES7vzIl46mk1eLcX1YFNs3WnYHF3K58byuK8RJarMUm+7SFcoo0skosfrbeVN3ValsD6GP8ts6h2c4bwCyAGAxVbdblSZm9OBPVknP5KLGZ28oUXXsct03oeFUWdCQZAriym6XdlW6ZRK74rv4QWdD3D4iIrt7SqNd+v+tyvP65yvRSgwMQ/eo+MYcjBmQGHPd05fZMYLAGGzFbjV0d4l5WJa9xjU9pDu0lgOUFhhVcvmHT0jpCwaTGaG3ndNN1kPUB8020/uqXeeWxDuANk38sG7hoU+cbu2uRvABM8/Wvl9AjTs1XN3aW0hLJEJ8JaFxuzq3bPhTwb5vv8+ODTScP0mcnhIHhWqL8GNkvMVAiAaNYEQwqOuUSCz9brn9fLIGBTfxT2qkYylGCcSgop8TEoYo7puSFnsDYsFauvGn3VhVKqAvAHfF3WOMad5WSAJFxbPe1m4MvaLl4CXgJfAmpaAByzWdPH4zHkJeAl4CXgJrJIAluy2MLk/l4pqL+yzkEClHDAvBSaMRm5tyjIm4DZJZELLJJMJOEoMzoUMFsXJm5XeqXSVElaQTI5LYtIVrxrzqujN6WoPibN4i2MusTrVe1+b/JZhGcq8A0w8oIQC8EeUnGWpFizvH1NikoyCECtn9qFcNOU29zDvEu7Fs0y1svodzXr6lb6Xv75HAhVYYV5AKHUnVJepi8My0nXj4x7FVyry7SP6/QMdw/rz+0ooaig7H17H16xXWwIoPmlDUGjLGShTiJtwkxpcFJC0rxbAjDa4qXq7XscBgbHwRgFqnmqnVLa+2i/2WnmegAvXjv+X0iMr/8OdnVDeFflf7S9jdVUL5WBlYH0nympCN6EEPqKS1PG8LygieSPgYuB4DsRLkQ7rt8IdxYAFeEngGYYHmNS1hfqWiOfq2hDAgsdx3ymdh0fGRgXVkYdFjNKZvlf3lR+CXHWcZ0eeQ3gsQCz8vu73tA4t6gSB7zhL5Gk9akmzraOfboX/YIuIlIvOrXEY/b897/V/yf3je938QFvuHLgCKB8RyuNIOcl5mLaX+uPFg9PZVHwkXb+rnrU2p7XacJjEtUYxFy6l9bSpkE1Cjwn2JIpo/dHrQ6RRUgsJOlFsILc4MOPlNQeEgmPO/4iHkntyIsINbYvsu6hrA6+FjkJLHZakjyS1eMpF05Ilv7wu3qn7Tuv7iXU+BgcWvpE7IgIzNDjO04/NjxT3nI+X5X6FiMKAAcU/AIFCccnboubGQpdohEBfZEYcP9C2gCsp7AkAVT5PPCbu3vK40T0AX0RO7YCPDNCpFLh+U954QqyMLlwuo7Bdu3Jgrv8dd1gO69ne2biYVz2pnFmcLwrE3E7JP1QBJBB9l84uke5NfjMZbWQ6Jwye117aIuOK4B14n67AC+PzotQOSQ6HBBTsFaDwnF4Dr6+3yQPj2mai5+C1EQcbBVasl9wX3HOC4FtKnDer4uM5h1SeY8oH4dRIGIr0KVuOTBt0TGAI3jPImzGXhcFzYFRPsvHdKcvO5OTXXgJeAl4CXgKvvgQ8YPHqy9w/0UvAS8BLwEvg7CWAlR6KXpQyV1STj7O/m7/yXEjAJoFMAE0BbBajWOgBWKAIZvJrXBUGVlymfZcqMekk1jpWdyhQUOxzDttMWnsXm2DyvLMNA3Wy9z4eCMZkGGUD1n7kjTwBQhCaAcWQhVxB+cR+koXCArhgos3CvW1ib3Gh2Ye8HLkn/BRVrO2T5dEfewUSqMAKq6PUWdqUSyT7d5XrqI5Zb0+EnUVZrj+g31i9okg0JUwLi/dXkBV/qZfAGUtAda6rOkybhFJuQfWSkDN/LeDiLq0BfC3SP23QiI7TtgKc/kXVzrg2VfcofP09Y/GfzQXF39tWJ2V9n2MI4/oBkvFdsI+yon+kPaLvo59YUkkCOuA10ZSmnmPiktDfIpNnRXilrhoIUgW/EWClvbRpKmcHdvAg+iq1VS6UIFwVqhuxIAZ5V0R4ZoR1ARSO49uFjHJW9OF+pZ3aFmgRHqhqEv00+aAPnBdOQP6yRr1VF4bQr8BLP6c7OGv9avlPUdg4+L/c9MXiE498ALoIZZAsitPK5cMBwt0H594y//35Nx1Ni+Rwf7i42Albw1G3q6hU47NLaf/0cDTdEjtLXfUXYCHWvxD4hsh8LK6SV14V9uCy4h/bhS//0rlsw3vBeWL3qAn0cCGVBNXsiaNwIq5FkFATWKoRx+G1WRb+pHIPyEdYLN4fa38W88JzvgwKE8W+5fGIwkSdsF8I3xu8KEX+l3U+5UNYpXcJIBhT5gAJ8NZ8ixLyvE7pezr+uNI+B1oQJqok4OZVFOKr8kSNqj6p64i5ATEwoAAAcCTV5mnRrW1sHJj41TcsyyvIsqH5r+wWjwW78PQo13htlONs7sUYjd/0eyMun4nqF2TiDhVy741sAHXoS3kHrqXeIS8S7VVKyKjuV4J90RHnbYGxB3UVQu3bYzgp9AQBDtzvXSojDD7wuL1H6QE9iHHUQSFeA9qmnDZRjDxLazxAGI+19FDy3NY+wIodVb5p81y9q/KllV+8BLwEvAS8BNa6BDxgsdZLyOfPS8BLwEvAS6BXAkyCmCgyycEKDWWwt3C+QHWkskBnwkgyxbv9thDDKMoI78QkFtCC/VjgEQKKUBbwVTC5BtQghBLXO3LFqqx5u8pG0k2AmVlb2Izz/eY8F8UR1vSEYMGrAiUDAAv1jvehLqIwRNmExSr7eQfWTLDJL8ojewd+98YxNxtICxXitCXn+8X8/Z1ShDpJvcNbS3HLo02EgypjkCwvKDhEFlpMq1wox2Vlolf2+lp0ASVAvaRtoj6iJMQDaEZ1lPapr4d/GyP84TxLUf5R1/G0oM1CmXdM/KgL+C6v5Ueb55x7RzwvFC7K3tdAC37TZ6DYpfExTieupa9TORcvqQfhOMQNAs6lYS4KWZpHhIeCXVrkyxlKXHlj5JSt+pgQAu8FnQdoAYe1PCsKhZaKG3I7KL0X6xpOuQBHXcCRXXrGs+7+USJC5XiD47fIuiLLdo0iIaXg3Aj1Dqp3RXzTUHSZwvl8zF5Iiuf/MJuG+961nYg9QfBrN32++MwTN2btopnPpqN5p2gIuwAh4alFIh6LOM8bw4vRUDOVw0hfOKcOs16fT4fr48n+vXHURUkeZlnRF2bFkLCKwTgJZUGPr0dFMo5E5Evg9PKAEhVCUVJ2V0sFbvRWtOVmXsd0zUFZCuwIuvmlKPtF4q1+wIEj6hsKATYhBjKMN1Gyz8sZpaljAB6Lv//YzyoqW0Y5MR5ggefC+nPklh2H54Jv8CEHLjA2yEU+XejbVHgkbZsRB56bP65ESKrHdPwlHXtCNYJxiHFe8WbcgzbggM6hTQBwwBNjiwMV4J0oHC9FuDBw61invp3+zo1HNu3/538yuPhN5cX8UNzYi3aCusS4jDUgBdeXdNt4P3Qgi3fvi7fDFvfu5L1sVwCByJN5pJpxBjLKa+9xNW6+++XgiWJObVEavKSnv1f3easytUHJnaeEHLjX9Ur3Kn1J6WEdVxgvl3/qEWNGyoX3duCIyk11OcArCKCPb8mFgOJ9lSgXC8Xmx1kShl+8BLwEvATWsgQ8YLGWS8fnzUvAS8BLwEtgtQQAKVAOM+HCpZ3JDBMSv5xnCVTgxGpeB/ttnhUGVmDNxjEmtKxRoplLPhNgFP5vVQK0wDIUXLz/zAAAIABJREFU6z0Wi9Vs9zELVANDOMesU481ozyz9++dqB7vPkYSTr7hqICv4FEl4ofbAgjDRJk8Gj8FykDujSIcAAMFNxNpI6W0vJsSi/e15+NdcWZv4c8+WwlQJ6lz1D0po1x7MiqC1gZRUUgloWuEno7ye0G/UVRRpiiITRFzts/313kJvCIJQPReeVnQRqGoO6Q6CrBK23pZ2ZaUzZyoCSIBFrRJeLuhBHShpJRou6jPfnkVJVDxXPBEwAvKwBr+0uJ+JRQi/Sh9jMo3xIKcdovjUgxLs18ovFMu4uo4koJZt4jiuhqtuhow9btOWy+vDPFXhJGs7qXczzOF95F3g9t2Uf7V0NXa8rJYkKE9nhXP69huARVHlERZXB9yMZQyh2tVMZiKK3UOfd9MEoXpQiaOg55lx1Jxzz98Mk8an53pkxI6TYs4/6XHW8X1gw8VPzb65+mlzZ0iAE+FPcTRSHJYGuc0zfJ4MA1qzSyTRl2aifl8OJhOJ9P1xZ6DfWELdEfOQwVhj0RAHgzIQQIlNYACskNmDVX3UUkApboLGUX1d0KtPoNeIKN0CnBeFdUfhwJ1JLH9ysxzurYhUGS84rIf1jEU8turMRC6kwUBFYm6B5WBolelKd+f8lOMlf2GI+lmDIHgUI6/jKNKoZHwNtijBxPyqOWAAECLWP1RTeOH2I0h1rsSn5fCPgxuUmkCWj2m0QQhCV9QOqLjlReNAyEBKSyUJmvAD+7DMkKBtmvXjC7Vr79aHhVps/P4juHWXy2FYaqQYi6/gBVTusdmPZ92ZELPG102R3FCU24AQ7rVezkSdQjc3bPMOGXY1b2SpBuPEOTBb+P9cA1T7cdd+b3Y+Xzw5WIpOEp90YEbhEXhXdKvVx8SH4UDUBQ2CuCFceGgzDkeVdEdict3570pE6sLELVTwC5ElJKNuRwsV53nwKTGfzK/k0pCfuUl4CXgJeAlsOYk4AGLNVckPkNeAl4CXgJeAieRAJOQzUpMmG+sJiNeYK+OBJj4MWFkgkqy8AdmuQY4wUTUxU1XQiFMYnJIuADWWN0RjoCQBzcrMSk2N32z9uVall5LOAMwWJ+PMFC9EmRSayE1UERArk1CccL78U54UrDNuzMRNgs+9qFkYpLN+RZ2iIm1eVgYWGIaReeJ4sGK3iI479uUC8DZNiXz8KnlFburlQUkxkWWUxdQEAGUUo8BSI3S9Lxn1D/AS+AkEqDtAHCgjtIm0wbTxm4jvr+FzunxGEJ5CWBhilSssj1gcX6rGO289VknChNk4JH1JWYJTn+H1TplyrYpfJ3SXOkzTj2fdX9Setmy31SbJbABoELq/C466pp+14izQzcjfICwT7RhgBtdeVYAtr+o6wBky5CbVJiuhlqd0jGDCx1hRBSJ3FlcGUW+Xvun19eDzlX94S+Z+GbS4DufPRAcnEuxzC+W5AOxVAtFZ13E6Q/m70gfOvL2bDyYzg//dxuCf/3Qh7Jr+h5J/2v6D460i0ZX/BTyohBpPEO7fGN7KJg+fElj577R5IgLwaQ2mbHfYamfGRdgqKJQZ66v3SfhMR68UscEOotTo4KA4KJYtkw4ji396vBRUoS78Go6dUIAyTCW/joH2V/CdyORqh8PxRejvyUPhoi6nWL8AGEcKw6kTPuXQwZW5YTHRQcviyp0VMC2QIslgRbPKZMzeiu+YXnN6F1ijS8S1Zm2U/fzEnX9ukY14TqdAWE3Y4un9L4P6Nj9Wv+wKjueSyr5KwA1yhBT4jsJok5t2yUHRn/1J1yBhkkyPvvHB+rZC9fqHCrHtP5eom2VrcY4kQOHEpcjwVrOt6IEH+wZ4ldRvvktmWs9UgEWjI0Y/7hQTToHoM3GhdRZrmcxL4qj9Q8EM50vB/eLkb4rKE1E78GtOs44sdYRH0V1PuN+vE3WSf5TermHtA3wSl02YxhO5Vvj2TYO43nss2+sup1feQl4CXgJeAlcDBLwgMXFUEo+j14CXgJeAl4CJgEmYbicM0GFT2D0+7tnd7/hUuaWfjnXEugh1LaJIEoxFPYoDNg2EkoLr8MkkbLoDQFgoQE4nxBQb1diMkoZWhxoCyllyh3uQTJrUzuv1wXhbNwRrJ70gge992E/igPiVaME4PnmKXK5tlFyM0mm7vGOWNwzYWbbLPi4H7+Nq8LACvOqQJb2fq7IPFjhxPCqLBV/BWVKeaHkQxkFeLZV7MXH5CFSkHNZphMXGxJ16gVlidKlKwv3VyW//iFeAieRgFkVUyepm3iAEcbl3Q5sq+qz4tVwC9rhm9WmSwkb0m6xFPoeYrw1vJTPvQR6+k/rY1bcXqrH9XhbuPKokmUmkweGWeeb0tWOQcy9Q1d8TZep/yxukBZ9RIUOGfOoQAdZ6SdCAFJZ7mcCGyDnxqI/dATGSiJ8JlSU+qmyPrh2TdtSTPeo+ZddE2C7FuABICLehKE4HLhjpFi3pRn8HcvQw3PF9758WEBFyXYt8CwEQFsQ2qEQSgSh6qoRHc+DPy6Kf3K/cv4/h0Xzs39Eu/pVMTdN5kV0s7wtunPR8KFDwYbnZ7pjL21u7kh1s3JcAXdC2R+XSu9SEX5Qf8l7v2AWPCyGiZAFVqNnwhJuMjVLewELJmq8IXrKveSG0P0KZDSusFDrI/FmpF2RmhfhDcJs9I0Vok4XXbkOEoZKPcZ1wne2wD2lRFiked2fPmNOxxm3kHfKMBRYsZyXCrjIPqF+6Nf2fe6QcvldXcv6awIvblW6UWDBVSrLDRpxiW1Ddyj9T3nHKSWedal+v1nX7NKaPL+g9de1H9cVhQZzYLzqhPaE0fY0mrg8i0cZd7llaPGrk2HWBWBI9K+jaykveC8UAqwC2Xhu6U0BmHVY+6k70y6vRrJtbxW5kGF4wkDQTYkRSmqT1qMO0CjH7o4HpZILb+TGirW7gqX0yeAH+XSwO1wIHivaCqeZB3dI1pDJDzV0R8l1XDXwerxPVEt/JM2Cx+SVsUdyBsAhfxaOE5DGxmPUF5J5Mr3sGzR5+LWXgJeAl4CXwNqTgAcs1l6Z+Bx5CXgJeAl4CZxYAkw6CM9DGALjPyBUj1/OsQR6QkCZdShjBibfTGoBLYzEkP0GYjAZZOII6bQjWVTiOEphLOTepHSTEp4VLL3eBr28FKY5Nq8OAzS45kyBil6gYPW1vd4a5JfwTxArf06JuNGEniB2NYk8886ANAAWTNwtPBCKDmfCqsSkmXtZqAbzHFnWAnmOiqr0L8zKFFe0JROq58QJv1plMqZtV0YVgLS6rphyGItfH/v/wpSdf+qxEqC+GqeKxbTnDCmXoSyQhlnavDLEmWu7tlVtD7Hdv121VyEgnkALD/qf+9plbc1Z31mABqCFhQ60/rD0PpSFvwr5eyruoypxeYChWKfPzaTkDTcIvFCYnpz6IQv4lH77GQEOu6W8XtR1Szq+4iG4AlKskECs5LoEKyrKiLhWi98wEmx651h266FusH+yFqz/8uHgi596qXiyLc8EuwzUQnl03phJXMzHhdw2wm4G7JBPSSf+mXlVzEwK6+JFeQNJma3H1OpBO4+LPa0tC/cXd83/yNCDmbLmPEtUhzVGKO9X9bPOw0j7eQ88RIbEIR6FUcXPgXV/2Q+LuNtZ/aPkd5iLQztU42nyS3yl3FXez4X/W6df6xwXDB4DUbBNJ+zXPrwK8C7gf58OMrZR3sIslJSlYJ9VKCm8Ange92tX/Qn9hoWGtDEJ5Zh+YoPjuzgqr4uHii8r9GQqgDyUUQdhoAKBFl1xRBQylugIDMDjoByJlV4QuYipF4Lbde4ByXWnjq3Xvhd1LuV9s/aN6LyuKDc2L/S/kTGYW/pbD3WT9OCVzpPDejqkjB8Ff0sIE/prSLzhxsATp+SECB1AtFh5W+CBUb5pCSeJJ736TS4jN24a13MGlCdAU9ohQKqGrudMx7kR9ovb4hb3+6DYWmbTR+V9Mi8gItUz82Bc4MSEym0wStz7b5BMBsTiQs6bKqMXXH6crF1d6fV8tTBQ5dtV4zQfDspqgl97CXgJeAmsbQl4wGJtl4/PnZeAl4CXgJfAsRJgWgTx3vur3QAX3mLqHNeSHstQs2hkim/xtBk7WBgoJqBMgkko97F028Gk0yaGWnMtSuE3Kl2lZAqNXgXZ8UAI9hkXBm9oXhFn+rYGInA/FAn23F6wBIABC8V7lT6tdF91HqAYChKuBaAAjMEaFUtB3hWFiCkKuZ9NlrmfkcG7d6sUhV4peKaldw7P7/GuoEzxrgCIurOqZwZULCsH006b8qKOU2+d1WxVDyhnv3gJXFAJADKoTqOoo11CMQs57TbaHnkGWSgVWX679oukuPvRlfK8QOH4xare08ZTz72XxQUtzRM/HKJuykjARe9Yh/Ki/4EEW/wTwXfUgNG3KuRXSPg6LNoh0qZ8m1rL4l4eFSj/40SBfuCmOFGEquPkxVwRpB2u5Wl020B4yS1D4S1LebAwmwbTD82HB3e14MfI4R/YpOeRN/pMFNMKURU0dQu1oYW8OAplqi2S7DAtiggwYVLXifcgDoO+Zr1opxvbncaGnYtXPC7985LiWimzsrkv/SF4H+o8gADjA+RAon3G2p53ZD8JIGefno9nJHxFeB2UuvVEQJ7IMHpxmp63pn/fp2NXBVnRJBqWnFX6s7TYIjCC5+zXNpIlrBbeCPLD0MeVRFGW5jXHt1GSnjMOIK/8xrOAsYOFjzQFuoX56srrIg1v+lxXYaIe1nmQbH9e68tUYnfqKji/btK7bFYaWA5EScgm/sXyukiUasFtOpfvG64Jwjr14ffQLi7L5gbfbZ6qwcTMH4rwXFkrv3pAB+7C1pL2AUpQl+DVwIgDQID80/8ZN8QKQGqjNxsBlXcsF4AiY14ptB2KWLwch9H/cg/rU8lJCSWtD9IkCV7InhX4c0TeFq1gTEDUG+RNcUMtDwbEENJqd50ny4DkDv9U5SkU0GFzPwCRjrJFBbf2jW3HXdGTuyqTfuUl4CXgJeAlsFYl4AGLtVoyPl9eAl4CXgJeAi+TgEI/5QoBJYvC5YXJioV38RJ7hRLoIZXs9Xbgrqa0Z4LJBJwJMZNwFAEoc7cqlSSP5X7ItI0MEbDiNiVc+/HEMK+Gk3lKmILNnnumXhUmCVPE9YIUVl+w7EP5QILMHQvCR5QAW3h/R16rhOKDfUx2mQyzjRz4DSiBLGwSbMoH4lg7A+cqIx6osBK5QOsKrKBcAdaI409YsmvjOGkQsr2q+y6MhLalREOZVnxf6x9o364qUU9aUhSfgabvAr2wf+zrQgKqi6nqNophvNpQFj/Bi6vu3i6y7Q2q22qrCizT3ZxP9T1I845Imh2ATPv1FG2a7rHk6/U5rzJmSX9O+oEe4IL+pwTHS26H0ouiBK6oC/Rp9MUcL0MSFgUKYpT8EyLcnhJAQMgoAAaIp3vBe3d65cho+V7pf0EXakXjJyejd6DHH4iD4Yfng4eeWRRPdp5LQR6KBFyx9KI40206QdppqSeEDFoAv0JP4d3hwAdX9/CuUOwy/U7q3aBWD4O2dnc6E3KDuK4b9H/712764uz9zzfzB+feknbEt1yBFtRp7pEop9oGUnB4M0p1tds60XFfu74ZOXGucS+IKFufQFYQQkoKbwc4rF64bq++oV26y2YBEf2AG4qsti7NG1tEEL5TsbZaovDIRWeP+1LkKEPEY55lru+AkLtPUaN0lciu5R0gEYuQ2+VP46JQXBlu/GCBnsgbZbgk0KKtMFGpvC3I80GBF4T4grx6p2T4gNLVunKb9k0pofyfcgGX+LrNNENhsQQHDK+wfSnWVf/GZK7v7dV7StOfPRhGA3qEfG10v5ZLofNS2as1+YSXgjqFlwVjHsZLJaMF/1aPyFabDfUet9FRyXUBgJHoDoq3qLIr5D0SVkBOGU6Ke8+FU8H+uBEcjo6IjPtAEGV7lK+WC311s4Q61qipTBOBK0T+UoFo/6DwtxEd6+rRcG0w+iKcGOVfQjFK3rPiZXXd7/AS8BLwEljTEvCAxZouHp85LwEvAS8BL4HjSMCs91E8o1TG9d0RM/rl7CVQKWyNrBBlB5Npm+ix38YMKBqYvLKgABlXKq3xSitGygTrTjwQmJTjBbOlOud0M2jTXZ57NovZ+pkVo5F2cy/yiUJnpxITc5TQWFRSr/Cy4D1R6AGGAb70clEYWGNWhqYIsSAIhGBZVmb70E9nU3Tn7RrKlfIEsKB8b1ed3+4q+IqZLSiT1E8wFrtwOs/rMOSe8JlgZTrj4/2ft/LxNz57CaCUpi1zYIUWhagprhIHy0YpUV3MfjOQJzyUqjbfwe2q31xjACzeGoAWHlw9+3I40ZWrvfpe0RMMuNBNHMAqzwv6ZMZD5v3Ib/pvC0+o4DmuBoh8WSwBWU6fNqGKQL8NQbcUyfIXkLvDMYRKvRWnyjEMFhP1sNEvHgF7ib88mD/83LwC+AShQgBFSsqGo8yQJ0Dm8IRRBWoak2p5vZ5BH8p4bUYZIrwSwIYorEUHwXWi3FAeGdOV3Apa7tyOPv9vbSzCLpFYfwBgoqzW4pLQpqnFu9pZenGukD0bBwOnz+k6kTsXGruE49rBuYQuKpeypLg3Y4JnJFYpwWv9c+1YuENjsK3QSu2877ooyA82oqUFpaXY0YWnWZJ3urGCQqn70D9dGYexbldX6hdi1NR+vPWGBZTIO8DF15IxhEJJlcAKzzNS6nmAC/3O5XGxOP3VwWcH86V9SZE9ofxtlcQud2vGVXBEdNSnZS6NS6nP2IvSh7KbAElRnvUFc6Pv4nmOmH3DwX8x21h87mhQcwYVKP1deSjBgSOQxgEXgBP0lZPampd8Mu1vOF+OCs2qJNYrt5cfsZGRmaAAWsCvwZK7gFQbdN9B3Zdx2ZC2KUfqZzMcUngupWhrcDRcFzxTPB3MyttiXhDsOgETSSLvHt3W1adI8IdjV8HbRUlvFuucVLIXgYuE/wfHgaWOeQH/w0vAS8BLwEtgLUrAAxZrsVR8nrwEvAS8BLwETiYBLPfhrSC+70eU/lBeF9/0xNtnV2kqLwCmk0zZDZhgQslEnnGCxf3lN+eh5GJyy1SU81GWGWDEJBpPipK8sbwnE9FXe7yB2sHCF/BsIwkHwLD6gyKaya69H8oC3gkQhnflHVAiEMbBeAsMqOA+7DMLTlOWoPA+Ruejc/xygSUgRSz1kPoIITHlSr3Fe0Yxyl/mLFGTZTpk21amKHRpbyhvHzbnApelf/zLJVCFhkKri8KRun2dmmrVX6fOxUNseamIuNlHODQUknwbeMoZSa2FsvOiPncSWG1/fu7urDsJwHB9mIALx4mgRD8FYGEeihbOEW+Aysp/2UMSI4MxAQl4Pwq4UHVwAK7ScXgtNjSC5i+sD2+2F3ipHez+xtHgJcV5Uh64Riv5QgSiqyjhBKUk6ZP2vhl0tT8XIhGGFrZHXo0hHheyrC9kJa+s15Xl8h5SuOdR7c9mkqyIVW0befDztWUw7WM3fd61xb/38PtxrtB2bO9t4xHaezO8QD7Ua/pykc5zpaidy31cJ48T990sLyIAb8kJYLc8Kq5ptQfXT3eGdXJ/1MnrE2mR3CjAYn8t7ByJldEkStt1gRfD8fThwXhuLizkZ6Ec5VKXF9Keswi8aMpTY724OtanebGkcQLfK8zdjI8YT5ErAA3yZB4NLYi6/6g8trC5e2jhfTP3vdgounBcKIyW69NqGoEN6DfjYVwo7nSq+S4E6wJLwmTo8OgvDx0c+UcyLMmL/tYPDtfTPfepg3vcBX8q2weAI4w1KBfkZ5xceKNQl8rxnUiv9RdQYTm0VK/Mjrvd62lBviyAVyUWSZ16V4a4Kr0r+DfqvEcgUy+9L/bHW4MjxZTAiiPBQ6ECVoUz8rqYEeTSchwWtF4tFeASNPMSuUODBFhQ1Of12zvl+/sTvAS8BLwEvARekQRebQXCK8qsv9hLwEvAS8BLwEugmlB9R2smaCw/qwSBqFcmnkH1qICKXs8Ds9BkAovSHiUWinsmlEyMOZeJK+dxHGUAMkcBgrUl8dONnJpzesm6z7fVrk2Fy5jZ5cSfSbXxDrBNXgEgIG2X5aQLnYHSwvJGfrnWwmEBZnA9AAeTeBaUGyvhOCqyzeoYq/P9nj2P8ptnIAHqrinwCNUl74ngklq9MdhFiVYp5qQ8Cmu1hmxlu5QjnjeUuxGod731+RlI3J/6qkqgCg1FG0eddcpZgW7zcVIbBKTIFAQeI3sAOnkQJVEYb8iy7lClMLXvIxG45+v5uSs5sys3DqNzd+fj3KnyvMDjwoAL+irK1votrjKVMf0bx2n/FMIp6gsa/TXiHjmwga4swQFA3SJAguqNYidFv7QhuuEdYyGKcbfcfaD4xlzq7r/ixmNAR8loLTW0i6dUem8k3FQGBGHYlKeHFNMZD5PCWmGpVEedejnP+pUnWd6Hk4oXNReFqfwEsnbxZ0ezTiqnhV8YWgEubv5Cr/dK/nuPfBDVN+8lz4awptvh5dDQmvafvr1U8pdPwpK/DJmlPCi3CjGlGFr54EQ7HBxa6DQHl7KBsBUOduRVUe9oeKBPqV56ijA2KmThX3TkYdGOw7xzINycDiYzL07UDuwejQ8dTsIuXgrLKnOJwbHJQAAuTgy8FfifC8RA6Y50NCYJZ7U2jxnjeUC60Yu1yfTfT76vu6F75PCbFp+YH84Wi9HOPIG3Ev17TiV9n+4vsFLyLTGnvk59W//s4Hvu0K93CUiZy6Lhe7N46JM6tlc1QZ4tlR9G+UxXikqUJ+Mhxn/iQamAn8KNmQjrxPgKsu4Vwm6DBWwU3gtU2Pbq0ZFdU4IU5HcFNCJneMrEenYkAKMbHBYx95FY5gbFRuW1FSzk+4JD+V55y8y596gJpciFlfGv9Kwo5RvUlOPOR1UhvJdFVcR+5SXgJeAlcPFIwAMWF09Z+Zx6CXgJeAl4CUgCFY/FJ7X5K5VAbnSTKA9YnLR+9PApcJ55UzBxR4HQ6+ZvBNtY32J9SVx0Jq5YBGLtBoDB+MHIDA3ouET7sMA73tiid/q6Op+909iTncd1lennshrAQBGUFOSPOO7GP2FKG9YoJlBAE6+d8D68B/diP9fZ4uJIK3E/syzE+pHJvCl+jKfCPDNWv4//vfYkgOIHAG6b0jrF67hcRpjrFftJ4SOq6odiTlqyNO1OS6l7UNojrNWxOqVOFB6sWHuF6nN0XAmgrKV9eybPs5rq8mZtjwmkgHTZhT+TWbc+gagvKqJr9RsyX4BZ+gHaObM69+J95RK4IAB2D3BBH2VejryNeUzSJ9LXlgYL8Djwu9tR2CYXQYdjKOa1F62vOFCE8d44HI69ZyK8y8Ty7GLx1LeO5nsFNVhwpvKQxR+jj1WT6tCysp0t+S3gznD8Gd0B501RjikISSVVubrXHALucKv2DaPc122UX4EqIulu1AR+fPZoW/vz6j2PKaWP3fTnDrRTyKhOiQEU8Fs4sBoIRuumtOP85t35VlDCsx6VJ0dzJh0fmk6nti7mA1tb+cDUQtY/0s37kiKST4WiXSGbuGjV9AtXEBlqhApFpCBFuYPBa628OZ7m9f6snjw3mhw+3IyW3PjCYTao0XmwCL9duCj9VP8Ti3tBdN3O22JI+0jKp9TwGpsor4tVmCTKkW9zcV9tfPFzI29BcAY+tcR5wfk7xXnxoNYqRzdma04PfWhqvv+u9/JcZW+gXd/+23vW/c4P19367zKdyz0paxsPuhdUYoyT6AjcI/R/hPmEwJsxEcfYB+DS5xgukJ8AA61J5Zhs1ajOlcVyZ+vOKJcK4NBxvT9kUtpnTo81x3bR51LXgSaQdsPY3hFkcjS+PFiILw3m8oMCLRYVdmtehTEjsGJOvxeCTAWfU5lj5UqMKn7xEvAS8BLwErgIJeABi4uw0HyWvQS8BLwEvASChyWD+5XuVHqHEpMzrOfPyaIQU9ynd/JWCCg5J/e+wDexyalZGjIJNI8EssZElAk200b2M1GF2BGPCibEKH7hpCC0DvfA+6AMqbBimXe+X5GppyPcrPLD85jiUmg7qzUhoFCCALYAusCn8ZjSA0p4VRjgYiGfuIcRX3Kcheewj/dj24i2XfACzb79FPh8l/S5uz/1gVBlWAa/U8ra6wspc7sdFS/KNcxbpTHSPtwtvqGyBdiibu9Woo5cEMXjuXt9f6fXiQRo3wFcdyqhIaT+AtS9U2TbV2cuGg/VHeVpR0rT5L1FltKH3qv0VSWL9V9azPvlXEnggrQfFiqKl5DXBYpk+i7z+iBPKMDpGwEUphXdSPTN8nwo+05xSMi1Ah8JKfObUdC8blAeD1jVV8sfv1R8Y9eSVMPulOMu6KnLUE1l7D2pkPO6gApFUqI7xd1A8ffgrICsu2qLtRtOA4A2wvdpHCIVdTkeMSMBZ1igd+pW7/iyhy+HjHrkg9T4KlyUuw99unlRUt95f/YNvdC6at0zS9eNdbL6evUH14RxtKWVNmKFgAqSWLGG5HgXaxgwKG7wKBdHdSh+mDCJxUEtzAJgR8zVWXPjkWCyryvei7SoPbW+vudFhY4Sr8ZKZCIkkVU85xV/EtB5fxRH/YpEOKHbTGm/PC1C8mbhN3lH8gsYyc3MIMNCYblvNnx30BYQsV9nHHj8iidGusmmX9feWyoBYdCxX2NZN3bRuQYNAF5QINzfQAzqhu1D3vShDILJE/Iz/jLOn9WdoP4eVwJUKCnF3UMotDBqR7U+BfZKxcPRpafliBw8ROtR5J0wUbyvMG4W3SXhESsxGs00pLwT5Y9BjHkLlePzWlCPNqqvTuUdsyiQYl41bFolsUs5UECr2HnsaLz2H3wfXpWIX3kJeAl4CVxUEvCAxUVVXD6zXgJeAl4CXgIr0yBHDGgLk6dzvXBPU9yUoRMuwmWVZ4WRaqOUwK2/Ugg4BQUKDFNq8N54H3A+k0QIqJkoMw0tY16Xk3y+Lzy5AAAgAElEQVTO5zzuY2GYzkRKPMeea4qUk11v1n88kwkrycJPMcFGufx9JSbVKKhRevBuHNtT5ZVrGP+QfyboAB3mWWHxm00p0xtaY9mjwpNpn0kRX9hzFeKG8ga4ukrpBqWtkcKS5J0yaDaKJDNDVuWa1fdyTwVYEOYMDwusz19GdHFh38o/3UvghBIwTzPaUxfWTHV6s7wtaA9VxaVyRoUr63mpC5M8c4DGtdW51PcX9c205VHk6/wrrGSlknptKEpR7EvBT/9p/Sx9Yhk+SVGQpOadEahwQEfr0i+jnN7sQkVVHpMbmsGmH58IbxOxw4LAi/6ZNDjyg07f4axGKCdHlO2AX7eYh4VcDnQ/PCNq1b7Sk3P5PH6pqxVmoX2ZUDSFfhJbt7T32kY5/qPK15AqKmEnW9VteQh9tuOQqsJfVQYFadb6mcljwCF5XJhXZv67j3zA9efKlI0Z0m/OvKc40p3Kullt7Eh38obZbOzdSdC5Io6LqajZTIJuS6hE3omKJKorOtVgOB0p+hPRnUJowoXHtAg9VYRREsp5RHKodYpobCYdvSrN40Y3rzU3N3c+uwJamJhWslnWE8EfEqW24yguhgSYyBMkGJFvSlshozo60NFpjFMspBVjUr51xkIKhfXTTrL8+4R23Dr8283B5JJf1OZHqvO47t8pMTZ62SLwgoVMAV6E+l1oTf0wgMBCI5p3CmOo6cr7Y0FnMi6EvLyvaIRxN0zqnTxpLOX14U5RG+oGwiPCUKHo8k5/3j6SSKbdMG4sRo1JwIokyFp9eWdax2aaRWcRcGP5yylrLaGoCBOlyGTE5qrCVIUKRxqpPsSqH0kwGw6qTIZF1I1/sGpd8bxQN2Aav3gJeAl4CXgJXJQS8IDFRVlsPtNeAl4CXgKvewkwifpTpQ9WkrhNXhG7zyHxNjNIAAsmgyguUVpedIsUVS7OjZvulYp9lLcACygDUEowieUY1mssdi7jAxL7OQ+FLyAFCge2AShQGJjlHdND7nn6ZIwrz0OJsGy1eQohm5milQdKFwAJM/Fkgk2+mKJybFeVJ97FJt68M9soPcyrgkm8xX7nHhZL2UCKzIMUpyiZNXi4Aivw/iFc2Qbqrb4J0b5SNZzCKNVvyrahqCULWv9Q6Qfa/4ISChgUZdQT702zBsvXZ+llEqBSo1jEO4i23oEW1Ok8y96g9UYXuIb47mFYl35YQVoK562m3wDTfCd41NEulkS7fnnNSKAKoVRIyU+9MI/B0ihDtu4VyQnHaPP4TT9fb0RB54ahcMP2vuDKdl7Wi+/PFfdOL3UOEWdIqu2S2N1RHJcea9VvVOiEN0LZXI1Ber0xdJ4QMy2QZGS6trwQACOMxHHRvUa/5nU/xiEiYHY311hBlMulAQV5of5WyvS43fjs0VQK8Lz7oZGXtdm/cdPnnUKeJAV/+Pu7fqt+MN20Xl/E9Y2odbvggjcJZHirPB36XEAhhRWqB4v7a0H7gMg92qO1+Y0T8cHJoXA6awUDYTtvdLI8Pqjr+qMoG46jolHEsTxIaklaxOPzCkaUd2OFj0rTqdr+Pf3JAuOlCrs51itFnhVObBSDXj+K46ghWKUhggv263t132RL3ytlUhlhhDPaD0E33Vmn8p9J6/GoYkz1wyf2G2VBuHHeZ5Q+pTGycVVUh16+Aqxw+SzXqYALvE7Nk8P4zDglnpeo9scj4UDeXqzLbUYeE3GaR4PtqD7Simrr5T0xlYbxsLCdeq42Rw1OdzFsHFQ8rHYqb55WWN/IO0u+862se0jAxq4oL14CtFgOEWUQW8l1UYUxA45wbZwI251sZnSkTykKRySvEVc3umrNFvUe3mPshKXtD3gJeAl4CaxtCXjAYm2Xj8+dl4CXgJeAl8DxJYAi+Vs9h/5Xbd+rdK6ABRToWOcbsTSk3hfNUgEV5tpvgEAZA7gEILCqRZFrRNoGVDARBnwA1EBxBTjBNhPDLdU292P8YETWABWAOqcLOvTK0YCU05WtTV3xrkFhwfsApJBP8sO7Qf6NchrFM14V7Ke+MNHnOJNXJrh4YxhQYd4WFjKDczxHxemWyho8T2CFgY7blD3qMnV9n9J6yFxLlYyCSKD0KgoUtYBb97rfKwTtKGrMEnkNvqXPkpfAigTgWVG9p+0CfKUvNHLhx7V9n9IHVOeJgwYQvy6SWlSeF9RvAF720T5exrbuswSRt5fva08CBlzozfC6WAneY0BD2ZfjnUP/Wr91KCz+7sbwdiQh34diuhvcs2Mp+NRSlgFsbFP7SfsKL0UprEKEDSyiJZDHgUI+sX1COdLPqr4qQlAY1RxvBvmAN0NODDo2rH20zzPV75K0u0wAF87TQok+nPWSQg61mncfSfM8ysRLUWQfXiHptlz802c/Kde67BIp/O/Ufd8j4OHt8mq4VCKRGnxA3hOCLjpz8wpb9MMkDr87Ee3ddePAd+6arO//0cFkbp1GB/lsOnT4xfb2vdPdqUURb0/Ug/ZUHvVNKRTUsC4P8rhvcD6vXfliKxnI8toDlyVP/3DFveTl8jDHFDAcri8q/EZSiBWxsF/7AdwHhdswfgOkAawox1CFlPOip9H24kC8GeToJm1fbk/Jg/TTIoSg/zvjhdBRAi0sPKaF44x21dcN7aytm9gfDW/sK7obBoPOllqeXi7AqE/gxHpl6hohNv3yfIjxHHHYS1ZknSiRx26oUFqOED2q4XcR1bN2JxlXfUn7i85MLUzbCh9l3jFlnu2X1adYdU4Pc34lZV1lbfWD8SFjvAPKO6CF9xg745L3F3gJeAl4CVx4CXjA4sKXgc+Bl4CXgJeAl8AZSgBPCnlUMBn5EyXc3t+kRFiLXhDjDO96zOkoN1HCM+Fj4n4xknovh3OoJnHOWlKpik/twjxxDkotJv5MfM3KFnBiq5JxQSAcFFuAHqYEYxvQg/XZgBXc00IznFidcWwpMulkIvq80tNKWImiLKGcsIgHbEG5gaLNTd6VmMRiFcia39zDPCtQ7JGYhKO4samw8VQc+3T/62KSgIU/Y6yL8haQ621Jrb6OWP5uwXK3JCCG6JW6fqUSoXOoC1xDfel4wu2Lqdhf93k1QBblLRxEcA5dI4Uh7aIUh1FDTkYQ/CoEDUbtUUMW5VfLAwOvIhJtH216XaBF5uv+a7s+GXF1FS7KXpa+nn7W8T19eH2wdWMj+AkOCrBIDneDz9w/W/xQ7SdjAQuxOKk2dMVzw4WTEjF1UsPDQj0ybW4VfG+ZlBu9uutz6X8XdL9F/WoGSQInhMCLTGMVeXnAb1H27VxQtut4j5Y8UuYNqXuEA7LKr0JFhktS9HeSMM+Su2dU1XPhB42g9b7+ovnZQ03RWmzX9b+sUE536V4TRVy/JOwbVGQiCCa6nSIP9wlreUqxqf4mTtL71ie7915afz7ury1d0mgWeAXE/e2ldaP9rXi6NfzA0c7Ig3PpWPNwe/S2dtF/TSPpNOqJ7h4kcsMY2TQXLm6c6Y7sGU6OzgBaVOHCSnlLAr2/S9wI0KY87MIW5o4Ind6qoWfX9KNPEaQaChfFeG6fzlnUGXkSNubX1e/c0Iwm/8AKUw4af360+/i3Hp373dMdZ72s0lfeFl3CRL3YWJc83Nw+Np33benEtZu7YfQG8YhfEufpaJJ3B2vi40iiYijJuuNJjAtOHvTJJ6UhOpM4KRKBLg1cJXSNw7QoVSFLirAVT3TD2lgnSPoloRkXUawCbUxOy+tKNpIRlcrqgfGcUNmQC/udd0jF0ZGb98jLXtDv8BLwEvAS8BJYkxLwgMWaLBafKS8BLwEvAS+B05AAk9xPKwFYsHxIIMb9AjPOpVUoCnlZ3QVfUXLu/Gtt6eGoYDJq0zi2USbgHYGynkk8v1HiA8T0eljwSkzsmOwR5/9HlFDcAgQY6SLnWEglC/vEvQBBXslyKqDDAAQXmkCJUCcQIkMmS6JM8JJgUgrownvZub3EmjwHYILzuMbCYXAu28al4Wz4fPinV1Kka+Za6jN13XkN6TvZoHK9Qlblo6lCgrMQCkp/pcBVOJLy+8AzB9AOJZgjoPdW5mumPH1GTkMClZcFFZz6i/cb9R9wmnrtQGdxV9Qh+wWw0PdQj+LaZoWH2lpZbtMG8t3QdxiQexpP9qdczBIQcAExt2sWlZY5rP75ZeHorcOhCBLKRUryRztFsGPnkgvRRB9L2DzaS7iUWbe1H5Jt+lxZvRdj+l0LIk5FCb/K0L3UzvM8PCgO6+kbFBBJgIWIuYtCIIUU8mEoTwJIuctb6A/jDojCzYiiDGfl8hHSn9PPzyv8UMtVcuVHmHQ3aLX6mn92ZErXbda+66Qt/+mgf/iqYHFWzw+jotMVn4eMGbLsOZHRP5IHdbnpFfeP1Q4//WNTX2gJHHhQYMFGYS+Xi4R7XVKL+kZrC5ubxczcOgEae9vbvr1/dtPMTDbSEVZxbV++0N+MWrByNBazgamZaGLdYG1uPgkzQhGuABUVjFARcFevEpqgBCxWsE6l4Ner6hN2XhW1NMv5vvuk+F8S8p6OJTcoT9d/SPuWw3Me7T7xez+c+/cdPbKhUFh80yvq/qpcP3bT52zfCauxrk0+UehZRT4hGV6h0r8dDxWhMrcK51kfxjUBKc2sXgvihuAHcY3zoLxepArDKG+IYiltRHJ8yXSFUFNwipoEpWsTAItI4aIo41zcOkA6DopYnSuDXPCqkMeG49Ao91H3LLSpeUVyNUAX/bszPhBwkXnQ4oRF7A94CXgJeAmsOQl4wGLNFYnPkJeAl4CXgJfA6UhAwEQmgOKBnnN/Wdv/UqmM6fvKFibE/1AJq+uvK51Ksf7KnnaWV1dgRa+XAhM0pnn077wDSirjnmCiyqQOq1sUs6bcZ3LHPQBnblW6RYkQS0bAzXGU/bjcm6fCWVvqnear2lTV3oUJJ2DFI0oPKRGKgoko5YNywkKasA8ZcK6FwiL/gBmsUWYYWGHhn+xZDqw4zfz509awBGQZTt1FkQPotk3pPUp3KQ11OzjXlEuJhgmsKFz9oA49VyW2j3qwYg0Xss/aCSVQEWYv6DtAmUyb/awSoZ60XShmv9tXfgNSIKflN/E2Jb6XLyih3OObIEwUbb9fXgcSALSgSlQp/9X7Z/L3ToR3yhKesZVb9nWC3/zCweJJkW7Tj3IuKEdFeu3GCIAP7EvVuBLOCeOH8aBWl0eEhh+phiF4Wyx7WbhWGLZp6tte4QaMT0RpIG5sxiihKJTdsuJxUGWFZzHOsVBmeIUaWMH4YFaVWxpzh4gICJF5P0AFvGdh+CPKS3+Q1BWCSIeTeqI8LQXpwkE9/xk96x4BK9/S9lPdonHk7278uBsjwQWjz4Vx1FAnzd+vV9re6mRyBCm2K3tHNjZ2fa8YCv7sy9M/972dc1s/0kyW7hitz4xN1fYEtbAxMheOCoypvxCFrVQKeoE/8ilAJr2mJiboUrZu/OOYO2w/CADXrjB0cDUyK4Q9xlONO+5sRhP0d26ZTZ/5P3YsfG62my8yVhIvxLJXqxl2sIbTw3mYrgYufvMvfiwZ29CfJA2RVZRjrk1y9rhGKMGtCpV1U5iEl4tzYzLr4vGiguuL4+6SmMKXFBhLjiBJnk0r3lN3IZRbRpHtF15BCK8hBeqa0++FpJM28rCmEI1RvZl3DjSC7kGF1+oIPgKOWKmNq0ec5W/yzBZAhckL4xzzHOYcxrm2OP6Snt9+00vAS8BLwEtgjUvAAxZrvIB89rwEvAS8BLwETioBwAks7gnjwqTtnQIx/vQckG9jkfoGJZQ8D1cToDVVFBVYwWQN5Sz9uSnombAxuWSiT2KSacexmjVrW85hQmwcEIQM4X3tfN7XeDBsAni+gQrzeCAcBUoz8oa1L0qCHUqE5+JdKGsW3pl9Fq8YZQmTV85BycDvkqdghYvALBeXrQy9R0UlzdfAquKu4BsAlCNMHJwml8dJMqqwN05/VRrjKuC3TF9zmZZr33e07/vaSZgx57njwYrXQGXwr2ChfQB6afeeV11/l8KiXUlYNL4Ds+pOajVIuPEmLImOy/ZyWt9TuwJAvDRfZxL46KaQ/vd/6n3tbhE8/fWjBYBESX5cAlokKhTjDRrXQ9puqYntFx4sS/9wv1AxkSTH4wIwABosrKTIuOG5AIwo6KvlDcH1rmvGawIlO/3/ikp/hdAbTX9T55AHNPiMVbjevOoAO6rGHkN8gXRhpDFO/naFqboyiOUMEIaDQbeta9MZARSPKg/ivcof0/o+hYx6Pojrc62fHSs+phtLoY8lP14Wzyp3X9KujVmWj+r3aFKPG912vlVuIbde2rdz7yULOx/YuXjFiHwGJpIwua3ZmdEAJh5cygb6NjT3dCaTxQ6k942+msQivXzuPPziSPG2XPgnARLwkPWGiVredrhNOXRxHNQsOlOeUuG62m2bFQ7Khe5i0Yt197bubc9nOwTUFEM6EyCHb5vnGUeXhcR0nqb/5tEPhd1uV0TqAi/DcEyU4YPK35vyPF8vCOGofCO26bGXSZ4bdGydnj1ClxpJnN2OoIxusU/Zx7+ileXR7noR7I6DdFYxuOp6s3ZUZK1m0RWzSNGOgqyoi+NCfBWqE2GjL28XfUV7pq/oTMd51gpzwoppLGej0PKlyqUciQqEcltWn3gryLhJXMU7leBZuV2iY3+jPxWxuMnKr70EvAS8BLwE1qYEPGCxNsvF58pLwEvAS8BL4PQkwETkG0oAFiy/pXR3NTk5vTsc/yyUNSjvWe5QQgG6VhcDLFDUG7G2ucdzjLwziecYnhMoIczCljXKfxQDABl4WZhnBe9rgIi52tu+VyKL3ilnaeReLmybN8RObWNxicKZMoZPYG+1jdcIAAUgBpNQJqucA3jF5JSxjcUvZnLuQvtwDsBED9DDZN8TMb6Sklyb11L3UYqhPKOuU6+Hjg23gX5sGXtDeYRnxYNKsq519agiuVibL+hz5SVwmhJAMUkbCBDnFJOq6zer4cPqvQe8K7e18O3QB2CVDHBNv4GSc8Ut6TQf7E+7eCUgow8yTwMJcfP7et7kj7c1gwNHuq6/pZ+1sQJ9sZG9s5/wTosCJ+ZVsQAV5DEB30UKufaw+11eP6Ref6D0tgjV9xc6rjBPec41ABmlVX8YUg8xOjjWA5Jz5FbgdkPW7e7reDUaDgQRKOBAlKJg3DOl+GfrFPDxSnlUjIgnQ628mvlOe1Zv+pTO+ZqOf1vXPyvXhx2tn1t/TGhReR64T+Zf3f8TC7Va7QFhBFvl5bBO1749kSo+7bhv5s36jhbeM3532M3jxx9vvflZKe3f0Mr6oqVosH8pGx1/cWlbvb9verY/aRcu1JMuVfbxRqkLEJBy3oXScip63cvxczgMx7ort1n9cK9Y4jtFFskFYrMZcgBWpHu6X/qLg537G0GUbRN5zZzuL16IgnHVUnWdEJ1CXlji+9DzBUo0lAYVb2pK510uQGJjvS8eby9kP65Hro/r4S5xaSi0YjDK9SEM7HnQSlvZwVzhtwReHEw7CqdFfsJ4LguDJ+Xisrcv7x4Z7c4v9WXtxki2GG7vvLSYC2JphfVmrUibjaJbU4yoZkv8FfU8TRVCSu41qjf04aK6cPWvF6VZqZCu4lSgRa8XNGNeM1yhDTTjFRtvcp33tOj5sP2ml4CXgJfAWpWAByzWasn4fHkJeAl4CXgJnFICFfn2f9GJf786GWtqyJdfOOXFJz+hNwwGyp2wmsT3XhXp+RdS4W1gAhM1AyOYNDPJh5AcRRWaB5S2KHCxON+qxESQyT9KBs7Hk4R9Bnac77GBWfYxGe/12GA/4Z12KaFgY5uyJDwPIU04znugTCbUCfsBI9jHu7CQd8qOSTn7ULQtx2E3vg8PVFTSem2uqAOAFZQ93hJwshxXOSHvCuoUdQhFD98NQJhZl782pePf6nUjAXlGZPKQoD2knQWIALwTF66Cy5dt5WqPOb4HA3/3Vd9Ef+Vlcayy+HUjxdfti1I/3t/z9rST/1YJ5a8F6zElMb8dR4CSgRhwR+DhwBiE9pj+Hm9I6hXnM97QeKTYol9JEMdzOnd3kKaXB0VXnqDynBCxtfgkJrSfcE+AydbPl9mCDwOSbMMxSnU0z6nGM6HqfLRVqv+tOne9AAkBH9Kyy6lOxNq57g1IIs/N8D4947tKT2r7cJBEUfPuI+7dsjzOuz+LPUe5/NM7/1vxfz/0U+onQtnpa2wVBnfh4SDPAwCHazTGuCIJ07veN/Wnn9z74rZDC+3hI3kcT4R9fWGa1SZ3ty/fOBofOLAtef5g3s351oyDAXk3dQ/GM326o5wQTveTE5mIeK4VDuo2y+eB9nfufXHxnmfzsCtHwnA0joORtFtMKGH8ISwh6NPd5QETPCb5CG8IrqvKCS+rG/VOfUk9Gmk0k/XdloAM3FkGkyvbS5mcJFRg9TjotiTELH9e59+r9IDutSNL1X+GwazuT/8biq5iXs9ZUvinYCo7Gq3vHo3lQSHS9KDWDDs11ZCmPFOoH/06Zx8oTVV+CB3wqTSugbGiZLUQALMstdKQZsXsBeCHto12rZenjCtKnpVyKeRlEXovC6stfu0l4CXgJbB2JXC+lRJr9819zrwEvAS8BLwEXisS6OWx4J0IC/WfzzYslK5lsoOFvi33aAPlee9iE6DzBlhUk9XSgsxiJKAAcLMtZx5ungQAEngdoJBiklcSX5aTMya/TOpQGjCBA7TAcpZjgAHEdGafKXQ5t9dSbbVCa5UYzugnsiJfKISZqPcSgnMj8o1lHEoNABXygccEYAXheoyPg/eQkiFgosyk2Pg2uKfdH+UJv13yIZ/OqJwu9pNNYUXdAfzq1/cyKEXIMe8VKxxUlnV3qG58r6qTKEf4DlIfAudirwI+/z0S6I3bTp/xmL6HedX7N0dxLCVr2YVJZUm/wnGsp2l/Af3pP2iTl/sgL9nXhQToe+lXf77nbT+ibUKLFRVBdw9SsBxiiP7Wxg9SMLvhA2MPYvG5sD/aNt2DhethPDKoCihj/HCPbr9L60F5QIjXQI+I5B1RFFKmF+KlCvc5e/plD4OeNn2Z6EFeFTYWKopNys0WBSxSKCrV5SgRVbWy19UwIcsWdV9AkAeVz8e1xsiBvAFc6yQRh+vMCI363UcdQFNxfAT/+Ja/KD7+4M/sCZPsK8rN1m4rfbdAgasUyqkfOozOUnZdFKQ/fkXf49OPL962az6YGAuzehK3Zgf2BZuuH46vfmZr33NP6loRlDtuDGfxT2glPYax51btGq014kj03M77ie+zXELoqKvNUhBx2Iw3Nt62TdwVjOfccrT75O52flheD4GAD7wnwobyN6b7Uq6TetSU7jMi4uyfUj4UIS5P9DwdD8bFRzFZa6p1iKMamH5zQOBEG66bfF5gRSTPkiPaflp56ujaXcrFt+hHBV7sFUVJvjCXtn/7vV/KP/GDn4l/7ca7l40FCMVUyrYMJxaXJO0AEi4cmIoWYnXqFddQjozjADf4LSJ3N4aV94zqS+TAltL/ogwGRoKI3OoXAjMPXMqUsSL3Zh9rHxrKKotfewl4CXgJrGEJeMBiDReOz5qXgJeAl4CXwKklIGBiQSDDP9GZ/7o6+z9q/RklFONnszCJemPPhX+pbSwHVy+na/52xnmowAoLDcD1TqtUKZRMsc8kDItZiFIBKwxsYOqGxTj7CKWAhS2TNfIL8MIkF5ACy3PADhbzKOmNFnzG+T7FBQZY8CxTbFioLX4jY5TMWACSR5RlWGPCUfLD6n0cuaQS4aEANlAqlFZ35UTUQkCxn/MyD1ac62Jcu/eTJbhxrZiywtV1RZ9YDgll5phRLLvOPKQOKW65qz/US/P+Wbsv6XPmJXBmEuBbMEUdStk5tYn0B3cq7r0syEve2orbRbHfw/X6Qb9hFsr2TR1r3X5mefBnX1wSYGxxpxJjC1ue0May4UYPQbc7LqW+9ek9wYvcIa6B38KRVStxb+oUFW9a+1FYT9IYay1y7OAJ7RsXsDAZ4AAXJQPyhpCXRPSC9ktBXhBmyjgYUFkTJIlxC7wFGk/kjHsu1fUaK8jDIi/koSElNqfkquyRwkBG8bxU9IwtnpHa/AXdb0mJ8EN8C5XBh/tGFmQjonyLsFtXV8BFwLv/+q13d37vkfcL/Av/ozwQInkkKHSVG3OFopMg1NVbL+t/5vmD2eb42e4tgmPqQa3TTdIo3PJie1tN3xtgukAa8XGXPBwK16Y3zgsMOUS0LbeHPB8W2ICnxbIRicNlygGiAxH1+hHeFeP1m+Ceccve9j33HOjed1RnjAiP7C8y58Eg2YgFOwQ0UlinOJjQvQbVD46A4WhZlIj66RezLs4xYSdPi/bCTCdu9EUAB4fTTrFbIIW8MaJd4u/4pmTZ1rvSpjjup398618cEzquF6xwkn23e471sd0KwDBuCfaTTzMCQkfF+FB1x40Xy7BOAl+quwBclGAIdUByElwBYKGOHYDMeWQgJ+N04x0sdNm5NMQxsfu1l4CXgJeAl8B5kIAHLM6DUP0tvQS8BLwEvARedQn8f3qiARb0bX9H6U/PMhcoLz/Ycy0x7Y+JZ1wd6/VEOMtHnfAy7m0hO5ziXQkLcKzvLLY4k3+8JAAt2I9VrHkvEEKBcE/cQ2EOnDcDE1qUBdznsmqbe/fGoz7X77H6fkzMmZTaO/GebANS7FTCqheLTCPmxJMCfgGUC5yDlwXvYJZzTJAJ4+MsFJUcV0X1u9cC9Hy/l7//2pAA3y4KMJQTfBe3Kl2eJPVGilVtz1KBgvY9Uceof3xDPrb1aZSlwCE7y0LTHSNe/eD7MwDUvnM7t/fbtGO9ALAp2bmneZnZdn4yDxhI13X8vIHJpyGaNXUKspBMaBcJE4hF+RVKAL8l2fHy4rZlVp1Mytz6Bm0TIgYvNspqQPfoes+jNVW05yUzMv6gj96m9H/2POBPtE1ffMKlAm7FaTEAACAASURBVDCcslmK/eVvtfp+e3kEaGONY8us6Wmc2Ue/LiV+cYmYp2VQoTqJZwFK9ii+ShuJyBrwwhChtxIAhnlFFAVjA41rCoEGAkHiZFQK9boQOSmxdZMcD460pdGBOCuKFwRoPCmwgtBOYr4WIFLoujBkrEd7RD7IE2MOXob+ZJmoGuCC9/3YTV9IP/7wB57SdZ/XcRToPwtY0eh3nhGTw+nc6PjSviJvZ3FHw5Y8GlFWwnQ6nYRDQu/hxmKM0UgOxKkMLOiPlhQwSiThGu8VChEFJBI5/wOHLZYUHdLGR2PNqwY/ctdIchWhPYNuPrewa/Ev07zo3sw9dI6AiXCLgAsBIuL3EP9EWSaFPCjimkARoR6R4jPF/fKayDsdoUTyZGgvpYRT7HK9+Dkek4/HE9qPochBnW5hOpGXMxoRx8fZ8j5xHXUCgwHuV3KQlDInMXZlMQCDhopzS24dvC46rsxGJMEBwRORcoQ3ho2ZuR/J8YGU774MmPl+ohKKX3kJeAl4CaxVCXjAYq2WjM+Xl4CXgJeAl8CZSEDhAoLfUPrd6qKf18T7bnlfHA9oONV9sciyicyXtU3IqdUTG5ton+pepzzeE/qJc43XwSZV7OPZKFYJ9wQIgRWfc+tXArRgAsoED4s9Jn7mQQGYwbugoGLShzcFEzfW3MO8G1Z7VZjC1gAZs0YzJePZemFwHcpkkyVrJrtMfgFVXlICfMBiD+UDoAUTZJQGKNzIF8oDRx6rRNky2WVS60I2KFke3bb3rpAUXicLimq9KvWcb4U61NC3hSdRk5AblQW5I9uGzlWKGqvX1KudSiiQOq83ZXclN2pJoXdfri3ab9+5Bd0orZjL9sWF8KgS35qFp6ON4rgplPg++Y5po/h2aadol1A0Wrx7AEi+Yb5/2rPS0rr8no08nfsbONlR3vjOXViRnmTtAQp6tl0b0Fue9q6vtzIGaNC7W3g92n6nHHWhZsrvodSCRi46DRbdKDnpX7Cq51zKD0t572UhIbzGF9rPtyvhgclCu4gxCN/oaS093hfL4yYp+U3hT32y73mFDLkk4uacGVXGhwQiXKOKuU0ODwIpVAfDcIPAiz4d2yww4oh+E9JJaulM9yLclMZHIeOiCBJvtVWFQglRsdHI40GRA9i9pG1CS+3XuZBNq31SzKdIDNxFynuTN4UaUiwq7o8XZyFjidCNQaj7Nu4oKo+S/NdvHm19/OGffkCXAEK8JG+Lm+SxcKVytqU/XmxONI8EAwtHi3ZbjiJZGMvBY3hdsvuOQ+2pRyfrh55TTjEugTeC/B3U1+i4xXS9+jInPtq6pjaH5VfCN+s4ROKa3CqieGhD7Y3XjNduxBvGLS+2/9tcJ5iWcUrR0L1pB/sUCmpEIavkneAgj5o+c9fKypuDqFtZHoowOwyW8J3QelbvsVvHDioPeGN19cxD2t6rY7sF9CiP5DV0qFRVlvI2+Wn6B4ALy8op15XHBS+Jt4VxT1g/Qx9iHGXUDfoJkbG7PohrFrStcnWgBZ42QoMks9SBF7RVABo2NjTeFa41b7NT5s+f4CXgJeAl4CVw4SXgAYsLXwY+B14CXgJeAl4Cr1ACAiYyARRYARpg8TPafrf2/dVZcFkwoZE1n1verLRVaVr3WZ3Lc2WJbeCETeR5DhOyXoUhIAMghYV/YhulPqCDCyGgRHgbAAHuwzHOQQGIpSxrFH4cX+0ZYpZnplwwF30md73Wz+aq32vxvFomvcDOarf73hBX9o4oArDkA2xhm4kmhNp4ihhg0Rvay0i0WZvS001GS5204/YgnIG3nFtdMq/939RjFOZ8I4nqwnYpYK+S8inOZapKmPBSKavTgCuydLf2AZRR/0hHLjYL8gpUWO294EKFVMm23WfR8z3bb7Ps5RhKbdvfa5Ha2w5wvlMw2ffHN6eLpSwMkTsx1Glj+CZRGLGm4UT5DSDB9vVKfOcopMg7bRtAJXHksfynHDmXhTaAtotn0j68oOcdVrlxLW2fWc+SLwORzULagZd4BmhNW73cpmqf4yqp9vOcXpnZb9Z2DdsWysQp5uzaXpCnyvNaXdFmAgDT1mIt/3iWpdcoLJTCzpRNO99HnikcTBQplE5+vV7+Kcna4skDInnAYq2W7jnIV8Xfxdjnf+u5HeOqZ85iHHVMjgRiuHZDin6+xyrs0jHAp4W0BGB4UOcAbH5IBA1jQSENO6GhIhTSufYXh9Tjiy1BHAgunJILc4RCW6GfRKqNQp5QZ1mHyiyldcGYQlwL4Q6l0uiBTiGHc7tyVVCl17kCO/QM9hW5vheFZwpDxlcGuJZW/eX37zguAC7+2fOubfr6v9j+93dm3fQOPfltus+b4mzx6rHk8NBofDicbY/qZRsioEiGBpLFN4e1+mIRxiKqTq/Utch8p8CKHXqy2kIXkq1f3x5tKWmjvs1J2j0dnxesSGikdYrgNDmaXO/Gqp18NlvKX8qns0cnwyhPZK4hXKccghEZSf4ZdHxOLHqnTOCEPn8FfSqKGWVsWq4dAiok6Tg8LBHuiPMw63YdCKP2VlBR4dpywAvCe1GW5KsM2VS2n66dFXDRazTinn86IEYPeOGAcAEYPM+F5VIyDgrjQGFMSJtPuCh52lScaKLbUMnQPi9qH+dQRvQhtPUWrmp5TOtJt13x+MVLwEvAS2BNS8ADFmu6eHzmvAS8BLwEvATOQAIo7P+F0v9eXfNbWn9NyfgZTvdW9I03VSejYDtty8LTfcCq88yizBRwTNiY/JlHAnnAUpwQN4AQJM7lvZg0mgU0EzOsZ03JxyQbJaKBFEz6TmcxBR/nmkUakz2LZX469zjeOeYBYQAJci0JOQMX+oA1IQGY/FOWTIJZG2BhVnIWXsKBFppQG5DigYqzLZnXxnUoM/g2rlUi/NlPShn7XgET9SxdcbRKaooA0mlTlwgZd6/SC0ootDIU9hdaAV15ATgAgWI5Xn6qc+x75Hs3xbqBl1zLO5oiHgFwvnmPWZtTKvlWQqpxnPaC+5glKtcZAMH3SvtgwAX353xkvl0JJSNtEAnwiPvZ/fH+ok1CQWdhVrg3YAbfOHHQKUOSgQnspz2gXQDEAIiFzwbFu70D9+D9sZCmrUTZZ20C9yLvtDW0lwa20ob0Wkzrp7sH+7iv3dNkzDHjArLQNY6LB28Pymh13ekBf1wZrBGvDvL8mBIeSMjxo4qW9mbFf+H93UKY/zipXZflHYAk5EY4Ps7frXea13ucK6B++Zl+Y81IgO/+f1TCSMMW+MDO2RioIuw2bwvjFTClNG1JzYVrynOFWCrwHBgLGtotIK3ktNDnFycT4qAomailYQ8SNTNZF0TaMVq4pXRd1X0L2o2nNTjAkxNg1AwyyvOWGax1ujCMnn1lfxIKvCty2iGAPvoJG7NYe8DaKdk/c/Cjez80+QdfjcMUr5Q99aj1C2P1mZtHatNBU2zU8/GoMtQIsmRgfb0ZfVg5+Snn1VBm+jalef0gj/LsKGgr1wlGyZQzCKZHeFWRXk/rxWeTpLaxFg73N8P1TpdTj4bjfd17o7YcSSqv3aDbyRX1SvhNTTfpAMAESVyPEoV+Oirp8E4dgR/P6v4aZznPjkV9/i09seN4MvQ4wRwDcRIVugZ+iFk8PKoxF+2khVCknec3AnR8H0o23gsEYhSnA1qUwl9erP+xNe04ZWKLlbTVpbIOQbodunyV3Cll30JerD80sNkbtawSuP/pJeAl4CWwFiXgAYu1WCo+T14CXgJeAl4CZywBWQDmshD8fV1ogAWWZ8Q4+frp3qyyMHx3z/lY/aI0Py9L5REAKIDSkcSkr5eHgYkgijjzmEAhy0R22cJP20y8mMihIHSTXCUUDoAVFgaK/K/2eFj9TstK0urcXu8Ks8S2kFWrrzWLblMUHi9sFPdncm9xoZlQkphQYr2LnFFk8v6m0DSPCgsdYWFoHGjRC1aclwLyN70oJFCRbaNsA9QDbLxGwfivE2DRRAFLVBA8LCJpfwRgoMzAcvw+rQl5Y4rrV10RWym1e78p46lBceesVnUO34yBBAYAUC723fPN870BPvDdl2FVym+L75/QWM9BoqptC7HEuWwDFphC3wAfvBy4h1mo0o5wDEUd8kJ+FmJug+4L2GjtEvekvSKx3QuGoMhqShneFEcCbZUDZcWZEMvUl/bNwknZNbQlfP/kw9qJBZXpAXkE0FaggCSMCse5F4AJoVWQJwAHylALl2eh5zgXuQJscE9rb9jvFHiS1Sa9EzJAOcm5ACAkFIkoP5E15yIH8hiqjJxCrPLmYBv5IjMDexZ1jOcZgOQ8Pl5lcMxALPKOQpXQLzerLLZpe72+jdhFz9EPLTX5zWxW0PyfkawBkrB4py+k7T5TA4Dyjn5Z0xLQ2Id6/Xalf9ST0Y9r++Gqnp+z/FegBVXN+nMjVeabLUNVRtEjaqw/JeDizqCbXe48EQpCQtEmpDgNNIPmAPwUK14SzjOC26qtC6MD+lL36zeA24taE0ZqhWdhGaiw1+rVXzv8VziCwlEpWlTQbRFuiHaOvM1XIAffs/GGOfDi+3NvWlKa+c1tH3t8KJ5BoHOLrdp7F9LBNws6GJf7QqRYTsFcNhpNd8abE8NHmomiNClkk/CWXEB6Nq4GYkOtEV0q3wf1XSLBTmSQoRBXgBWRHBvCbiw+i2CyFjfqfXI+6YtpestlOn00zOM2Qa4I99SVaBT4UKThWTGve+FpsiiSiwW9C6GUlP9wVqfiQYHcFW6KvsDJwTxV///23jxYszOv73vf97739t5Sa50ZSSPNvs8wg4HAgDEUOA4eYMAhgFPYhQsbyqHKxDblpJJKxUnAGwU4qVRBErwUmD+IzZJAoAqzw+BZQMxgZjSj0ag1u0YaSS2pl3vvu+T7ec753T591d3qbVp97/0c6en3vec9y3M+Z3ue3/f5/X750kBROPYjhIzLIsfwasizEuHj8xFdHsv89QgbeGC0s9eXahcuI1qUsHDJHhfxsiivtrpOysOrBJF6d571JIxjSfbNfsvrrsKJNt+S/reF3hVbl41fJCABCdzQBBQsbujTY+UkIAEJSOAyCWD4/pcp352CMe5fpSP+uogZlxrKAkPTDw72ec1GF9aot77TVOFZKjYvBjSMfHT0agRfhUshzAq90ko+WJ3HykeBURLjYIUPwBuDkc5ss7wZLhUj267R09Xxox7lxXEh0WOrY9rvqMSPsgKU8RFDImF4jqdgKKUTjLGCZLD8hjGNDiYGAIyJ5crfEjumbHV6+++Xelwut7sJcK1y/TNhKH77dHXfvo0z3cBgxIruMyNNZ7Nn8zfXG8Znrjeu7/nlhIMaJJxum+33e74Rm3Wf16j9WpbPMrbUb1zbLfxHyp15XpB7g/ohPtQIZwz7JVCU1xPeDKzLMwCxpp4hrMOzgNAiH8gnxmbuYwxviAMY4VmXfXCv8Te/lccD+8XAd1+/T/bHdng+sT7LvnrfgUO3tMStCEMtJ0JnNOS/zvbVDIi9qSiGuVlvM+xi1mfgdDeqOSY5jIJnl28zR4cQDzhv7RymTGPwWz8Tm9tyyXPkkRSeG2wUgRrBgucKIb6oP6x4DvLsYFkYMCFsYXCsMHQYNREk9mU/r8wnz8/j/XolwLDNj6ZwjjBUVk6OCm+DiNJGMafclPodzbb4zjsJ8QNxpc5/O+g+F0cTL/p6DQ1051xPJW5caR6OPvl2GfpaOJuUh3M+PpN63h7GK0sMopk528TeuzJZ27f/i9bPnKKu74FNSvPsIxTZ5dwv/bH5cWMT4Lr+nkEVud5/KIX76ZpPfZ6L2m6JaRsJscS7n/tmI54UP5MHxvvi+fBlEQ++JrfJnc0FCF1tMj2ah8cdsfKvoEJn+U5wRpQYL3Lvj/GI4L7O82p8Ihc2yby7/ZXZujPL93Xon1Htr745gxiykVsaF4jxmGcJ9eq8sJYx/rPt7hnNs4DnDd9P/dDxH2eZj/xXd//Pjz747Gs//9Tslrtmo4S0QsjMs/LpjcPrjz5908aLkz7i4P45YkRE28WBfOY2HK/F8H8LdV3ME9+IPS2X83g4LOeRAyJmLKbTyBzrhxe37n87z/o2PXDqJzafPP3gfJJgiNQxfhsRd1teihNx4ngyj86IseMnkgeDZ9E0UZ34m2dgTS22X8+jAxWpZJ765n+ShfPr4dSw5fpInajtyTi8PJpK78t+nswxtDw3WXAzx1HPr6rjVt4jPC6A/HxeF32YqK4miMl9novMbwNj8ncJI92Amu5UVnu1vIPbYJdaZ3C8fpWABCQggR1AQMFiB5wkqygBCUhAApdGIMLEZgSKf5qlESyYXpby5pQWnP0SJoxbFQ7q1/P9Z+jsXMJ6512kFynoRg0Nlbx7K5RTeVfUKF7+rrAodOpek/LFKXTQ6HwTCuUVKc2omUIYAQyVGBH5LNf88ta4kqoPE2Oz/oVEivNtG+NddVDLK4LjwKhIR5lOPSFJMBgzv0JbYQjFgFYu/xxvjWSmE1yj44bG4fMZiK/keF1n5xMobyCM2BiG3tHfH+ceWWew6i3oTSDkem2jS/t8EBcMw8SKg1BMbWR9f42WKFihMGp+G6bbX+M8V6hX5VxgnQotVJ4dXP/cewiUb0pBOMDIXQlEuXe49zHMsy2MZBjGEDPLaI+xHU8DPARKfMQK9o0ZKc+oeraH0IDIWfluykhewkmxLG+puqc5HupW92YLlxSD9kCYgNL5phIvBr+V8bCfxej+s1N/a2+tdtb5ZYajSLcuLO7t68OMyruxvZ71PCKXz/CY+M45w8iIeIWh9JVhdSisOLZK3I0IgTcHz22eVyWK8Myt4c08296fwjMP9jx/YczyhF6qc1EGNv7ensCc88++OM8t3FTPox3sIFQY9eB6LSh1PZ+TYLxft32UyNHP45rh+CoHUgd72/lgFkJUJjwrfieliXu9NxP1H56w4e78vsMIpM3Etcj98c5B1X8g3xHxrusUIWMR0YL7CAU0OSjGeHg8FIv57+XzVfn7pVyt+ftI4hylHbRM2KbmLcCzjVw63DtpK2VdGmArK+SxiPUfq/vwluGwnq9ps9XE6O7f5HvpVNmWyPtw9sU9zv1E26wGn/C85j7e/KlP//31/eNTHzw5P/wf5pMDeS6M7xttnB6dGa89dmpx+HPz5cojs/X1yALLW7PVt+07tHqU9Bvrp2Yn4nXRnrsb6yQJ54jJQTF6dra5fGp1cXhyy+rbXn/n2lfwnEn+iqc2T2w++AgHuZiPSY6d3BPt+YFIizfFGmsnPNR6ImmRpLrTlEu4OfcM10GfhdPNYf/sD2GA8FBxGBntm65Obg6HV8Q75GR8NPIeGh/P4seT2PuJiBg873jP0K5jK5zXSlx+2R6NvVfEsN3Hd55DPDvrvTRsb9cgl3OP0L8kIAEJSGDHEFCw2DGnyopKQAIS2P0E0nHmIPFyqBF3W52T8yS9vhAQRsF+ZwrJIpm+P9v9GyTmvhjBPhwUwkG9G+kEYci6bMPMQKio0Ej9kL2tTi0Gx/KI4DvGIwyodOZqlC6GRWLDY6BkHssXG+rEKOcaKV0hSMrYeL6QTJdyAQ2Fled2XC+8haGRs+LlVyeVTjOhZB5KwQByvOfK+Si3fVjTma08FXzS8T8Va+uW4S5caz/mq7iUs7kHlumFBoxFXEtl8J03q8W2sB8MIe2TCHO9sUgZ44dCWxsJus3IW/dT5XiAbI2M577kfkT4YJtc99zTiX3ejFr8jcBYBuIS3+p+7kKgnE1eynPgDfE4uLMfxVv3BoY4toGQwTrNKNbvq8Ii4TFxa8Iu4SnQ26AzGHmycmhz4wzPNpY7nL8zRDeHVAlne8sVyZe70OWMNu4eBS0hc28ST9igcO6sXISP5zeM2t3A3Ocz/vVHeZUfFd4r9V+NuJDS17PZELtHVkb3rnIMZ7082rWwtlXHrePOSezCUzF6eh5u8YpgSHMXQowJj5Bsl3NYYaQqJB/PKM4VO4XrF6VwHbQ8Iow6zk9cN5x7nuOcqxIpWI7zOQz3xTyeeQhL5d2CEbaEKdYvoyHf6zlLRbmm8HzY8tYoD4j+Oq6QfiWilTiVcdMtTE6XOr1/4nPsg7NJHduLua9/hey6YiG/35YfNw4Bniv/aFCdf57v9/fX8+gy2l7X5Ih674t5hAtuRK6zGMNnj+XG/nQeZniNJSxREmIvF6n3+JYu1FPzFsi92UzxfO8ExsVifwSBtcxbzXKsl9m5/FEGKoTUc55dw3ERHFL/PMRQz/8k+55Mkishz/YWpqrdODwjWli5zG9hLc8sDjx7ZrQf436SfEcoION1VntqftszD55+0x+9+sCf/d6+1Y+fjmdTPBdG/2G2Pn9pDP3HIlYk3FJ0jQgPeRT1Az+W+Xv8ufFy9dTda+/4srsOfB2DVdr0+c0P/O5sceq9yUfBwUegyP5JRl1h7cYRTxNCK9vtEmW312B/v58VLeISUc/+fsMcNs/R7rnAMyMM+6dobSMhmOIZwnP4wHRt5WAEjKNJ5n335pl5cm2Mnsxi8WjMsUzaeaw2X3uj/PgHmqdF/6Aut5bn97yo4y4BI54WJaCe7yU0FDiuyfXpRiQgAQlI4PoRULC4fqzdkwQkIAEJPD8BRnCRMJeODYaaihHcYthGVMAwv06+igttKr/NstzvDn7/a/n+f6T8wfPsng4ZI+aOp9yX8qvs6/mrfN4luhF554ZkYh7GrBptXXkr+LsS1DJSlw4WhjCS01IQLpgY3QwTQh2wnTKWUe8KF3WF1b3gMWz/YbuIwXmoedQDQwEGLgyqnCs68AgVjJJkpPEwfwXntAzAlTi4kvoOjXkYDOlgN9Gn/7yWx+m2djYB7qsSFGpk+2QQgm3r6DDSJDxGRp+OEc4woAxzRrAc1/PTfage/mY7GGPK0Mw1XaJmjRbN6NglAkElBeV3Rtm/LqYdxAWMzCVYlKjCtUxdS6jkGKhPGaLvSlLVw0086EOI85G45L2AkNV7o/LWMhxbC820OBt2qT/y2ZIQP4mGPhrfzPJEVWnGs+E0MOKf18KTmYQH2T6dFYV6VeMsbW7X/q/eKjbYx4UvubKgnbWksWwd5zkCxQW05Jj7zi+gXGD/2Waen+MSJ54jdEV8OBZ+x5oIBIMy5PXH1wz845XXd1rO2WOezyN2LBYIHIhZGDTrOuI8M3K6nnfl7cJyLb9Efz3gicbznr8reSzb4DnKu6me+xgnuQfKy4fcJ7NetGA+1y2FyjXPmBRq+yxx6HmmtmM756T04b269Xgv8i4e3msXPoX+smMI9N4ViG1fN6g072quwxd0inDBJdmEsYgXXMeEqWIQSe+FOj6QG4/rk+cqJfca87aEaNoX+/LAo610JMsebEm6mVrUunbFn33gbIWMKrt3u9G7ifueZ2ayYjeTfXfTY82nXngZcA/TbmG73JudRykiyWiZB8F8o+XbyG26vjy0/6GTr1n/5eV3/NE33/5vPnto/Mzi4PjkkflidlceDHfzPMqWk2NmdCKF4+Pdwjvr0Vcc/LZbX7L/a//bsydmeeb07NF/lGf6p1NXnvG8U3i414AP1r8j1cc7BA+Um9o2YZRXAcffCxUk7WgKRQm99axtCDoO7SHRMOHCkbwbmxvdUyOpiEbTfSsH1w6sHEwoq7tm64vEuhp9Os/NnK/l54MubJZ5hjUB41SjFC293/Ks9wgZhsc7e4jP822Qj0Jx4pKpuaAEJCCBnUFAwWJnnCdrKQEJSGCvEKhRYRhnGElHoZN6ezrWdAYZQfxYvmPE2biIcMHI1P8z5W/24P7HrPNNWf5iCUMxIP7XKff16xCT/Hwjts57LraFfyqjUI3cxkBEh7ZG89KBLg+LEh4QIwgtwPyX9QVDJ2FHalQ1HVcEAI4Dw2iLA38dJzqEdHJbWJIUzlOFGIEfxgQKx80ydJofTvlYXyqhNvWn7nSuWa6MtRjyMNrxO0m1tw5tIFpcx8N1Vzc6gRhl8YYo75x7U19EvtXmGbBtIul2LloMxSQS5jrDmFOeDlzbGGW5ntke1zCGscphwAZrpD33XoVqQmAlPBHXcuWY4JN6IEZyTWM4q3t1aMWvEEFV0ybKpUxnm32uB36p26Ct+RybDPch8cS3PAyec+BttT6vxHl/HMyse+48IYKeb9X6veWc6IKvb3lfNJHkebYZz49mCNvycMihLiqp7qXu/JzleoPj+bltLdk9uy9s62qeJxGLukWIK9OslhVqqtvOeCAAbW2qfeEZXmrO8Ewyvy7SLbNo5pWXGfOOp2A45t2AwRKhgncE4afwwiAsIMtz3XK9sg4XDgIHib55rjKP9w7vEa7fEtqoMCEGeTb/+c4j5Nypf6exD0KNsU+e36x/7rFvX9G/dwSB3qv0Dansrw0q/O/y/d/25/mGOQ5CRaUyhIviuk2eiuZRUc9onuE16IHnOtcn13MNGmlh/9rfq2v7kvsif/GAbWLD8Fp+nvbeQMDgmVECbjy9mscFdWiPhwgWy+yrCaHZb6trCs+3dXKGb744ssAbjp9+1dF/8Zm/9/DBycnZPWsPnXzToXc/ftP08x+8be1z9TChbtXW2nj1oe+eJwxUEnPH+66fFsvZX5uOD71nMV7nXud9VmG8uE85bt5VbCfJwtszA/HxjtSPZdlPeU6sxQuie4eEdCJSRdmJqjEGFrPi+zF4gNf3swJyMnafniU/eQ43Gw+Nlena5CWTlZU7I2xsRsRAHE24qvHxbI42/TSP1c5juAthxflsAkpyXLDL9vB8vjwXxcFPCUhAAhLYnQQULHbnefWoJCABCexIAr0A8al0pOlEYSgkXjEeBiRBpTPJdzpdGATJV/HJrMNItnOmzNvIb/9NZpZgwejBL0v57YuAYdvfMfj9kXxvBiVCIvThqtrP/I0Bfdu2avRpxafnbwqd6a6T2BmY+F6hkCpOeuV4wFhK3oqv55BlKgAAIABJREFUSsFIhFcFxia2gcETwyciDuvRQX+Okekixzf86XzWuQt11ocGVr7XKHAMv4zERFygY069EDAqmS3CBbHf6ZxiGGP+MM58jRqs0cFlSGsxjodiRf5uI4CdJHABAlyTXDeMZueZEcHiuZf4IraXiBZ357e/mGV4vnDNcd2W+Mc1ipjBfc/9mtGoGZXbXbdc5/xeeQrYAdfuq7MMxme2x7JNiIwB+GhCDHXeDG0a3kb8OUxM3S/SX+JdiPSzYYkuZkvv1zydY6LOB7KXFuyki/nRDQIuMaPLSdDZzjFODQP/IDAk/BE7rgTf+wi7xPbbNpoZqjuGLgl2HtHUt8Iwtb8z6nYjtrrl4vHlfIHgezRr8KzCoP7yldW15hEQI1a3fiby5ZbXR1gdzywY35r1ygh/93R1bQ0x42z9uzpdyOOkyQ+NO+FROk+a7DPnBTL5tdWbr4MwUr3I0g2Q7sSJc0Jkjdqoac492+EZf+607Xo76xFC6Jge+2CN7vSco0T1v44P1DlL8mvEMN4B7LuuP95/b01BxODdUCGjuP4wAAKW6xJ+GC95Tt+TwvuNHXJ+mY+o/9pw+ZJcb6tnr9OuGt0A9Pb6w1uI9fGSW+8FwssOkzg4dL/eOAS4Xv7Otur8L/310WZf73BQz4em97poD9VevOBarPwvXPclVNBW6jwsCNG0TEgm2o6zzTzrkx9iGa+H0TIhjiZdmKRlwiWNx2ftItu9sba3P4b3e/+oJVN9L0EeSKCkzvOVl05XB1TPPPDyONq3b38etvfE2+/2ExtHpycmx858ZuPu6Xue/WqWneUYm1odw30JKouvvuVfM4t2L+3Ymj6T6Hd/+M2v+Y5nsmyJlTwn+F5c2AZJtwnn13mANGEF0SfPs4gGi/HKTcuVtbWNzZWVM/ODB04vDx0l0t9KVJ21lY2NiBZN+MTRdd/kzOmU9ZXlbD50yqpnJvnQwYEjS55j5LtYifSxtpjg1ZHk3Ms8s5ajl0SIzvrjef5+JkvyLGrCe//ZxCkKCbojWlxYTX6+C8bfJSABCUhgRxNQsNjRp8/KS0ACEti1BOisMLKUEaUYEzGyMIqZv+m0vSwFY87NERJ+JZ8kZDyTzvWwY4PB5v9O+bae0jdk2d87Xy6LzKejhDENkeLelHLpf45hphcrCvxwdF43Uq3rJJdYwTzqj/HzvhQEC0Zdsz+OCWMTBiUMSPyNceptKV+ZglcFBlC2RYcRY1mN8sZQhbHhSqfiVCN/2c7FFAGWY99VDz45P+9LwcCICMP5wWDMhEDxnhQSttIZhQvHjXGgtkHnGeMbpcKVNKNgOrLncFesuNLTvGfWw9hRBuULGlPnsbvE+H1PDPMYYLknua655xIPvRmsuDYf7q/Te5MKYv/KdNpsTskBwbIY4bmeK2k1827NNjtjehMh2Gpn7J1txEZ2OULb4Ol1idc892wZeaj7IQz7sQXFFrbM82+5kqrwPOI32vzch3kmxV9gsZxnd2fdAlAOuucRhXWOxZDNc4ZjYrkyKPGV7+UJwP5RARhajKGN9fECo/C8Yx7P7WW4v7z/rNwNPB9LjMWg+N4UPAg4J7Cmvm+M4f52hCPCc3X1b5ipA3/XvDqWyrHAfitp+UrOIXXhuOqZXexYHr1nHpGFY6pnN3XcH4Erz6bm9VEGwDyTUVsubkPbGnlcOUAAOZguxYEl28DQua9yigyEjC/OpmqEeZeUN8ySmuRAQom1a25jnQgsSxg2D8UcIAxhwnHxvuEZ/drpdO0lubabcHTuNbclZ3GgXBucnxaeJ6KFBsRt53On/Zk2D9c9gyO+dVD3n8v3h7e1o27YQ+vFC67pzYgXXJ8VjrIGRtCu6ATn8bi7T+azPNOS0yJ6Z24UfqN9Rtvk1iZYdEp31xbafpMOn+XD7y3E3kCQHsdav7Ka51reKQxsWS4QUea5KXP/RCyZ5paeL/IOmYf/mOckbSmeo+0Zk2NBtMBQX4b7DJj51zwT/3bKIBzU6K/nb+5jPBHafRoD/8DV6xyPK5hw/3bP3PFobbFcmc1HK8dOzw7efGrz8E0nZjcdODm/6c7ZcvWuyNfzlfHszHQ2PzMdb5wuT4uj06cem4wXT0wmc3i3JycfvT6+pWGDZP0Uec+758rKatSclcnNEZlvnm0s7s088lowMulJ3lH9s30zT53EL6y8He3dsZljmuX4hsfVdu0kAQlIQAK7n4CCxe4/xx6hBCQggZ1MoHIZYHjCC4FRpBjFSUSNIEGIqG9PwSPhd9IJ/+N8PouHRQoeGP8wf399CoabSlBbCUSHXDBe/qsUxAqm/4d1hqML63vvWVEj2Fi24vDyTq3QBNVhphNKfRFZMP5hVKXjjMcInWnqUh4KjAz/ihTECgx7ZVirDjTHi6jBdq7Us2J4zG0gcsqluC6wTIUDKeNwnRsMlDUinWNlm5yr4ykYy7oRfV1nmePn7wqVVRw5LrbBth29OzxLfr8UAlxHXFsfSOGZ8JdiuD8ameE565JEub8G39L/WAbvGgf/+v6eWJnPNvp8EJ1NJgUREbGiwu+0TczY5vYRt5dS68tdpnk6bNmImmG6hVEakbR1gvdIRraujtZPP8t99IcpPCd4XuDthBdIvLbGGOzwhEIYQEgoHvzNvcy6GPdLXC3DP8vClonnKd5V3KuMwM+zYcn6GN54LpRxqfI2cP+z7IdS2N4fpHwshflvT7kvhTohcOKVxbJlIP/FfJ/mucszlGckx1M5IHheI17zXqhE1Z0A1T1vqCf1wrjPMtS/wnTxN+eTZzHbYzmOiecyvxF28HWr+w68Fptc9IwDEaWaSLwVIoo/mhfL4Jy0eddm2vL0GEaO6p7W1AO2/IXBlWnahLXmWdIqxLy6XmukNuvAhmsYlmubmxdO08SA8dwAH85yv53Ce8tn87U5tS/oVvpQUHiW4U3B/VDTD+cL7YwdN5V4gbE/la82WYkY/M18bo48J8YIl9zzHDvPFYRK7qPcVyiMeAaQeqJ5aaVcahOpsGUTeXf03lxxOZj0IayWT+T7rWgB2Q1txT/fPC+65w5tXIREnmOEvtoKDfc9d2Wh5ej1cYobihU/leX+ZHtY1PJG6D0uqHyF2eQ9V56IpyNKHHp0/SW3LJaT+TPzm6ZPzW67/VOb971lsZzedWTyxGRtGneLuKOkns+ujjfPRLDYjICxnnQ3iwMrp57dNzrdCRZM7GXYWh1cPSWC4liymDWPtrZ0MiodWJmO44k4unW+ubx9trnk+fJMlq92LsfPO4FyKseznmNrgqmTBCQgAQnsHQIKFnvnXHukEpCABHYMgfOEIaBT97l0tOnUYeTCII7IgNEFQxydGmIxf00KSbfpzGH4eiDlu/plfj+fz+l59t4Vfz6/vTEF48z/lfJLKWc7ZD259LXK8FOjc8urogxIlZS3C0XQGZboKFL/MtBhKMBoxHFgUEKc4HeM/YycxQDH+kx07viN/bE99lef/SJX9VGjiS+2kWJGRxKjJZ1GOr4YATkGOpYVMgfmnCM+MVxWO4PfOZYKqYOVrIxfNYqwfV7iyPKrOmhX3nUEasQ9xh4MH6vxjoi5JXlO+7A/NTq9P/JEO1rpjc99aKbO6sw/uW7H0wgAMZKfG5qpC3GR0rlRtE11xuwufFMfRYQYR13eimbx7UIMtf1HUKhQSKzb1Yl5XezwYd6Ns/XtQjH1ybQ3s1fuvxY2KOucysj4Pg/BnMDn2eMcwxuVw/up8g1w3/KciVF+icDwcAriAEIhRrtj/VDYMuqxPPdwF4O9e95SWJb7lHv8kRSOE44IFuHeQnvw7Kok0nWPM+8z2QeJbzl0wgshbrAc54xnIs8GBBPqVEZHlm0Gtxwric2P5ztiAhPPF46dedSLdwAb/2z2QzLe8hgpi/yJzH8089keQgYTosyX9OtxPDBjgiHbf3RzY/2RiBUVdonnXZ7Py7x3xrelPgmTstzMqdvEA4QQYHV+Ky9GhSYbXn91zWy5KfTnvrsGKtF6q0fq3pbqvfbyvcYzt8TCOdxoVizQcmy0a639VddUCc14iqzkp35ceIaAj8cZ1TwMidU95rv9TxLHhXD/+3MPEXS/8SIclIJFf4Hs8A/ex3hyfsPgOL403//sInnBdsQhbwsZ1bwO+op3ImrXwOB+qrZVd02Px8Tv4z7HeyrJqReH4o6X531zSCN2XfdZN227Xfqm0XO86LhPBwvGnyLbjxgxzjN0eSx76GLixespG7kv86hj2rFjnoVPZv7nu+Xbs3B583REEu6fqBOQLf/sxmL0P+ybtOfweaeBcFGqS3nFrd//1JeOP77+8ptPLY7ckf28LhV5acJC3X5iduut47Xp4XlejYdXnonbw6l90SgOzRcrm9PJ/OTaZP3x2WJ1PFtMk9JiPMdJJW/M/sGxJVK3cHkdkrPN7f65tAWlybysPBmvJBzdLTkteae1QQfrwbyeVU/l73rvwIWwVzyT8bbYenTuiIvSSkpAAhKQwBUTULC4YnSuKAEJSEAC15tA35luo64iNGDwwp2e/BT/WcpXpyAAIGRghKKD91spv5mC4Y2OacVnH1YdYxfhjJgQOFiHsAiEVem6Xc0u1cSKSuJYyR7p+FcybfZRIQhYjWUYDUxnlI4lRkJG/74qhXjiGMtYvoyAbB/xhe3VxP5r7Npw24NFnvN12Jmr4YHbhZqhUHEpwwcrrAvHgDGTOtEB5pjZB4ZRjId4jJBThBHdzMfwx/GXaAP/rdAi+b4lVmwPA3WxA/Q3CQwJEKImCYa5lrjmMGp8PGFuMMhyz0wRCs5G8Gm3RwbLz4fh3GpzjK7FOMK6XLPYpLfuj27EezO9nHNf1SLdZxuWyzMqhvWEBGnbaFGMiCo0WzbL11Zt+F4iQT1bqMvQmFb7q+cI9+KLsjWWxysATwpC4iG2xitk8yXZIc8UjMzcq5XMFI8BCsIozzmSKPOMQiy4N7Xk2Ykhj/sTQxE8axQ/93VvzGv1hTH3PHXhM/MSJ747Fkbvc1z8Xb+zzEd6az5cYVweW3jF4HmBsWr4XK1E5cAjTByCaeXBqdB7HB/vgC55a1f/j2c/laiWfXC8PIdRhjiOEjnYHqOr+Zvt8QlDnlH1TP90BKF356yyTdZlW1+eY8UL7o19GJMW1i7fb4tAxvOwris+h544nMdy+aF+FboqX9tyrQwut3pflYGV5fqpCROdVbTLa96u0aHY0Y9k5vhbrou+rk38YvHennqOVZVtkNsE5SzX0cb68iQsEAD1fBvQ3wVf7+mu4/aMoL30MynH0+bZVSPYI17M46mw6EUMcl60Z0l//rj/miDQ33unmmjBM2SxSFLscJnPjiSWEQI1N0xTB7upf/yf41XX7p7+98GizCFe4DKi52TyWLJRvzyfq1EEkTES8m15ODddRIyUzU0yVic5doSNLpzbky8/MN782mPjv5UtRijtpic2Rz/7Nz+0eOIz66OV/vguKCT2xv35O37jXyw/dPqL9p+cHzlyZnbgvuz/jZPJ8i3xx/tzq6MzR6fj2TNJtH0iqmaE+psOJ0XF8mBQ7ZsQOTADSUbjPJ/XH09T+ImEhMqzsOUEmaZeU56sefrGG4Pc3O3ZOanAWltE+pZ0HcM86ZJwQumQjVeS8+LwymR8mKfgrEVfRKQeRaRua9Szkh8qgXptyk8JSEACEtjFBBQsdvHJ9dAkIAEJ7GYCvXjxVISLn89xYoAr0QKj0Rel/O8pf5rCSLX/mPJv+u9bWLIuBrn/MuU7U+iAER6EDlcJFGUIKqNQeThgiMcwhwGL75VYu0KfYLTHUMR7tgxXGNMwkDHS+c+lMNKZqbbN58Xey5ciLNSx0bHD+EBHtsJTbR33ZX5hW5W89aP5TtitCqfSj65uo6UJa4BRj31ifMMAWQa6MoSUEbMMYBrCLvNkuPj5CTD6O6IF19MjKf804ZwIBfe1ESvuS5z+lvwaY3DssFyfGNwrP8xwg9xjCImYUjCO51nSXC+275TrmPt6KC4mHNOEfBcl5jWDTvIKrBKqCftvXzdEBowu3CN8J2waAgFiJfvmfmVZnh8YrfoYP21/3E/sE8+y8jRDsGA7NZVwUInumc+++BsDP/dshU+qXD18ImYwcdwIrOyrz0/R6sN24VPCUP1WAsxQMGI57nnA8Xvd58xnvVkvMvUhWtp+y+hWxvsK68Lf1IXfERnKy604l8GxjrOJVP2+y3ON53TFcEdM4vipH88r8maU0MVxMr/CkjCfZzb1ZH+wgTe/88zjeCrsFNuv42A9RBJEoPIIYd3j/b4wGFMqdw/LJQfFyp2IW33YssrzsZZrGMV8MGp7az+ckxJ2+t1TqyY68Bv1RpBqo57PM7W8SPGmOICoxz4IMRaxj7r+Se6ZX87nu1KGIvMFNuXsnUCgb/Pgyclz5P9NQbgk7FqFh9sJh3HJdSyxol+hRMNqozC7xOezAuJ4XM+I25tosVzwrD04mq7Fnyn3FulsSOPTJaXf8lu6aKXGyc2wXJ7MC+JUbrAD2QZhoXg2HGhiSEsp1O7TtCfJrbF8cSr05LfcMT58bLXlrmhTXOw+/jOfWR6PWFHeb7M+f0fzINl2vFtV+veff2fEgOWX5dnwl7L9Y+PJ2ism08mbZ4v1Qxubzz4TwSJqzvyxKA0nZ8uVQ8vJ0TPj6SZeFXlXLePMMT+RZNsPHJs+/omjK089mzcd9e3r3ySLYXuPdvWFnjk9s3OxgXLG8yefnV/i6EDm0bbmOVrPc94D5OkgPJTeXpd8F7igBCQggZ1LQMFi5547ay4BCUhAAiHQCxf/MR3xj+RPjE9/NYXRg3gxEI+e0btvTUGM+N0s9xtZ54l8YoAiLALLs+7xlHetrow/+IYXH6YzVuGe6l1Z8+jol2BBp5HvFSscoxXGLAxBGP0wOiJssBzGSDw58LBg+UvNQ3E5QgXXBPWsvBLst+bRwSsj4KVusxKCVzgojouOKAbWSoiO8Q9jKCFk6vcyulYc5hp13I/G7jwr8Fzp6+eHBK4FAa4vDMh/FOFgGSPsM/FqeHPEgsN9uKXy9sEDgSTFBwl90w1WbwPLxzEWc62yDa7p12Qbt0yTeLvdRF34p3GSd1dIEWZzLbf7KfvkvmBdBEvCLx3JUPXXZ7M8MxAEfrf/jfUJB8I9czyFewnDOM8K9s82MZqxrTL8135YF0MR9xjCx8MpGHKawS1Ti4Gewr3L/DLwl6dGeR+UoMl+2D/3NeuVWFNCyfJ8oYAiDm0bbrxl+GsjmHtBgk/+rKmN1q0/+uTN20d18/tmtl+LbT2r+m1uDdq9QL3KE6TW52+EgTKgVUg7focfv1e9ikHVMWFJCOPSmJQ3WIWagnuJX5WDh23Wsw5DG6J0XSsY9PA84/fKF8KxsH3q96ZcP1+eUDTUgeXw9mAbL8o11+UUSdiUXIQlnrAuMahWuYZbuDEGOseYGrFunmv1Y6k7QsPrIkKsRgzJVwKxtATiCGgcM+f9sVzPpwhaA6P5KHl4c01m/fdlY7+f7R7P3+Wlw/E57WwCtFd4PiFS8PzhOXdmpyTavhr0GPNj3C/xtMLOcQ8zrwRYYqJ1Am1C7uXRcDSfhzLvcG6sg2m1kEibZ+9qBIyuOi1UFGXQnBmGieq+8wzJNhdRBlknybfjlZVyLHfevsxjn308tlXUw9W15fq+o9Mt79+2q199fPm//eJjzXOPZ0vVnfu4rU/ui3acv3CC58xa9pd3yvil+Xxdln579vWVo/37Dy6nq8cWK5Mjy1Ozp+aLtUfnk+mJ6Xjz8ZXl5uN5wT0Rl4pNclgcWTmxSP6Kw2vj9Y1bVx/9ZAQLcllwQE086LV83kc8gJg6EJ3nRO+Q2H0/F8m5TdDyWyzPjPYw695xPBs5VyXMNvEiokUTnxQuGnMnCUhAAruWwKUaLHYtAA9MAhKQgAR2D4FehMDw97UpfznlZX2Hh1GxdNK/KwUh4Qf7v78tnz+Q8v/lhfi+uKTf/+o7Dv7J2pRxXq0DS8eQDhPvyxotzN8YFukw0qHC+InXRCWcxgCGx8fHUhgli3ByXwqj9Eiq/VUpjKauEbn5ek0n6o7BizpXHcvjosLO1KhCdjz8zt8YpzB08YmQg0ENcQXRAk8LCt4U8GQ+f3PMZdSrUYwVMmbLoJtlWvgbwz9d0/PtxgYEYujmGi/vJwy9JE0mRnaFA0EoeGXKq1MQDlsIiz6mOMYWYo3fn3kPpsTavozI2EIscT+V8R8jf41gZ37LK5P9fLjPs8A9gycS23575h/LfLbHiHXWrdw1NTqf5wTPmxIrOAbuGzwAKmwUBqJ6DrHvEiAqsEYZyssgv+gFgfNeHwPBoYkLe+kiOt+xDwSSJrL0y5RHSJ9DYkvYqJBOnKMKC1hCAstyLiqEXwkyZeSrUIH39dcQIa04hySB/08JPZhrhfcH1w/idgnc5Gji3VbXHaeMfZd4xXMVz8AS7d6d33iG875J2t7x/i5MFEl+W44VrsNHUrguqUN757F+lkWM4f3Fc/2J8GBZp11AIG0knmW0RSq59qm9IFac79TFuM89WaUEzbqnGexRrHiOH2ziQuIltXtuMkk+nhUEQ1RCXJo6m0q7xQafFSYKkWM8vi+//+Xkxrgp6jbr8dz9o6zEvUpC7uYlwbS2MpkcGs9XfvqNK99962obbDM6fmb0rn/wkflPfvxMxOjx+GQvkJBACW8vzifPmi7M1TKhplrbc5lBO+MvyTJvy1yeJXeMjhylLnkCPLueevxBKvLRhIc6HcHik2vjMx+6Y/VTH4wXxeiVBz+0+upDf5owUkePxqNiesvq59bjicG7tcTyMGnCO+/ZBHJqz54k0h4n1FXeZ895q1Cts6an56T+6LH1ys8yv+e5M0aMoc1Om5b36jApfAsrqGhRV42fEpCABHYfAQWL3XdOPSIJSEACe55AOuUYjb4x5S+m3JfCqGNGtRL6CWMhcdNZ5jUpvAt/bjoZ/8ith1cfefHRfXSCmDBCUliOUYkYqTAAVVgoOm2IFHTWECXo3DKPTieGSDpYGBzp4CFoYCTF04NOI8uVgbHf3TX7oMNdRrLyDulGw5VxtjN21v63CxawoQNNYlyOl2Pn+Oi0lxGVhL2MziwDKqP76ChTML6WUa1GJXNwJfikI2rz45qdbTf0HAIxNnPPcu9itCF+f5KWxojS3Xfcswh5GH/ruiWOex96oiXdxmCLMZc8FFl2zD3MvcSzAwMN9zaCHesTcodtrWY/J7If7hnmY/DF0Hsk8+/oczAQfqXyMPC8wPhS+RzqOMpoVcJfhVwamn/K62J4I239vtcEiC/kLTAQLrY/J9kt8yqEVfEvUYv5FcqEeeW9wTyMoVwzrMM1wHm8N+V1/TWEkY5nNvO43liXa7beQW1UfArXJaGl2D4ePFx3PH8x8LENntl4GbIv9sFvvJtqXf7GEwdDYAvXl/2f7r10qBe/m2w7EHbL1IeEQkw7GaGiQjbulsO74uPoxQvWr7YR91q9M7r3SSdWdILFeMw9xTMcj4sDyQmxOloN1hbbKHb7OWl92Fz/iMZSPx7znnlHSnJkJM9OVolg8FCW/eMs9uBoPN2IEJKwSLPxKw8sj/yVO8av/6bbCeGUG3Rz9Mmf/OTyl371c/MH45p6Jutj/W/h9fIdwZF7nvuVNljcBpfxqli+I+VtTShZ3Xdn9hcPrflK9kEqpWdH62d4x/1sfv9DcvRElNjYNzn99Jce+a3P3bn2qcWrIlgcmZ7YP1uu8h6cRKzgXcRxc/3wPcfenk/kZovLVlMjbtt3cIp4P9o8k5QWSdVBiKd5sjcto8+06FdoOlnyQoJFn38HFCzJO5TjOw6GdrxncwNxvKcjWPDcc5KABCQggV1IQIvBLjypHpIEJCABCYxG6ZhjnGR0KV4NfCccE4IBnUw6PhjhMV4+niGt/2zfdPzrdx/b//ihtcTXOCs8gJLRiBg+6bTWKFo6bC1cR18wHLFdCh06jD0IJOwH4xRGJYSKl/brnc/4dbmnrQxkiALVycZwtd17ooSC8nQoQyiGUjqDjIrjWPidkXoYVSkYbTF4VSJzuLAso24xjtFBZqID2YU7OBv7fWgIqfq1EeGKFZd7ml3+SgjE0My9UCPhuf8rpAT3M/cp934JFoycPRoLCtd7JbfGsMs124X/6K7vyt1Sxlyqxvaah0W/vQqlhFhZSV3ZXwmZ7LM8uLhvKENRou4Xtk04pis5fNd5AQlsC2dVI7hLIK5Qg+WJUaIH1yPvDp7JXCP8znXDJ9cE7xzW5dnKdcVnefhx/XyWROy9JxHrM49rE2PiQVK+d6JZ8yBiXZ75lSuF67nyd1QsetafK369gBfSF2DXaRe1vv9e9aq4FKQRL1hs6FFX75Lyusi9urw5b4dOsGghkCYIEISPitfBfP9odX/M7YgXudUqZNQoYaVGo/8k5bWx4t82oqk5nz0a8eAD2Vu8gCN2x4p/++ryyD955fidrzs0fiMVyQNi+UOfmP7L3/zc5qdOL5brWWbeLP/jMV4MCcu0QMB8Ktugnng98KzoxJGV6etTtyQPT0w4QlghpMw2PpkcHA+MFhFKlgkNtjLNAJRstzvmxQ+/4rs3+hhM/J1KLnm/9TajceVsQyzh+UPbFw+QzQgSPMtuXlmb3JyF90ekQMFIYoqWhHstoe3S1I4zY99K7RxMWhzDrdPSUHWuGXhYxA2lhTj8WPZOmxMRtt7pLIP4z/PyVJ9cfGs7fpGABCQggd1BQMFid5xHj0ICEpCABM5DIJ1zOjcIFV+dgnDBKFUSXtPRap2wvAgfTk7TX9g/nfxa/rjr2MHVzx87OD2TnhUdJYyJ5TlRI2cxIGFcYvQrIgRiBB1EOqMYnPgb4yZiBaIF+8HojydGGZ1KbLia93AJEOU9Qb26QOVnp+GobObSKaXQySO3Bx1d1qfTSZ1Jqv2JFEZIxW47AAAgAElEQVTd0metUYRsk3Uq/FOxYZutw5iCgatGlzN/6MGBsWxQLb9K4PoR6EfJV8gP7pMa4c5zoO4j7lPuT/7meq4wOPzNSE6u/fJSqmUrVFqJEEMxguu/Lvra9zAXAtut8EPbcz1cPzju6boTQNDow06x73pmlzBWMfabwNs/V7lWarQ31xXvJD7reVsiA/MxKFa4QT4RJsrzj+t6GKIKoQLrLM/+EsouGkrsusNyhxK4AQhExCihkXcH7SXuMwRB7q1n+/BML2p5KcYJIThZId9MnBZic0/sKIz2+cy7ZxkBcZzk15PX4EIQ4eCZCA7kq/m1LP9Y2qLLeFa84e/eO/m+Ouz3nli+5x8fX/zWZzfGZxaTFfJc4JnBZhPNqWndp/r90y59SRPfJxPKF0U4uTVPkUXcHWjtLvIbYaB+M+Gofne0Mnlf1r0/OgLvuvnGf87qz51+/P3vyA6zr/asmnAMTfwnR3a2eSg/0L7dbOJJBIUIDggYaTs2YYV8Fnl24ZGyPJDjW2mpLRAmome0n3M8XW4dFi1dhHosn43MysCYT0TkwKOR5xfMORfsi+cXAwNORrDYCqd1A1wuVkECEpCABK4RAZNuXyOQbkYCEpCABG4sAsQCT43mxz9/+qNPn5lP8/ebY/2hs/me9I3S+xo/MUliwQgTD+Tzc8lfcSwDxF40X2SE3GiMgRJxg04RRkzel3SWMPAzj+1g5CEXxRenMDKbThzL1Uhu5lW839oGvbEyRF0rC36FgGLfQyNpnZDaD/tlGepNJ68SbmIwI455HRfCC4ZVOrEcAxPiC8deiXyHo8IrDBTrt1A1vThhB7LOgJ8vKIFhcucYi7kuEekw9tbo9/JQqsSrlTei6s09VtdzCYRc90xc80MvIuaVl8X24z6vx4ReFC/o5XHdd17nu/9s11V/XXaJd89O7XsvbvDcpnDNcu2VNx3LNPGrv6Z5d9Uzn2Uq0ff28Hx17c6yfZ/V1/0qcIc7jAD3D8/+8kbi/UE7kPZeeUk9Fst7l2NhuaD9hFhIG/FFCfd0OGGZZqPZmXhULJ5qXhfzlJXpodFsgectQsfTh1dG81tWY+jvpw+eXP7pz352+d7PbowSYAnpoV4tJO2elXDeiRTj5vHL/mh3Hk6ujISxWmzGy+OZrEeYqOTJGP9pNvOr+bw/esFn8jmLGDBNdSZr//ap+cZ8ZTH6drSY4XRm+QNv+fftOZNk1z0HwlFFfDjrXcsKJbYyoAUup1Mn2r4IGhzji6JJRMhpAwDWxpPx2nJ+7pgatogHRu+U0jw+UmDNRMXKWxG+52vvbqu7f0pAAhKQwE4mcK2MJTuZgXWXgAQkIIFdRIBRWzmcKhxZGxn32afXD544PbsrAsXywNrKWrwoTsarYj1e6ZsRKlYjVLwofac7M+/A6kpz3aczWKPpMNAz0guPCTpieEvgYUHIKdz2awT1dpJ04Ia/VSLq8oYoL4QrOQNDDwv2U3kxypDFNs/3nscoxmi1d6WQVLvye1A3jrcMYoy8RbDgbwQORpjzidGsJc/uP+uYWtLXKzkQ15HA9SYwyE1QIuLwfjlnlPm2ZYeGYkLmXO+quz8JVFLw8vor0QJBbOsZfJFrvISQEjokKgEJXCKBPmQUbSOM8RXarXJedHlrlsvkmSDvRfNSvXs0md7WEnUvIjIsl38hzaqvbJ4Kq/sybGb9dESM356uTB54+7GV0ffftfyGu/e3/Gqj/+6h5U/86bPLJx9bbyGbmGjn7Y/QcFOs+ngx3BoLP98x5if00zTJwCf5nf9oj40/mzBQH0nBC4RBKsmXMf6jlEfyN4m78ZJIUossm5pk+Vl8HXoB/pnRmW/FYfjc6cff/01EekrJUJ8mWmT9eFv0TrSLxaLVcYV05Cm0o8vz+M4sB7cIFstjaS8eW1kbryxmC3SYZfJdxOMixMZLvDVSluupHu3uD2c7tDu75OedcIRgQdtVD4tLvG5dTAISkMBOJKBgsRPPmnWWgAQkIIHzEohYUQlQ6/3GJ50nOpYYaXq39jZKq7wmmE9nj1jfjEwrN388LJh3XwojWjHg01GiA1a/IVqwzqVOjBSj44Uw0Dp1l7rieZYrw9T5RIIywtbI8PKuYDMcC/H5Sa79QMrx/tiq88fxMTFSsEKFlJEWcYIOYokU8GgjdxUrruJMuqoEJCABCUhAAjuCQJ+ku/KdUWfachWuiO8Y12kn0Ra7LcZ3BrlQaC9+eRMsVpLHYjKdJqcEYZqO33Nw5aF/9qrxm+7d38KKjk7OR8/8nQ8vfuqBk8unM5iG7dAOw2uj29YYb4ok8ka8QDdYxGVjdS0yQYbhzJKGYmV6Jnk1Hoz+8Cf5+7HU4eGsl3wVGXgzTvtumfbdMvkpxoSqahOiCAm9ew/alpMiJerLt6I5XHj60fu/ZZwIV/1Aoebd3IddbRkrKqcG7d6WKDxVffHK6uQlSfVxZJZ03bONJNdAYhlNIlIs8cBodUgIKYSJj/V1Ky9i2p2VYLxyWOgldtEz5I8SkIAEdiYBQ0LtzPNmrSUgAQlIYECg96qgI7Q9j0OFaKIjSQeyYntXbHCWr/wSiBCVOBejPB0gOlq398u8PJ90FisMAJ2zCpl0qeejRuNdjWfFcF/DgQcVH784sBydOrxCKokr4sLxlD9OqZA4JGfkWAn3hJBBZ7DEnXLxp74Veorf2ddWCKhLPXiXk4AEJCABCUhAAjucAG2kCg9YA2FaSMwU2p20Exn8QduJwSAkr04Zs8z7U2g7fk3EBOavTvftf/FX3Dw/fO/+5V3F5UcfWf7OR08tJxErboq4MY0QgXbAIBpypyX807gf+IKzQ3YznU7iSXEmy9E+O5P8GJ/K9h/KcrTrmEd7FjGk2ny07zIwZZk6RVhYLmgTnoj4gTdthaej/hsJFzVLjosLetD+3bf+wjLhoqrdWGFP2T4MaPeybQbB0I5cjTixHj+OU/ON5UsX85bUm7Zqa39yNI3buLXXYVwDkdgeyzGQZnv4vMLmpwQkIAEJ7CICCha76GR6KBKQgAT2CgEEihrR34sVFQ6JjiPiRAkD1WEimyBeFBXiiA5Qxb+t0E/8VoIFHbZKhsq6dCIRNNjG0CvickMg1X6rY3c1p2zoRcJ2KgkhHTpEGEQXEmsjWMABJuSiIF8FI9ZYBjGmEg+XAMF6fC9xZysZa+bV9woJVfkqruY4XFcCEpCABCQgAQnsCAJnvnUrQXUzzsfjYujNWoM+WhLqdkBxHeiyM8TQvoy3LuGXlssID4uXj9f2rd42XRy5aYqg0U0/9enlZ9799Oie9QUG/4SDms9ZF4EC74q7su6ReFPka2bP1pcRKrLdSUJLzR9vOTKSDyPLfC7fE/5zvJ4k4PlYHk4VED6SfDvJwMdJ4L26SqioWcJSEd3pZNZ7tIsIRR2TpLsTHE7H9eH0vn/31Gz9rwxEi5/OoX/X2TEzSXzNeolh9fXLM4uD/aCgrTChlQOEz/1pv2+SZHs+WxJO6qb8vQiTp7I0Hh4cazw/WlsblsWTdRErED8QYCr59uW2w3fENWYlJSABCUigXqKSkIAEJCABCdzgBHphglrSSVnJ3xjh6aiU+3mFQapk14wmI/wRhneM8/Qw6Xx1LvqdtwQdIkI90QmqBIZ0GnEzx3WfzuF9KSQyrHWHpC43tOIwt8blrrv9DFUHsLbDsSJIEPOX4yFe8e/3x1cxzj+cvysJK5wodAYZAchnF3+5+76V3bH/XqPmqIchoLafDf+WgAQkIAEJSGDPEegFjGbpj3hRngAY1XvvgGa47+Z3YsWzyWfxhuSwmO7bt/LSWyfL6Xfc2QbbtOmR06MXPT1bEvLpiZQMImkqQvJVjCtkKd4WBIrqjPjz2ROjxSSDU5Zp3y3TDhwjOCCOJNQSKSey2CRixcpq8rNFR2EtRIzV/UcjXmRW4jJNVhAL9o9m8857IaJCPiOSjKfEasqszRwbIkw/cOXEcvTzT1XbMvkuaGIvR9/3ptYkLRFhI54XbIc2aQ3UmTHiKLrJSrwrNpN8++RkMqG9Ps/x1GAYtlGhn6hPefnClFLzqh+w5645D1gCEpDAXiBwtcaSvcDIY5SABCQggReYQC9W0GGpmMF0Avs4u1su+CUGIDTg9k5+CTpILMvINArboIPz0pS41DcRgtFaFTKpjPgMXWNfBO59ZQpJuM/nWXEl79HhaLArWb/OBnVGfGDiOD6dgvBAx5BPCp4ij6QgXuBpQaGziWcFx4+YgzgDEzikc9xCQ/F9GLaqPCtafc1XUafATwlIQAISkIAEJHCWQJ+YuzWX+kJbi3ZlH7Z0eWi0WL4uYZy+8i1HJl/3D+5ZvO1lB7o25h88PR7944eXo8c30uyarsbzYDwfzZKZuss1EemA8E/Z3OYsqaoXT0b4eDyfn8pPn8ivtN/iZZt1uuTfNNjYLEIAU0I/kWMi85jPttpQlOxrX7wiFvNnRuunaC8+md9oY7Jy365s67WcESlDL5KNiBUXzSER0WLIooVTTbv+QPaNJ8XBtCkrvGq18REw2C9t0mrHsw32XzkumlgSz44mFDlJQAISkMDuI3A1hpLdR8MjkoAEJCCBG44Ag8gyVV4GRpfRkSlX8YpnO+wMIi4gSLym7+jQEcKjgmVqdBa/3ZeCiNGSRqfQUWJZts98OniV5LBc9StGccUsrmTU1LGEiKEXxXaeta8SAy43lwXrEweYDiOfH09BXGDf5SnCMRILuMIRIGp8pC90QGFYoaBqJCB1Zj22+XQ6jyznJAEJSEACEpCABCRwFQR6AaPLzdC1RWlrHrx1unzV9949/r5vvH3y7bX5v//QZONdJ8ZryyYmtHwUq6OVJNPePINAkZIQTiurJ/L96YR3eiJhnh6N0Z9QTk+SH7uJFDV1YgUzZpnPuggV2X/L0j1otWZfa6nSfDYbzTcRBSiIEizPNvlO+/PJ/E1bkzYobUzairRBGShTXrmLCBjPERF60WJE6Kgff/87iVEFh8ozV2IOg29gwyfhSREtWi36/bOfyqE2z7YMB3X2bPtNAhKQwK4jYA6LXXdKPSAJSEACO59AL1LUgZRYQSemPCXq/UVHiU4NIgWl8leQa4LOEJ0Z/NRf1nd46OzQySJxIXkpajm2NwwtVfGIqUN5VrAeAgkTy1cdKlTSMC/FhQYEVBLri4kaFzuBdBoRKfCUwHsCYYIQUHCgPnQe6eDBhH0gvlQHj984lkpkyHJ0/Kr+bJtlaiTexerhbxKQgAQkIAEJSEACz0OgQkb1uS5aeKh4VGz+Ty9fefK+A6O31ervPrH85AeeWn9iuXLgroRoOjBa33gkQsRaPCxuy2dEiiVttuSnYH7CSo3Hp0cTwkYlf0VryfX2+4w6ads8K1503sWTSZefjDQRTbxgoRYyahnPCv6YZhnazDWYZ6V5ZODl0YkUt+Rv2p60MbtBLuPx5zOPLXUJshNKKsdZYUVbNTj+PsdFf6jEoWo5MqgPy3bCTNdeZT8IGNUerYE+lWeNuihW9CT9kIAEJLCbCShY7Oaz67FJQAIS2CEEBvkpqPHQhZ4ODH/zWTkk6MTQYUGgIA8Fn4Q3wouC7zX6CldyPAnIQ0F4KDpAGPAJGcX7rxJgM7/2UyPE2OfwHVliRXWkKiF1ER56V3whqdOZeziFZNq4/pfgQH05DupHCCjCQzEdTaHuiBMcL/VEdKkO4jBecOsE9st8IY/BbUtAAhKQgAQkIIE9RaAXLuYIFz/66snkzrXR96bxluTb3fQHTy1/7GQCQKUpFmEgngadQIErBG28myMGPJF5Cf+UtiwhotAlFot4QyRh93KByDBtibVX01xOHu78ViGhqh1N2zVhobY7QBAiqoWQ6n+IB8Z4zDbbD22dyfRIQkalDb0kVGp5VTBophsU00JNpR3aiSXVZr7AIBiampPO86Nrd1LKY6M8USo/Ri1TIaD0qthTd40HKwEJ7GUCChZ7+ex77BKQgAReQALbvCiGIZLKe6HcxctFnGVwU6cDRMcMbwoECpZDmMBr4iUpdLgY/YXbOsvgRYGYgfGe78xjG4OEiF2PLBMhkVi/EnIXofK4aKkKUyo5dYkrVf/nC7XIcrXO8y07PDt0DhEaypuCY6PTSievhRbov3PcLItwQSeSv2sUW3UOh14VNXKNfVUP1s7gkLzfJSABCUhAAhKQwDUi8Idf0pqMtF0ZUNOm+XL0yyvj0S8uSCwx20y7dwNPCAbZICSQBPvm3quC9t9d+btrpy6XGZCypJ3MYBzalQcT1ulI5q9GZEjOiwgIzQMiTTu8Ks56YZw9mt4ho+2rm/Cq6MQKNAw8Msb5Z2W6lrBRGRyz3J95DHyJqLJYzTZpm57IMrQ9aWOWQFLt0XM8d3/gLb88JLlMuKhK5j1sF9d3vSmu0XXnZiQgAQnsNAKXYyzZacdmfSUgAQlI4AYl0IsV9Q6i51beDpVHohLwsQydMoQGvjOai04SLut4TSBEVM6Jl+f7W1Iw3iNskLsBL4RbU96agpjBdumQYczHQE8nb5hMG88Etk+4KOpSdaQDViIH+6MwXc17dBhCqt9cq1sJB7Vt6kMOCjqEdAY5tgdT/qz/m/pTHwQNfkN0oUNLobPI9kokYVub6YfOe6+W2sfSRNp1CvyUgAQkIAEJSEAC157A/Z9gHElri35tyk+mMNiG6TtTfu7L34tbRBsYQ9uuklAjblRhXdq1fDJohRBNJVjg6XA0hTbsrUnOjZiA2IFQMY6HxMUOiOW6dmkX4qmbunW773ySWwMBI44cbZptoIIkl8aY9vMns8zn8z0CRBKLj8Y1eIj2cwta9XwJui9WQX+TgAQkIIG9RUAPi711vj1aCUhAAjcKgaFnwjA0Ex0wSokF9Rvz8KLAdZ55ldeCDhzGelzU6fSRbBsxA+M9Xhgsh9jwyRS8MQibRI+tQkCVZ0QJBWyH79uTYbOdqttQ4LjWPBFSEBkYbYbwwnGQs+L3++8INBwX3iKMzHssBWGCDitiBoLEcKRa5aeAd4ubnNIEkV6g0JviWp9BtycBCUhAAhKQgAQuTOBN+elXBj//dr7/Hu2zbfku+lBJJL1GJWhtY9q0TPxducdoB9P2oy14qM85cbCFhBotTyaiVDwxFvuSF2MtCbs7r4lZbWarFsMBOOcbUFPhpTrhYsGus8pkMh5Np2l3j5OVY/0laWk+ntkIFSxQdaTeLfRTwmGx43mO0/and4gEJCABCVyUgIKFF4gEJCABCVwXAgOvimGnqDpgCAkY4ksUGIoWjMzid0aMvSwF4YGOEDkqmBhpdkcK7vB4GGDUR3igp8a6dJx432HQp9QotRIlWo+uL+yX+m0Pj8S8ocfF1TJjfxwDAgWiROXlqM5d5ZnAQwSxhSTb5eVRHVPqQz3xqMDzBKGjBQbuj2UY+qlyUyz0pLjaU+f6EpCABCQgAQlI4IoIMKjme7at+aN9O29r9rnCBR4LrW3KgJnmKdv/XW3X+iQRN7/RJkwejAXtxLSVlxkAg+fF4uhoMUtuiuS86PJddCJE86JIc3JBzgq2vM15ePvfLNu8LvqxR+PJSsSQg5l3cLR5Bs+KtEfHtG/zPfttA2uY15J0r5/5lpuaWBHxorVXFS+u6DpyJQlIQAK7nsDVhLLY9XA8QAlIQAISuHYE+hBElUyvNlyeC4R8ohOHYIA4QRioCt/EiDEECcI6vTEFQQJjPJ4HLHtfCqIFYgRhk97c/12dNoz/LIdxH6+FSrpd78ASLPgsjw7qV14XJQJcS5GfbSOuPJryUAqeEtSHsFbUlWP+aP971Z/jYz7iRiUNR8yg0DlFuKCuHEN5sNQx1KeCBWfWSQISkIAEJCABCVwnAn0oKNpn35HyM4Pd/ka+/xcpbRDOW+/Bvn/hqTfyl3hBW5B2dbWdKzcbG3lRSg3uoU2Nl/KxiAprKYfjGZF5USyaYJFNLGaEgjrXi2K7UHGhajVPDmrS9IduI3HqGC3naa8uabcmROv4sfzE4Bvaq+u9KFKeFwgyTcTohZrrdFbcjQQkIAEJ3MgErqXx5UY+TusmAQlIQAI3BgE6WcTarZBMjMDiO50pRInycEBYoPA3YZ4qjwWdPTo1rIO3BZ4U5KZgmxjyES7w1GDiHUcHrZL9sV517ra7u1fnbxgKinmsS8gltolnx7Wa2HYlEb8/3+nAUXfqy0SOivem0NFjvzBAsPhECqPUyjOF9fDC4LdKoF1BikscaoJMPCvKa+RaHYPbkYAEJCABCUhAAhK4CIFerGAJ2q5fNViU9twP9m29S2IYg35ry0W44LMG1PBJG5iJQS+0rRnAQxuWQS+VE6P7ezym7ZwBMknWjfvzcjlPOZCk2pPmaVE5Ky6pRlmoCRtbEUgjVtTffW6NJXXK9pdLBifdkyE1qduY9i0CS5XNOrZL3a3LSUACEpDA7iagYLG7z69HJwEJSOAFIdCHf6p912h/3jkIC4z84pP5dNYwyNN5wvMBkaI8HyqZNF4VhIOqnBSERKLTwyfbKiGBbfK9RAe2Q8eNUrFyK9zT0MOwvleOB+rNviuJNZ+VBHw7z+qhMb+O80LMy/uB3+mgITKw7UqMzT75jkBCku2PpeA1wTGxHMsjUPC9vEJO9OtsBSMehHwisbZCxYXOhvMlIAEJSEACEpDA9SOA18P3DnaHePGBeFVcdj6HPowSOSFKuKicETV4BdGCibYpv9F2nEdMQCggVCrJsg91rWNUingvL+Y35XdElcubnhMyqpx6W7N4X2qQ9j8uFws8qdlzEnMv+wE3LTF3aw/nWCp8acu3ZqioyzsNLi0BCUhgtxFQsNhtZ9TjkYAEJHBjECjjfX3SAUJQGIZ+QljAcwKDPJ4F9Z13Ex0YRoKx3mtS3pKCYIGHAYZ9On2sPxQbykvifATOGf41WI9l+a1PbNg6deXBgXBA2CbqfaFE29W5Ot++hx1QOoN0Hqkz3/GKQIxgRBzHwvHDBgECoeLhft/sn3n8zT7Kfb7yX7RE24gUfcitc45dr4rzXQrOk4AEJCABCUhAAteVAO2/vz3Y46fz/VMp5RV7RZXpjfpNIYjBv9qz5W1Bm5HBPeyDgS20Q2lXUtJ+TKLs+EP07cvT8YBYpNwS0QIviWE7ftieHQ74GdR5++z8XSGmyHExHt+U1i/t/NRleXM0EgYqPZL5CBeIKNU+Zl/UcyPH0zykDRN1RZeGK0lAAhLY8QQULHb8KfQAJCABCdw4BHrPigpFVGGPeNfgOYE3BEZ5RIjykkCsoCBGMK+8KOhssc7dKff0y3Cgd/ZHOxQQqiNVXgdDIeNS4dApQkSoBNgIAtsFlvNti+UqN8b23hr1QmyohNp0GIlRTAxfclZwvHTeCG3FMnTYHkmp3BVsm/mIEpWzgr+HZV4eFSbTvtRT7XISkIAEJCABCUjguhJ4RfZG+KeafihfEA6u2VReF7XB3vuCNirtSdreLclESuV1Y/8IGbSBWYbvfFZIVparvGiEjjrrrVxeFU2UYI8X0DH4iWXaciT5zvbmcxamDVy5N9hPJROnvuWFPfR8vmac3JAEJCABCewMAgoWO+M8WUsJSEACNzyBgVjBu6U6RiVOYJjHFRxBgg4RnyTPJtQTIgadKAzzdGLowOB1QE6L16cQKqpyTtCJGU7DkEzVkdqen6KWv0hvqi3CeogB1I96U0dElsqJcb5zwLFWjGA6X+V6XyPE8AihQ4hYwW8k2WZEHd4bMKGDxnqEgkLIwLuCdfi93PzZfnUya18bESiualTe+Q7GeRKQgAQkIAEJSEAC15QAbddvGGwxSahHP5/CIJkv2NTnhMBTocJFIT5UDrkaTFOexc/03g60VWn30janDUzuiU60GCer9iRKRSXZpuYk2t4SJLY1s7dEjUqhRtO4jTeK+NEOezVbpc0PH7wqKuccC9Xgo/KQ/oJxcsMSkIAEJHBjElCwuDHPi7WSgAQksBMJ0LmgI8RIKTofdELKk4KE0nR8+B3jPJ0h5pEwm/mV04GOE+vhdUAoqFemVOxdtjtMJF2M6MxUb6hc2C+XH+9D6kFnibohmLC/i4kcdLdYj04fLu0IK3Tw8NQoAQaPCbwpWKbmEQqKY8KjAhbsA08MwgOwPIkSa9RdiRXw4Rj5e91QT5d7el1eAhKQgAQkIAEJXD8CfbJt2nh4Cv+TwZ5/pW//XXbuiiup/cDzgpwXFQIVgQBhoPLL0UYtjwva4QyqYWDRsQgS/B3fiMmB0WQly88GokU1k/tDGSbsLsFi6I2R/N4JB0UuDdq0tLOrr9Dl2OgGD5XH9JUcrutIQAISkMAuIaBgsUtOpIchAQlI4IUi0HtWVA6HGr2F0R8DfoV8QpyohNglZpS3BAZ8Okl0WvC4wKuC0E90lOjMYMynY8XydKD4pEOD8Z791mgxEDyfF8WFMJV7Orkktm/zYh4bJTLgHUFHi/oi0tA5rUTd5J8gzFMdN4zKRb9yUXCMhIuikL8DgaKEGLZbHcyFYsWFTqHzJSABCUhAAhKQwAtPoBcrqAhtvnv7NmBVDMGiDUxJwu3rWtmIF5Wou9rQ5SlMu7PCj9ZAGjyfT0ZcoP06i2dFknS3/BO3jqZrk9E8TdjlgvVyjEmqPRQrOKr6+5yk3E3YYD+0lytkLPNoO9P+pT3Mfp0kIAEJSGCPE1Cw2OMXgIcvAQlI4GoIbBMreKdUJwRjfbmU81mdIOLiIjowDwGjwjBVh44Yv3Ts6LjwGx06OlUY7Bl9hQfDcNruUXE1gkXVv7ZfI72GOTGoS707ER0QGB5KOZ6CtwQdMHqfeFQgftCRq3BP1K04DJN8c1wcZyXhZl32MxxlplCx7cT7pwQkIAEJSEACEriBCVSY0+8f1PHH8v23+jbeC1L1Ya6LgccF7fDKV0G9aJvShn02ggXzNyJOHE7LlAFIp0ezjS6c63LJMocTLop2e9dy5ZtW8TkAABqrSURBVB/ECsJF1TQUM6arrLeW7a3mc5Lts2AN+KmcGogktLMJadVCoPb1fkGYuVMJSEACErj+BBQsrj9z9ygBCUhgVxAYiBV0NCpvBR0MCl4PTBXCiY4PHR6M+S9OwXuC5Sp8Et4Yb06ppNqEWMJwzzrkvmD75XXAdq+VZ0Wdi6HQUS76CA0VIor9l2iCGFOhrcg1QV0/nlKJAslRwegwEoaXwMFxM2qMHBYIE2wLNhxfbZd1ynOkiTQm0q7T46cEJCABCUhAAhK48QkMvCsYpPPdKe8c1BrvCjwJboipFwFmEQXK46I8pqs9Sl27fHHjMaIE4UwJdYpwcbCJGYtF8ltEgCDHRb5FiOiODc+Kym9Rf/M5TROaPBizDRJ5b2S5CkVFe7gGPlWo1woPNcxZd0OwsxISkIAEJPCFJaBg8YXl69YlIAEJ7AUClbuCjhkjrni30OGpBHrDEVt0OMrgz3zECz5Zr5JyI24cT6FThKF/uN0arnWlnhSXcj4QRkiI+Mn+OF6dzwrdxH7p1JXnxO/l+/0pdOIQYBAwPtiv/9p8VsJwjoHcFBxTiTTlDs/2qlSeCuP3XsqZchkJSEACEpCABCRwgxAYiBW0V1+a8r8OqvYj+f6elOuSu+JykES4YPFlhIsSBpp3Q0p5Gdcnv9O+Z5ANntIHIjh04sZywUYiXMRjYpom7iyrL6Ne8PdKH711nnmb62nzjhFCPp3faDfTxmaB8rpm+5UUvDypbzhml8PXZSUgAQlI4PIJKFhcPjPXkIAEJLDnCfTeFeUhQCcDEYKOC52Vys8w/MRwj/iAMEHHBAM9oaEYodUSSafQacHwz/YQMeicsCwdJr7X/OL/fKJFdW4qtFJ5ezzf+cMD4sGU4309SnChLkwID+SswFvi3Sl4WLwxhXcqy9CJw8uC4+eYqSejxyj8RkeMujCSrDwsWJbCPMI/PV8d/V0CEpCABCQgAQlI4MYkQPsOT9uafjFffjqFQTltut75Ky4FUwkXtEcjXrAKDdJq79Mep51agkInWozHzE/IqBb3aX8+k5R7vYVxyjRtSbsX827AEcss5k/EG4NBQY9kXfoADPhhP9Xm77bX9Q/K00LB4lJOoMtIQAIS2EUEFCx20cn0UCQgAQlcRwJDsaLCQPFZuScQICoZNp2MO1LwpsCrAAM/y9KRQ+Dgbwz8hEyig/fKviBy0Hmh00OniLwXJT7QgRnmlriYhZ/12Q77HgTUPWeEWyW4Zjlc3UmSTWeK/SFg3NKvj+hA+KcHUj6cgscEx1ACBNvhOJmP6EGHCzGH920l02ZZ6g+jGjlmjorAcJKABCQgAQlIQAI7nADt369P+dnBcXw63x+OSIERfkdM28QL2sO0p0vAKM/g8jhej/iwiCBBP4DfTuRv2r8M3Lkp3heVlDvrjx/JPNrItP8rt90wt1vlrmNeG8izI4BZSQlIQAISuKYEFCyuKU43JgEJSGDPEBjmreBdQueCnA90VMhDgdhQxni8KjD4M4/1EATwTqDzQ0cFkaA8EzDiswzLsx6dFEIoMZoLkaNyYQC6klhf6F3G7+yjltsuarAvkmZTr+pgfSLfESLoWH4sBeGBjifeIOy/RpUhYrA9xAo6Y9SfuiG6sAy/s27lqihBozqqQ+8PjsWRY1BwkoAEJCABCUhAAjuXAG1D2oz/ff/JkdD2+6UUBr3syCnixZZoEM+LGuRDG7cGKJVHBG1i2ry0iXHRoNwRIYO2dDeAqAsDVZ7F1X5mwFJ5XFdY1BIrlibc3pGXjZWWgAQkcFUEFCyuCp8rS0ACEthbBAaJtkuMqPwVfGJ0xxOCd8uLUvCIoPOxPYk1xnw6Kxj3CQmFWMCyrFfeB4zKojDR6aHzUvFta4QX81mHUFSVN6MEisozgVcFnaBh7F22SQerPDv4m+NBYPizlA+kVL6J8vyoHBVsF5GF+iJW1LERIgqhAtGGevHJ3+URUvVqf5tMuz+zfkhAAhKQgAQkIIHdQ4D2JoLFlw8O6a/mOznPdsXgFMSDPkk3bXPaz7Spu8FHXQJtBvgw1WAkEnbTTq9QsTU4iTZ65a1gO4gerLMVIpXvvafH7rlCPBIJSEACErgkAgoWl4TJhSQgAQlIYECgPBVqBBRCAgb9ysdAZ4MO2+0pGO3xYiivCjopCBbMZzncwklKiEcF7yS2hcGf7THRealE3nRs+Lsmtkld6BhtT+xNh4n9EooKQaO8LSqJIAID3hR4eiCMUB/Eifen4GExzJeBkEGd2Q+CBfVhe7elVO4NlqlcG7UPltkaHdZXWrf2wQn0qwQkIAEJSEACEthFBO7NsZBcu6Zfz5f39e3FXXOYvYjQ2rR9rgvauxUeqkLFVlu62uuVS64ECdr9FWqKPkEJH7tC2Nk1J9sDkYAEJPACEVCweIHAu1sJSEACO5RAxa4tz4HWV0lBFCh3b37Dg4J5eBogBCAe0FHBo+IVg2UJx1Tr0dlBaEBEIN9DjVJD+ECsYN8sy1Q5LMrDo0SUGumFgMB+yxuC5RE16AwhVCCUEGqKztVnUshXQd4KOlXUmzwUHEfF12W75a2BuME67IMOVoWJqgSD7Kvi725xMpF2f+b8kIAEJCABCUhAAruIwP2foNna2q1flfLO/tDw2v1bfRtz1w5YGeS62Ix4UcIFbeMaTFR9h2GoVtrH5U1R4aHaIJ/yqEAI0btiF90kHooEJCCByySgYHGZwFxcAhKQwB4nUKGgqmPGe4RSCbcrXFN5OBAiitBPiAMsg0CBqzyeD6xHZ4aOCh4M1WHh+8P9by/rl0d4qH3SyaFTiLDA+hUOqkZsIUJQ6CxRD+pMHdhuFYQJxBS2Rd3oaSKU0HnCu6MS/bEfPCqGo704JrbNVF4mJZgMk4K3dRQqelJ+SEACEpCABCQggV1GoBcrOCrauHhY1PQ7+fLMTkq0fbWnhlwXERpq4M5wMFH1HyqM1NDzeauNPRQoFCuu9my4vgQkIIGdTUDBYmefP2svAQlI4IUiUJ4N5fFQo6eqI1IxafmbfA8IFHhiYPxHPLgr5Z4UklsjHJRYUSGfECyY2C6dP0QOvuO5UPsijFRN5emAmMCEkIGggRfE8ZQHU+7v9/OafhlCTyFg4HGBsEE9ESuo38dTyGPBMhUKCu8Mts88vlfnqzpkbJbjXpqjYuu8+EUCEpCABCQgAQnsdgK0O9+e8g8HB0pbkTbjnpoGHheGdtpTZ96DlYAEJHBtCShYXFuebk0CEpDAriWwLeE2ggUhkhAsykOCjhnzECb4neloCmIDggC/IQogCBBqCcEBz4nylGB51qNzx3zWwfOhwkkhSrCt4fLMY3mWYZuEomJd9oWXBKGeHkjBLR+vCOqDdwXLsTyCBoJJJfRGkOBvvC34LHf1cl3nGCv0UxMnUrYLFpnlJAEJSEACEpCABCSwRwjQvvzr24711/L3nhMs9sj59jAlIAEJSOALTEDB4gsM2M1LQAIS2MUEysMAIQBDP2IDHbYKqYS3BAID8xAZ+B1jP54LeDXgbfGi/vdK0If4gaBxZwriBuIH+SII28T+Xtlvn+VKbKAzSBJtxAm2fXO/P5YhLwXeFczHVZ/3Xi3LdvGwQKxgXyVKMK+SaFfS7MzaSgy42BbmyRFk0HGSgAQkIAEJSEACe48A3hW0Y795cOg/lu/v6tuOe4+IRywBCUhAAhK4SgIKFlcJ0NUlIAEJ7DECw9izfK98ERWqCQM/ggUCAPMQKsqTgr/xbMBrgvVYBtECjwhEA95JiB8sh5DBhBhAgmyWvy2FUFIIFAgkeE3gWcEyiBx4ReA1wTbpPOKhgTjBui/pt896CBUU1inRBZGCeuFRgRcFn8PE2eVNQZ12beJEDs5JAhKQgAQkIAEJSODiBPrcFbQjaXe+MYW2JxNhRX84hXaokwQkIAEJSEACV0BAweIKoLmKBCQggb1IAK+ChIUqbwI6ZYgTiAd8VmgkOmcUvBkQLjD6E1oJ4YJ3Dl4WiAYIF5XQmm2xPMICIgIFzwy2iSBBnovKG4GHBcsjOPxJCuGd2A+eGAgN7PtT/T75m/0jiJQYwn5ZB4ECUYKOJvut5NksX/k06rgqL0V+cpKABCQgAQlIQAIS2MsEBom28az4qpS/N+Dxz/t25l5G5LFLQAISkIAEroqAgsVV4XNlCUhAAnuOQOVrqATYJVQgIvBO4ZN5GP35jtBAOCZySrAOggJCAsIB4gBCBSGjEBUQEZjPJ9tCuHgo5Xi/LOsR4ol1ECyYj0cF6zKvPDgY2UZIJwQHOpKMfMNzg32zze25KRAstuelyKwugTZftoWAYpaTBCQgAQlIQAISkMAeIzAQK/AUviPlu1K+usdAKKhfTqFtOXrrPTRxnSQgAQlIQAISuFwCChaXS8zlJSABCUgAAogDTIgQhHOqZNsV5gnvCQQGxAGM/ogQlVCbdenI4T2B8PDSFEI24fFQHhyEd/pYygdSEB/YPttjG4gTLMu2mYcoQjgnvpPrguX5m20hVLAc6/G9vCmoN79X2CfyUpiLIkCcJCABCUhAAhKQgAQuSoD27lek4BH8TYMlfz3fGThjm9ILSAISkIAEJHAVBBQsrgKeq0pAAhLYgwTKe4JPRIAK84RogadDhX4qEYHwT4gEhG3iN0I3VYxffkNMQGQg7BNeDggJfJJA+yP9Jx4S7AuBAw8J/mZbFfIJMYT9sa3y4ECIoDCfddlnzcvXtp92LBEqzEkBEScJSEACEpCABCQggUshcGvfHsWFAu/fN6T8SMrvpzBAxkkCEpCABCQggasgoGBxFfBcVQISkMBeI9CHRloklUUlqy4E/I0wgPG/RArEAwQDvCEQKm7vS4WOKi8LkmojHiBEEMKJjh6eFwgZiBd4VLB9ck8gWCCOMA+vC5atRN61X5alHkOBgn223BR6Uuy1q9bjlYAEJCABCUhAAteUAG3SB1IYEPM3Ul6c8usJAUVb1EkCEpCABCQggaskoGBxlQBdXQISkMAeJVCeFggKlPJmqBBNeDtU8uphfgtEhvqb3/GkKO8IEmrzXkKoQITgOyPYbk6pUE4V4okOIb9XaCjml6dE1anlpegFCpZzkoAEJCABCUhAAhKQwNUSoO36oW0bMQzU1VJ1fQlIQAISkEBPoJKnCkQCEpCABCRwWQTiZcHyJT7g9VChnkrA4He8Lirx9Z35jgDBcggSJONG4GAiFjCj09gO8yrkFOszj7BPn+3XQxxhGwgUCBGV+2IYrkpPiss6my4sAQlIQAISkIAEJCABCUhAAhKQgAReeAIKFi/8ObAGEpCABHYsgUFoqGGIKESGKogN5K8g3BOF0FD8hsiAVwSeEiTI5ju/szy/sw4iBl4UeGsgWFRi7eY50W+D7wgVLSeF+Sh27KVkxSUgAQlIQAISkIAEJCABCUhAAhKQQDMEOUlAAhKQgASuiEAfbqm5WkS8KJECzwfm4QVBqdwWiA54VvA7wgWeF3hLIFaQ74KJZWvd8tpA3CAkFJ8lULCN+k7YJxNnX9EZdCUJSEACEpCABCQgAQlIQAISkIAEJHDjEFCwuHHOhTWRgAQksNMJlFBR3hYIDEMRo0JF8XuJEHhPIFowj1BQlfeikniXJ+Aw3FN9r/wUO52b9ZeABCQgAQlIQAISkIAEJCABCUhAAhLoDUSCkIAEJCABCVxTAn2oKLaJlwQF4QFhYrv3BCIFQkYJFfPea6PVp8+TUQLIMPSTiQ2v6RlzYxKQgAQkIAEJSEACEpCABCQgAQlI4IUnYA6LF/4cWAMJSEACu45ALzRwXOUpUcdY4kPLObGtNI2CEtFi1zHxgCQgAQlIQAISkIAEJCABCUhAAhKQgAQuTkCLkFeIBCQgAQlcFwLn8ZbY8pigAooU1+U0uBMJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACFyLw/wPP817hSR4OTAAAAABJRU5ErkJggg==" }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO3deXxU9aH38c85M2f2zGSy73tIWEPYZRVBQRY3rNpqpbW2eLXtvb1t7dOnvV3vc58+9npre7vXVq3WfSsqCFcR2QKyBghkJZCN7JPZ9znPHyMRC8KAUbbf+/WaF8mcOWd+c0i++Z3fdiStVvuSJEnXIgiC8BFUVX1LUhTFGQ6HrRe6MIIgXLwURXHLgHShCyIIwsVPvtAFEATh0iDCQhCEhIiwEAQhISIsBEFIiAgLQRASIsJCEISEiLAQBCEhIiwEQUiICAtBEBIiwkIQhISIsBAEISEiLARBSIgIC0EQEiLCQhCEhIiwEAQhISIsBEFIiAgLQRASIsJCEISEiLAQBCEhIiwEQUiICIsrhEajRaPVXuhiCJcwERaXucyi0fz7757mib+v5y8vreOPT7/A9KlVH/u4i+/8Kn94+iUqy/JHoJTCJUFRFBegisfl90jNq1T/+tpb6pTqcR88l1uq/v6lt9UJlYXnfVwlKVP97eN/VUsnLVB/8YuHLvjnFI9P/qEoikvULC5j9333p/z+h19j196Dw88NdLbw61/9hptWfOa8j1s+8Soadr1Ly74d2IsrT/ualKx8sjLTz/s9hIuPCIvLlDGliDJ7iG17Dp+yLRDwo1WU8z52Ucko2luaQQ2jSsopd6lKyizhv/7wGA/9/jH0mvN+G+EiI1q8LlPlE6dSv6fm1A2yji+u+ife+cuPzvvYaVkZHDnUh6SzIoddzLzuJjLTkoe3V06dz1BnI7bCyaz8yn30OwMf2t/v7ufN115HPe8SCBeCCIvLVF5eMR3tdac8L0kya554mK1b9pz3sW1JdrzuAdIKihnsaMPrduHUxk68AyXlFbz91MNMu6mUaDiEc2jwQ/sHva7zfm/hwhFhcZkyJFnw9536S6lGA2x9991Tnr9mxb1cN38av/7Jt+nodZ752KYkAp4AY6+ayuHaXeyr2XDSVpnbvvIArz7/AqPm3cG7616hud3xcT+OcBEQbRaXq5gKUuL3vM4pKECjNZFsM5/1tYpRRzgYYdb8+dRs2vThjbIGQyyGPyaTkWGlt2foXEsuXKREzeIyFQ4EMekTb8R8+lc/5XWrmSHH2X+5tToNSlIO5Wkqh44c/9A2SdYSUyMolnT0gV5cIdEycbkQNYvLVCDgQWc8ey3hhFgshs/rPeV5jVZHano68kmVFI0sMf/mO3nn1b8RPSULJEClcspsDr236R83CpcwERaXMkkmt3gUM+dfx4zZc8nNzRnuxpSI/5VP1NhZy7hv1coPPWfLLOLXz7zGjx95lB//9IcfHFvSsHDBTF555Q3KJ87i7i99Gb02/qOkxiKgarhm0RI2/s/aj/8ZhYuGuAy5RNmzS/n+zx4m5umlsb4BWWfkprtWkZaSxKa1L2MrGUPzO9sTPl5aTj5Bb9+Hnlv5jR+w+nc/4n9qGnjsuafRyhCOgSzLrH3+UZJLpvK97z9IfesgC68+wBtvbYdYmIDORlXBEP99qG34WBqtlmgkMmKfX7gAxHDvS/EhqT/50yvqvKuqT9lmtqWqt676X+q2pl71/vu+qOoVTULHXPqlB9XP3bJk+Pv0oir1zW171SSdrGp0ZnXs+PiQcZ0lTX25plktz0xV//u59eqY0lx1xX0/Vm9aMju+r6yoj64/oH72lsUfHF/SqD/5w/NqbqrlIjh34nE+DzHc+1IlG8jP1LNt+95TNnldDpLTs3n6lz/Aayzij8+tZv68WaeMsjwhq7SKf/32N5EkiZiqvn98LQ989wdIxNBqNURDXuoOHARJwwP/9nNSrTJX3fhFOna9xqGWTvRJZgKe+MCrhbffj+LvYcKU6cPvMeW62zF5Wugc8Iz0mRA+RRqNRvPdWCymv9AFEc6BGmHUtCVU5lpoaGggHI6g1RmoqJrG1773H4Q7d/Pb3/yBfTUb2br1PZav/BpfuGclcizCkGMQvz+A2Wrn6uW3883vfIu//voh+jxww9L5bN5Uw93f+CnKQC3b6geZPj6fPXv2k5ZTzNd/9DCKo47usJUFMyfyowf/BV8wQlpuOVMnlmHMGsPnb1vEP6+8ndm3f51MYxhb3li++rV7+fG3vo7HF7zQZ044TxqNJiQpiuIKh8NJF7owwrlRDBZu/cL9TJ8xDYNeRyjgpfnwfta+9AxNLUdPeX1GXimLbryV6smTsdvthPxuands4vm//oV+hwskDXd9/d+YP3c6Nete4LFHH0NSzNz7zR8wbUoVHkcfbzz/GOvXvc3sZXdiDnXx5vp3AJB1Zr70z9/BiJcn//hrHE4veoudz937AKkWLc88+ms6u/s/5TMkjCRFUdwiLARBOCtFUdyizUIQhISIsBAEISEiLARBSIgIC0EQEiLCQhCEhIiwEAQhISIsBEFIiAgLQRASIsJCEISEiLAQBCEhIiwEQUiICAtBEBIiwkIQhISIsBAEISEiLARBSIgIC0EQEiLCQhCEhIiwEAQhIbKqqiIwBEE4I1VVZTkWi2kudEEEQbi4xWIxjahVCIKQEBEWgiAkRISFIAgJEWEhCEJCRFgIgpAQERaCICREhIUgCAkRYSF8qpJTUj9ymzkpCa2inHF/e2raSBdJSJAIC+FTVVBU8pHb8gs/ehuA0WTGlmwf6SIJCRJhIZyWPSOXsnHTkeVzH+ArSRLjJk4mJS0DjeaD/RVFRzAY/Mj9tFotkXD4I7dnZufS3dV5zuURRob2QhdAuPjoDCZmL7mLMVPms/rxn3F418aE9tNotRSVlJOemcWQYxB7SipJViuZOXn093RTUl7B4QP7hl9fVjEGa7Idl3MIo8lEZlYORpOZYDBINBohHAphNlsY6O/DZDZjMBrJKyziwN5djKuaTFdHGzn5BfT39tBQt/8TOhvCCaJmIZxi9KS52FIyiISDVEycjVarS2i/aCRCacVo9AYjOr0BraKQW1BM7a7tpKZn4HIO0X08XjPQarXIskxMjVFUUkZ3ZzuDA334fF5S09I5VLsHg8FINBolPTOT+oO15BUW09fTTV5BEX6/D6stme7OdqRP8mQIw0RYCB9ittqZtmAFBlMSO956kYqJs0jLKfzI12dk5VA6ajQWqw2AcChEIOCnq/0oBqMRx0AfwUAAg9FIbkER0UgEAEWnJzMnF7PJgs/nJeD3k5Kajts5RFdHG5Ikk5aZics5REpaBqnpGRxpbECWZYLBAG7nEIpOob+3B6dz6FM5N1c8WZb9gCoe4iFJkrrg1vvUf/vTRnXy1TeqFluq+rWfPafedO/3VUmWP/Raqy1ZXbriDnXCpGmqRqtN6NiSJA1/bzSa1DkLFqv21LQPnj9p+4l9Tv73dNvE49N5yLLsFzULYVh6TjFTr7mZ/u426t7bgNc1SMvBHVROmkN24ajh102YNJUvPvCv7Nj8Dvv3vDdcWzgTVVVRVXX4+zFV1QT8PhwD/R88f9L2E/uc/O/ptgmfHtHAKQxLTstCUfTU79lEwOcGYPfGvzNu+kLGTLmGrtYGlq24g/TMLH7z85+esefibA7u24PeYBipogufAhEWAgAarY7qOcvwuBy01O0cfr7v+FE6WuqYcNV1pFog4HPz2O8eOaUWcK6CAT/BgP9jllr4NInLEAGAnKJKysbPoK2xlu62JiA+CMqSZKVm3bOMKi/CnpHH35978mMHhXBpEmEhIEkSVbMWEwkHObDjLUIB3/Dzik5HJODEpJeRzLkYzRaKSkeRnpl9gUt9+TGazEy5ag45eQUXuiinJcJCIMmewbjpC2msraH5wPbh5yORMFnZudx8+128+LfHKakYy3Prd/CtH/5fLEnWC1fgi5DBaPzIbTqd/qz763R6/H4ftbt3kJKegaLEx7ZIkoROb/jI9h2D0XR+BT4PIiwEJlx1HYqiZ/fGV5FQsdlsFBQUMKm6mmuvX07v8U6mjClgjNXF1jdf47tfuZ2jzQ3IIAZEva9yXNVHbisfPe6M+8qyTH5RCTqdjuppM2lrbSErNw+AlLR07CmplJRVnHa/klGVH6/g50A0cF7hFJ2Byuo59B0/iqOnjfz8fJYtW8aMGTMwGAyokow95RroOkRo3yvMkbyoEwz0OT0MBKDXD0dcMBCE6GXalFExdsJZh5Of6BlKTknF5/UQen8OjEajQeXMJyYWiyHLMiaTGadjEAmJYDAAQHZuPvV1+087Wzc7r4D2o0fIKygiGotyvKP9fD5ewkRYXOGyiyrIKhzFxlceBTXK4sWL+eEPf0hqavyHMxaL4XQ6CRTn0aaT0fS3U5GfhU1tpsASDwhfGNo80OCENje4wpzl1+PSkVdYDEBuQRH2lFQCgQB6vR6D0URTfR3FZaPoam8jLSOTMROq8ft8SJLE+OqpdLUfY8bca9j01ptcvWgp9QdrSU5Owe1ykmRLJuD3c7SlEQBJlsgvLiXg85GTX4DH7WLsxMlEo1FSUtNxDPRRXjmWcCSM1ZqMqsYIBYN0tbeRkZlNks2GTtGTlZvHvl3bKasYg8ftwp6SRm93F1m5+QwNDnCkqf68z4VGkqTvq6oqQuMKJEkSs5fcRXpOEW8+80vKS4r49re/TUVFBZIkIUkSsiyjDXswhF2kmLRYXa1kOOsp1ToYZVWZmAqjbFCVBlPSYGwKWLQQikEwBtHYpR0c2XkFaDQaSsoq6O7qYNSYcWzftIH0rGxikQiD/X1IsozNZicSiaDGYpSOqmSgr4eUtHTcLidms4VYLIbBaCQUDJKSnkFBcSlN9QcJ+OPdxxlZOWi0WoLBAElWG3mFRXR3dqBVFExmC73dXUy5ai49XR0UFJficbtQVZVYLEp2bj5ZuXlYbcn4vB6MJhPhUIjklDTsKalEoxEkSUKj0dDXc/y8zoMkSRERFlcwvdHM1Td9iZ62Bo7s38z4ceNYsWIFFrMZjTb+I6GqKqpGizMs4ZKM9JvtdKZa+Hv9Lp4/EubpJtjXC4EIZJthchoszocVJTA9A2w6iKngi8RrIZdacJSUV+AaGkJRFDrajqJoFQb6eykoKkVvNBEKBbHZkmk4dIBkeyoajYZQKMjx9nYysrLJLyymv6+XjqNHyM4rwDU0RCDgY8gxQHdnJ6oaA2B89RSONB5mfPVUDtXuQdHp6enqiIeSqqLVKoSCQbSKQltrC0k2G3q9gdT0DAC8bjc6nR6XcwhF0ZFbUEQ4HOJoSyNZOXk0Ha5DZ9DjGOg/r/MgSVJEkmXZH4vFxFC6K9CEqxZx61e+T/ueNyjKSuK2226jqKgIrfaDvx2qqhKNBomhoqLSdPxVBno2EDiwF0frHkYXgtcH3YOwtw56joHqgjwTTEiFsXbwRGBjF2zrhr0D0OGN1zwuBYqiIxwOkWyPXz4gSUQjESxJVgJ+H5YkK16vh3A4jKIoaLUKWq2WgN+P2ZKEz+cBFXR6PT6fF42sIRwOkZKWzmB/3/D7GIxGAn4/er2BYDCA7f33s9qSCQWDRCJhzJYkXEMOotEoOr0eo9FEMBggGAigVRSikQgarZZkeyrT51zN2ldeIMlqxeVyosZiyLKGaPTsQ/NPR5blgAiLK5Asy6SnZ/Clb/+cysoKsvVuqqrGYzAasJgtQPwSBU6Mv1JxB8P4AgH+9srLDITrSC9qY+t/rSXX5CbZDLnpYE+CigLwemFbLWzaCpogXJUJywuh1QXbeuCQA2p6wRGEQPTCnYczMZrMJKekMtjfSzAQuNDFOSeTps/E7/Nz+MDeETumLMsBcRlyBdHpdOTl5TFp0iTuufcrfOGu26gqz6astBiz2Yxep0dVQZI+CAveb8uXYlH219byp24TO//4Nyqn3Ym28Dhrn2/H7VXRytDvhIZ2ONYDKclw72egOwh/roG32qHUBgty4jWNUTbIM8cvUfwRCF9ENY3islFk5xbQ3toy3KtxKTFZLHS2HSUcCo3YMUWbxRVCURRyc3OZP38+99xzD3fddRdLrl+M3WpGp8QXoZEk6f1Ljij+QIBAKITu/cVzJaCnp4df/uIXHLCV0fnmk4wZu5zUwkw8mmNsXNPP4XZweiEYBqMBAiFoaofpY2HpbHh5F7zYGB/YsygfDgxChhEq7TDGDnknelYiELmADRvzrr2eaDTKgb07iUYv0mrPWTgG+kc0KCAeFiIkLmOKomC325kyZQqLFi1i9uzZ5OXlkZ6ePhwOsViMSCRCd3c3jY2N1NTU0N3bS3ZWFvOvvhpVVamtrWXz5s28/fbbRNKnYS2w0NryGtbM66mYUkZDTS+tewcZcMHuJsi0w6i8+MPjh6pSePWn8IsX4d16kDphVjb8oQ5GJ8cbQUfZoMwK/YH4uI3DQzAY/PhtGxqNJuFf+uW3fo6m+jrqD9Z+vDe9TIk2i8uQLMvY7XYKCwu55ZZbmDFjBnPmzEGj0ZxSi6irq6Onp4eHH36YY8eO0dnZid/vR1EUUlNTsVqtuN1uHA4HXq8X3Yqvk2oYpNi3nyVf+DID/bVgbOKl/6hlsC+KX5NGLBJF6m/HpFcpyYJxxTB3AiyYBOt2wsGjMNcOySH44bvgC0J1CmSbQPf++r7ucLxNo8MDza744K/QOXbDmswWVFXF7/Oe9bUz5lxDXmERLz71l/M655c70cB5GVIUhYqKCiZMmMDKlSuZOXMmJpOJaDSKVquNh0RMJRwO8/hjj7Fx4zvs2LGDnp4eQqHQ2ReVSctD/+X/h/lv/8LNX/4S2WVJOANv0R3JxZk0Bk/AQJ8/hb6dB3E98TCxqIpegfIiDbfdlMTyWRIHDoXo7Y2QJ4WYYFD5/S5YfwjwQ7YBSpMg3Qjy+80mMRX6AlDvgDoHOBKsYReWlHG8swM1FiV8mrU3ZFkmFouRV1jMDZ+5k9/+57+f28m+goiw+AcWA3gurYbvYRqNhqysLCorK1m5ciXz588nJyeHcDgcnz2qKIRCITq6ujk6KLF+7WrefOFPNDc34/f7z2HlKQnN0lVI6flUO48w75bb2ejrpiS3heiet3B39oOsQZ39ORzPPYrP4SetwMzoWZl4BgJoPB6m5IeYNV6i26VBGfRQ0jtAS0+Ev9fDzkbo6gazDJkGKLFCkhK/VIF478nO3nibhyv80UPMzZYkps+ZT1trM831h077mszsXAYH+vjqgz/g9//1fxOqgVypRFj8g0VTYN2uC12KcyNJElarlaKiIm699VZuvvlmSktL0es/mOkYCoXo6enh5Zdf5rhbIr18Jr/4zufoams+jzeUwWhBs/x+lGlLyM7Ox35oM13PfoObv10JqPR3BvBNuoPK0DqMZpmeVjeHt/RS9+5xvEMhpGiU+5bDF5drqDluw1iSQc6hVoo1QbZ1w/4eaD4OB4+A3wdyNN6mUZwEme9P7vRFYE8/HHFDj//U3pRrrr+B9MwsNr+9jkgkTNDvxznk+NBrSsormbtwMbu3b+HA3kvsP/5TdsV3nZr0ED6p7WvxFNjVEP9aI8P4YugbAo2iDF/nn6A3GBJae/KTZDKZyM/PZ8GCBaxYsYJVq1aRk5ODJElEo1FisRiBQIAnnniCZ555hi3bd1EwaSnNh/exbd1z57mIjQqqitrVTKz1ACXJyVSWjqG97jBbnt5ByBsiqyyZQ+ab8L7zOkd29uBxBNEZNGQUW8kYV4CSV8S2eoX1G4a4rtJHWlKU+rJxvPLGABPNEeYUQYoNcnMgMw16vdDkgPpB8EYg3QI5yVCVCdWZUGyFSAzcQQirkJtfSH5hCVs2rOeWz66k8dBBMrNzGTOhmszsHByDA4TDIcLhEFk5eXR3drBw6U0M9PXicbtG+r/psnDFj+AsyYKcNKg5FJ/DcMd8eH5jfJzB3Algt8DLW+LTj5sOH/xQq/rYqsnU1e6+IOVWFIXMzEwmTJjAtddey2233UZaWhqxWAydTkcoFMLn89He3s7TTz/NW2+9Rd2hQ4yePJ8ld32Tx/7fVzl+9PwnFAFgMCNlFmOZMJvJN9zL8fYmmre8Qex4C2pfO8rKnxJ94n+jD/WTkm3CVlFI2g0rMJtiqK4+VFs2rsPNdL+6msWj3Nxxh50N0TIe//YuKsxh7psBZTmw2wFdfrCY4pWashxIM0HQCYoLjCoY3v9T1+aA5/dAnTyZ/Qfq8PgD8bktWoVQKD5eIie/kAXX30A4HOLtNavJyMrGaDLTULc/PkJTOC1ZlgNXZI3ihCPdEIpAeS6U5kCqNf51vwuMevj7tvjrTtQq0jKy6O/tBkCrxE+d2ZKEz+v5VFab1ul0ZGVlsWDBApYuXcqUKVNIS0vDZDINl1FVVbZt28a+fft49dVXaWhoYGBgAFmjMOO622lrPkBP+3lcfvyjgBe1qwlvNIy3spr8MdPpaq3Hl5YD0SjIWuSlD+B/7TccN1TimPNdel76JSmO3aTm6rGkmrHNvIGkhZUc7uvlh4+5mDGzh+88OpWM3btwOsIYClSWjwFZA9ooNPfCoQ5Y2wT7W6GpDaQITMuA6gyYXAjfva2S41ELO3UBXAEYDMaQCdIwBB0+aDl+jCf/+N8kp6Sy5ObbiEVjvP7SM+/XKCRAxZyUhMFgYqCv5+Ofp8vIFV2zOGHhJLi6Cn7/Otx5Deyoh40ndbWPHj8Rl3OInq4OJs2YzZHGw1SOm8jxjjaKSsvZt2vHJ/qDpdPpSElJYdq0acybN4/ly5dTWFiIctIdx1VVxeFwsHfvXh555BG2b9+Oy+Ua7gXIzC9j1Y8eY81TD7PrnVdHtHxF46Zz83d+y9q1z9J4tAkpJRvJkow8eTEYTKhDfUReeAi1bivEwugMGsx2HdmLF5JWnoGueTOSDGoMiifaKbBrWPfL3fidQXoGwSzB8nEwrwIqsuOXiBop3hgdHAKdBxxDIMdAXfQg0t5fUZEdoGZn/DJTK4FZAYsS72HZ0w9/PAx7+yEjO5dbP38PzfWH2LD2NfRGIxmZ2RxtaSIWuzQHZX0Srug2i4xkqCwAoy4eFn/fBk2dsO0Q3DYPDnWnUVYxmoDfj9WWjEajISMrh7ravRSVluNyOrAkWXENOTh2ZAT+Up+GoiikpaVRUlLC0qVLue+++7jhhhvIyMhAq9UiSdLwjYZ37tzJk08+yRNPPEFtbS0DAwPEYvFWv/gam0soqqzmrRd+h88zstVtv3uIyVOuxhhwc/iNJ+KXIj43an8nDHRC91GklCwkexZqOETU7SLgDDLY5aNv9N0MrXkJk1VB0kh4h8JYi1LRZlk52i3R3RmgZyhGTSusPghvt8KmY/Eu1PYQNIehQYXNLlgfHsPuHg2/W30AjR6KyuCduvjEtWMeaHLGH1oZvlQJs7Ngd7ubN9/ZjM1up2LsBABS0zPoOHZkRM/Rpe6KHcEpATotuL3g8kHdMchNg/1H4qMO/cH4kFnHQD8arRaD0UhQktHp9diSk+PDn493kWxPITe/CI1WO6KNnVqtluzsbHJycli4cCHLly9n7NixmM3m4dfEYjF8Ph9NTU2sWbOGLVu2sHv3bhwOB5GTyhJfdFdP9ZylHK3fy2DvyN+FPOj3cXj3RiZffRM2mx1Hbyeqsw/1SC1qdglS2WSkJDtSdgmarCJURw9qRwPRtkOEjBn09GnpX92GMUkhp8KGX5tO0Y1LKRttJHtXDV0bttNx2IHXHWZfS7xmYTZASQ7MmayQk6VlVJrEddNuYcfr/4mzHH6zHf4lG4wV8PS6+EjRbBPYddCvwvr2eLfscwvhhSMqf9i3lbqYjqWfuZN31r0x4ufocnBFhoUKdJw0rf9YD8weB19ZCjoFXtwEN86EDXvB7Y/Q2txIOBQkFouh0WppqDtANBbF43LhGBwYsaDQarXYbDYqKyu56aabqK6uprq6muTk5JMmdoHX66Wzs5OnnnqKnTt3Ul9fT2dn54dCYvizqiqpWYWkZxey593VxM5zivKZqTQf2M6cZXdTMmYKu3s74z0tAS9q6wHUrhak9Hyk4glIabnxy5SUbNSi8RDwIo+eRXTXWjxemdb8u+kuWYhzzVMsmu/gQHoqRVNzyR9to6PByfEmJ5IsUVKdytRl+ehsWrr63Ewuuxo12MSC27OZ1OXl0NY+2gZUPrsQdh2D9XtAB9j18Wnzlcnxlb2OumFBLlxfAG9IVai5aawd6n2/9UI42RUZFifTK7CgGn67Oj7FWqeF44OwYR/Mq4I174FWq+B0DJ62EdP1D33350OSJEwmE2VlZUyePJnPfvazzJ07F0VRPvSeHo+Ho0ePsm3bNjZv3symTZvo7+/H7z/zzXoqqmejqiptTWdeR/Lj6O1sxTXYy6iqWezd/MaHQynoQ+1oQO05CvYspKxi5PxKpCQ7ancr2i/8FPXqOyA1B7VpN64f302tqw9dSz6VX7gRKWUUJn87VdfmYDArSDI0vtfH+j810lk/hM2WhuH+LB5/5FcU50ncdEsKFTMzadzSzdb98MgD8PDzsLMhfqn5Vhe81xcfs1FujQ8rX5ALt88r4M1NT3NnWfwyp8kJAwG4iCbEXlBXbJvFCXol3rLuC8ZnTN44E2pbIBSGxo74H8jislH0dp/fcmRnoigKVquVadOmkZ+fz/e+9z2+/OUvM2rUqOGh2Sd6OTo7O3nnnXf42c9+xrPPPsvevXsZHBw8bW3iZDq9kcV3/gvtTQd47+2XP7FGu1AogN5gpmrmYvZtXUvQ7zn1RbEoeJ3Q24bafQSG+iAcRHUPgtECHY2ovceQ7JkgK3Tu66KhxYg/qxr/nhoGu3z0t3vpanDiGQyhM2iIxeDWz97P03/+PX39bjp7VbZu95O7oIxDB7w4+kIoWlh2Vbx7fFxR/I/CgAeOOaHZCQcdsM+hYfzsRVR2rac/AAWW+GxYvSY+oS14hSeGmKJOvLU8+P60gZgKdUfj/55sbNUkjrY0jdh7nhiaXVVVxT/90z+xcOFCHnzwQcaPHz/cDRoOhwkEAhw9epTnn3+ehx56iNWrV7Nnzx7cbnfCMyPkyHMAAAzQSURBVCmrZl3PxFlL2Pjqn0emy/QM/F4X1XOWotUqNNe9d4ZXqhD0w1APas8x1GOHUPvakdQoGJPi7Rs5pcgFY4gZ7QxK+bQ++TJH9/TiHQoRCaskpRkxZKRSfc01mNNttB3bQTQcJRyKEg6pdHcFKZhbyOvP93D4GFSXQ4o1Po0+Jw1GF8RnxwbD0O+GMXOXsWFfM50d7dxeGp/1qpUh3wLltvjcFNfIzvq+pFyxDZxnEjnN7+CZbiBzLiRJIikpidzcXD7zmc8wb948Zs2ahaIow8vBx2IxBgYGOHbsGC+99BI1NTW0trbS39+Pz+c7p/fTaBUmzl6Cc6Cbhn1bR+QznElPRwvNB7YzdvoCNr3+BD730Nl3CvrilylD3USP1CJlFIAtDTm7FCx2JI0WuXI68uwVxJr30NHaTrfHQN+cB8jKjLCkvJQNxzZRsvI28neuZ7DTS2e9E8dxP/ZsE7ZCGwfqnXz+Z/DST+Jdpw0dUJoNYwvj42s6+6Fi3jT+zw9+xM5QfIr8v0+D39XFi1hija/09T8d8XaOK9UVX7NIxNRZczn4MecOaLVaMjMzKSoq4utf/zqrVq2irKxsuAtUkiRCoRA7duxg7dq1vPzyy7z++uvU1dUxNDR02lmTZ1NcOYlZ19/J3i1raDm4/ew7jACNVmHCVYvwOAfpaKlLfEdVhXAAhnqgrx26j6A642tUnmjjwGxDM/sW5CX34373TSwb30TrCfDeS39DO2kBBkcTFptMVomVrJIkfK4wE6/Lpb6mF583xps74PYF8cF3T78NihL/uqiklIx0K5nSHtKT4b022NUL/zwO3BHYPxBfqEcG2r0X16penxZxGZKgydNnUbtrx3ntK0kS6enp5Ofns3DhQn71q18xZ84cFEVBluM3hFNVlfr6ep566imeffZZ1q1bx5YtW3A6ncNjJc75fWWZhSvuw2S188Zf/xO/131exzlXQwPdFFVMJL9sPPtr1hGNnHvIocaQQgFURzdq9xFih7ejmXA18tiZoDeiNuyAcIg7brqFF158me76dgZHrWDw3Xfxdg+iN2pRdBpkjURRVQrW9PiYQ18QVr8bYXwxfOv2+Bib3iGYfv0qKniSpVODpFgg1QZBDbx6BOZkwGgbvN0Vb/R0hq7MBk9xGZIgjfbcT9OJHo6JEyeSkZHBN77xDcaPH4/NZgPiAeH3+3E6nWzZsoWnnnqKtrY2mpqa8Ho//lTp/NLxVE6aw+53VzPUP/KNsx8l6PdSu/VNlq38FuNnXHveo0WHe4FCATjeQvjnnweTNV7LqJxOXm4eTq0Z95j5yHnjCRtS6Q9l0negla5GF7Z0A2kFFrQF5ZgXzqW0qI3Cxt14ul08U+fiiXfdTCsJM3+yhc5+ePpFJy4flGRDkhGmVUCwFBq84O4Djwo9vgu75N+FJmoWCbCnpKEoOgb6ewHILyzB43Z+5HwQvV5PRUUF8+bN4/7772fVqlWUlpZiNpuHeziam5t5++23eeSRR1i7di1bt26lq6uL0AisnajV6Vl297fQGcy8+ui/E/R/uus0DPZ2kFsyhlETZ1O3821CgTN37SZEjUHID45u1LZ67rphGa+uW08AGSkpBSm7BCm7BICw24dnKIxjylfoSL4Ge28NlqxkfHkzMA3Vk5pjxF5oo92lw17+Vf70p+fYvGuQluPgNFgZfX0xE2alUlJpQfUGMeojWJKhzwVDV+iSF6JmkaAdWzay8r5/pvHwQQDmLFzE83999JRLBI1GQ2FhIaWlpVx33XWsWLGCwsLC4TaJSCRCOBxmx44drFu3jg0bNtDY2MjQUAINgefAnp5DUWU1uzb+HfdQ39l3OJ0Tg8DOY4Jc0O+ldtub3PKVH1BQNoFDu945vzKcjqqSbjUT7e+kf8MLYDAh5Y4CgwnN5EXQ34k84WrkMbNQu5rx/PKbbI8NsPKhKRxTPo/fmY1pqIHUXDNjp1aSPz6J8W49k40TyB1lw+MI8vqaDh5rdJCsDVGeFSU/Ld6TUp4H7X3xLtgrkQiLBHg9bvx+HzZ7Ck7HIJYk6/CNcCHeeJmSksLkyZO55ZZbqKysZMqUKeh0OiKRyPCYCa/Xy/r163n88cfZvXs3fX19590m8ZEkiaqZ8RWq97y7+kO1H41WQaNVMJqtaLUKJmsySbZUQMJsTUar6EGSyCsZg8GUhKzREPB56G5rIuj3EIvF8HuchENBggEfbkcf0WgEr8tBLBohEv6gVtS0v4a+rqNMnLOUxtptRMIjt6T+Z+6+l+f/+ihEQuAJoTbuJHq8BcmYhDzjBtDpUQ9vJ3b8CJo5K/AfPcBff9ZK6RdayLhuIeMiQYwWheriz3PMvYaKGRn0tLpp3NHHkb0DdBweIuCJ0BVVaWiFlKT42if+K7jrFERYnJEsy9jsKaSmZbB+9UssvvFWXn/xGSLh+EAojUZDeno6M2bMIDc3l1WrVpGXl0dycvLwMRRFoauri9bWVn77299SU1NDT0/PWUddni8JifScIqLRMKMmzqJkzBQUvZG0nEJyiioxGC3oDCYUnT5+j7FYDEmSCYcCaDRawuEgPpcDrU6PLGvwe90UllehMxiJRiMoOgOxaASNVgEJopEIQZ+HYMBHb2crPe3NBANeUCESDpGeXTjckDsSyivH4nY66e/p/uBJVQXXAJE/fgssNkjOQs4qQkrNBWsqmsoZBEITqTusQ+fJ4NCr9ZQVlTE4upZXX1xDVmkS6eOLMKQXUTxFR8E4O4NdPrqbXQx0eOlzitmnIKaoJ8SclMSC629ErzcQi0XZvX0Lfo+L2bPjw6i/+c1vUlVVhdFoHL7cODFmorGxkeeee44NGzZw8OBBPB7PJ34/irFTr2H6tbdhz8gh6PdiMJoJBny4Bvvo7WghFPQT8HkY7O3A0dcFSEiyRCQUxO91Ew4FgfjaGLIsI2u0GM1W9AYTsVh8BS6LLYXsglHoDSYUg5H07CIsthTM1hTCoQCKTo/bOcDhXe+y+fUnRuyzTZo+i7p9uwkGz7JYqiTHG0TzKpCKxiIlpSLpDMizboH/+QsPLpnDz3/yvwl6PSjL78OUmUqmbxe27hqSrCqKTkYFfM4Q+9Z34Rm89G42NJLEGpznQKPRMHPeAopKSgk4BygvL+Oee+7BYrGQmpr6wcrZ0ejw8Ow///nP7Ny5k6amJtrb289rrMR5l1erYDBZiEYiqGosfo+QaGT4+5EkSRKyRht/yBpQVbQ6PaGAj3DoIlgBWW9GyshHyipBs+JfWZQUpKurkwNhI1JOGbG6rURe+Dm4+tDpJSwpejIKLWQWJxEJx2jZ3U/fMQ/RK7grRIRFAjQaDTabbXity5kzZ5KZmTncJiFJ0vDoy0gkws6dO9myZQurV69mcHCQpqams87fED4lWgXz+Fk88NAf+WXdADGfG7VxZ3xuSjSM2naYWM8x6DmKFAuTlKJDb9biGQzid1/Z/4ciLM5AlmXS0tIYM2YMc+fOZfHixWRkZFBYWEgsFkOSpOG7jfv9fo4dO0ZNTQ2vvPIKO3fuZHBw8FOtSQiJue3ue6k7uJ+6hgYwJyNlFiJllyJZU5FkTbwWNnAc9cg+1I7GeCOqINbg/ChWq5UJEyYwY8YMli9fzpQpUzAYDMOrZrvdbux2Ow6Hg97eXnbv3s2aNWvYuHEjfX19IiQuUiazhfyiknhPCoDXidrfgXqkFiklB6liKpItHSktJ77eRmYRsQObwXcFTwg5iQiLf2AymaiqqmLZsmXMnTuXzMzM4cuNE92QLS0t9Pb28vLLL9Pf3897772Hw+EYkQFVwidn2Yo7eO3FZz785PvT5lWvMz5tPjkTuXwyki0NNRQAoxl8LsRSOCIsTpGamkpxcTFOpxOXy0VKSgrBYBC3201bWxt79uxhzZo17Nmzh0AgwNDQ0CV7t+0riTXZTnZewQe1itMJB6GvjdjgcTCYIRqOT6UXQQGIsDiF2+2mv78fWZZxOBxs376dtLQ0Nm3aRHNzM62trXi93uGFcoVLw7VLb2L1839L7MXRMHhHdlTt5UA0cP4DRVEwm83k5uZiMBgIBoN0dXXhcrlEr8YlzGA0EfCf23ogwgdEb8gZaDQaYrHYp3LzIEG42InekDMQ7RCC8GEjN2hfEITLmggLQRASIsJCEISEiLAQBCEhIiwEQUiICAtBEBIiwkIQhISIsBAEISEiLARBSIgIC0EQEiLLsixmRwmCcEayLEdkSZLETClBEM5IkiRVXIYIgpAQERaCICREhIUgCAkRYSEIQkJEWAiCkBARFoIgJESEhSAICRFhIQhCQkRYCIKQEBEWgiAkRISFIAgJEWEhCEJCZMRdXwVBSIBWVdW3FEW59kIXRBCEi5eqqm/9f/X/HNdwOa1eAAAAAElFTkSuQmCC"}
,{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"QXRtb3NwaMOkcmU=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydB5QU1fZ3/z5zzhkUEwqSxBwxJwwYnznnnHPOOWfFLGZQDIiKoiBIBkEBUcEcQBQDoqJ+Z8+r8iuanunuoQeGmV1rndXdVbdu2HXHJedX55z/+z8PCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAIzmMCsM3h8h5eABCQgAQlIQAISyENg3vnmX6DRSo1XXXChhRf5+acJP/7z999/C0oCuQQaNlpx5VZrrbvBqqu3aLXk0ss0mHW22Wab8OMP42sbqUUXW2LJ5VdcufGcc841N/u5ts0vO59FFlt8id8mTvy1Ns/RuUlAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISqHECoVMseNnN9z7Sb/T3fwz6/Kd/sJ7Dv5xw7BnnXzbbbLPPXuMTcICZgsCOe+xzYKfuA0akeyT7+eaQ0WNPPu+yaxEJZvRiVlh51SYPdHy1Z3Z+L/UeNrrtrv/db0bPLd/4q7dsvfbAzyb83XyNtdatjfNzThKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEpguBWeK4+/HOr/cc/tVP+xx69ImrrLZ68+at117vlPMvv27AmB8mX3fPo89Ol4k4SK0lwB658Lrb26dC1lmXXXcbzv/W62yw8QZtttim3V4HHHrDfR069f1k3O8IF+tuvNmWM2oxRCq8PnDU1517DB61Zdt2u6+4ympNmc9N9z/ZmfnvfchRJ8youVU2Ln93zG2dDdtsXtvm5nwkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUw3Altst9OuOEu33nHXPXMH3WXvAw/j2va77LnvdJuQA9U6Arvvd8iR7IOLrr/j/nnnm2/+yiaIOPD06+8O7f3ht78S5TAjFnLmJdfe0uej735batkGy+WOf/kt9z2KqLJsw+VXmBFzq2zMi2+48wH4LrTIoovVpnk5FwlIQAISkIAEJCABCdQXArPUl4W6TglIQAISkIAEJFDbCVx/72MdqUWw44YtVvonjtz53t+xa4+55ppnnn2233jN2r6Wujq/BaKoyJrrbdSGehHxhP755qvPP+v91huv/vHH77/nrnmOOeacs9Xa621InYn4Otf4ceO+6/tO924/fD9ubHX5vNBzyEc/jP9+3EHtttwgyppUWdeEcZ96tfeQDu3vuPnWqy8+p7pjVuc+IkGI8Hjr9S4vXHjK0Qfn9kGNltcHfvT104+2v+uGS845tTpj1MQ9j3fpMXCBhRZeuO36zWqVkFKdtZayV3le/Ldn1abNW807//wL/Przzz8NGdCn15iPR42sztjeIwEJSEACEpCABCQgAQlIQAISkIAEJCABCczkBF7pO/zzm+5/4vnKlkEKnf6jx/8ZdYvnnsmXOtNNn/ohpObq8/HYSbl1I0694Mobche00x77HtRt0Mff5rbFIV7dxc89zzzz0t8hx516drF9NGnesvU88847X7Hty9WuwfIrrMRc9zv82JMr6xOBjvoW5RpzWvv5z6yzzkpEyDV3PvTUtPY1I+8vda+Sdu6p13q/l7tXB3z6419RUmehGbkWx5aABCQgAQlIQAISqH8EZqt/S3bFEpCABCQgAQlIoHYSWDjS0PwVR2Wz6/T4Q/f1792z+++Tfvutdq6gbs7qP3FQP6TNVtvt+PGHw99//slHH/j6y88/DR1g/oUXXWzx117s9HR25QcedeLpJ5176TVEUtx7yzWXfTxi+LDZ5ph9joXiAY98f+jg6lL6fdKk3yZP/vPP/8zyn/8U28fwoUOqLZAUO0a+duxlzle1n68+//TjebN/WsYp570rrNR4tTnmnGuu94cM7FfOfqdnX6Xu1dbrbrjJnY916hpb6j8dOzx476B+vXvGFvtzwYUWWWTixF9++fmnCT9Oz/k7lgQkIAEJSEACEpCABCQgAQlIQAISkIAEJFBLCLw24MOvHn6+W+9aMh2nkRA47PjTz+Xt8/OvvuUeHMJVgaH49cDPJvz9yAtv9lkwvPblhvhw5zfevfmBp14oR79LLr1sA0SYcvSV28fyK67cGGYnnHXRlTXRf030uV27PfZhzmutv/GmNdH/9OizlL0a2c0WeX3QR9+8MfiT74jEmR7zcwwJSEACEpCABCQgAQlIQAISkIAEJCABCUhgJiFwV4fnX+s18ptfCjnFZ5Ll1IlpLrVMg4akgbr7iRe6FYoG4LlR6JpUUERe1AQAiq8PGPPD5NVbtl57Wvs/7cKrbnxr2Gfjp7WffPfPPvscc1Dw+/ZHOnapif5ros9TLrjietIgVVXMvCbGLVefpexVxjz78utvR1xbe4NNNivXHOxHAhKQgAQkIAEJSEACEpCABCQgAQlIQAISqCMEqE3AG968pV9HljTTL+Osy667rd/o7/9osFyjFQstZsu27Xbn+bXdba/9C7Wt7nVEkYeee70X0TirrLZ68+r2w32Hn3jm+cx3oSR907T0le/eOx57risCHGmWyt13TfTX/pkub3V8o98HNdH39OizlL26eFSN7/vJuN8vvO729tNjbo4hAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJzGQEVl61aTMcyLz5PpNNvU5OlyLXPYd/9dOF1952XzELJArjubcGjqR4czHtq9uG6A0iOd4d9e1E9sq2O+++96qrt2hVan/t9jrgUPbbsg2XX6HUe4tpv9dBRxxH/5tu3XbnYtqX2mbW2WabbbNtdmhHZEGp9+a2RwjiWV9yw10PTmtfM+L+UvcqYlX/0eP/rKlnPyMYOKYEJCABCUhAAhKQgAQkIAEJSEACEpCABCRQZgI4ol/u/f6YMndbZ7tbbImlll5kscWXqIkFbr/LnvvicG/SvNWahfqnHgTpdfY/4vhTC7WdluuIIW13/e9+z7896EPmlrXzrrr57lL63ufQo0/kft62L+W+YtsuutgSS5K+6tIb736o2HvSdqs0adai0D2X3XzvI8z/2rsenqLoeaH78l1PxcI99j/s6OrcX8w9c8099zzLrbDSKsW0LbVNKXuVvjv3GDyqXLVQSp2r7SUgAQlIQAISkIAEJFAVgSqLBopOAhKQgAQkIAEJSGD6Eni501OPLd2g4fIzc+Hf6UWMmhL3P/vK27zJXxNj8vb+mI8+HDF86OABhfpPowh4foXaVvc6kQSPRjHvS0IAGDV82HtnH3fIPkfvs/PWD9x+w1X9er395nfffP1lKX1v1XaXPVjb2G+//qqU+4pt+/247759t2f31zfbdsddSqkLgSDzxCs9B8022+yzVzVWKlSN/vjDEcXOqbJ2zVuvvR7Xhg3u12da+6rs/jMvufaWmkrBVMpeXalxk9UbNlpx5Zc7PvloTa3VfiUgAQlIQAISkIAEJCABCUhAAhKQgAQkIIE6QIC30qmZcM2dDz1VB5ZTo0toseY66/OG/Rbb7bRruQcikqHHB1/8eOoFV95QTN+8rf54lx4Di2lbnTZNmrds/fqgj74h5RTfq9NHeg9rO/2iq28i+qGmhbHNQ6zgGe15wOHHFDtnal889Vrv9wq1Jw1So5VWWbVQu2KuX3DNrfeSYos0U8W0L7XNHHPMOWfP4V9OQLQo9d5C7Uvdq0QB8ewXWHChhQv17XUJSEACEpCABCQgAQlIQAISkIAEJCABCUignhO46o4HnkC0IN1RPUdR5fKPOOmsC3CGU9Oh3Jyar7HWuvTdZqvtdizUN07ud0Z8/fMpF1xxfaG21blOJMHrA0d9TUHoaVkrTvNtdtp9r2e69RlG/YKd9tj3oOrMp5R7YNO134gvSHVWzH1EVfT5eOyksy+//vZi2perDUwe6Phqz3L1l9tP63U33IT9tNUOu+xR7jFK2auMffsjHbt0eLlHwaihcs/T/iQgAQlIQAISkIAEJFAMAVNCFUPJNhKQgAQkIAEJSGA6Enj64fZ34rjdZe8DD5uOw1Z7qEKpe3gTnqLGxQ6w0CKLLkb0xFLLNliuqntWXrVJs6+++GzMD9+PG1ts38W2W2uDTTaj7fChQwpGTTRtscZa88w773wjhg4u2LbY8bPtiIaYZ9755z/h4D13rM5amd+5V950FxEaV91+/+O/T5r024Htttyg89OPPVid+ZRyz1+TJ0/u2OGhe6kR0XqdDTYudC81HhBWhg0e0Leqtog4jVZuvFqh/tLrc8w511yVtZ1v/gUWXHGV1ZoOHdy/5HRQc0Zhimat1lyHNEtV79Wmzbg+bHD/KtdV7Hqy7UrZqwhIrdZef6MRw2pmr1Zn/t4jAQlIQAISkIAEJCCBLIFZxCEBCUhAAhKQgAQkUPsIdOo+YMRc4Qxtu0GzFf6Oo5QZbrLltjvstu8hRyIS3HLlhWeNGvH+VG+3U//hkhvuevDJh+65vSrnMLUHfv3ll5/zjU+6n6NOPefiVVZbvfkno0Z8cOz+u273zZdffJbb9oV33vv4tRc7Pc1cuEa9h/8edMSxkZFmkTe6vNDpvluvvTy95+BjTznr2NPOuzRNzdOtS+eO5514+P6TfvttInM+7cKrbiQN0B9//P77GuF4/SuOQX179eD+yeEdHznsvUEP3HHj1fnmu8GmW2676z4HHb78iis3jvIKX995/eUXvjegb2/atlp7vQ3b7rrX/jGlRRln9ZZrrr3kMss2fCPGz/aFYPDw3bdet8cBhx4dNSWWg/EyDZdvRGHu/r17dJ/ww/jv0/bM+d5brrns008++rCU55dtS/Hpp17tNeSmy88/46G7br62lH7ge/ENdz7QZqvtd+K+vu+89Ub7266/om/P7t1K6Wda21KQ/OXew8a80vnZJ8494bD9cvsjQuDIk8++kGdJmiKeRcrynzgmTvz1l4fvuuW6jz8c/n567033P9m5ZYhaW665ytKIIvnmyB46+OiTz9zr4COOW3TxJZcaMWzIoKP3bbf1j+O/H5dtv0GbLba5/dFOr1x+9klHrdasZWuiIHjOV5xz8tEwq2z962+y+dZX3v7A43CmDX9npx2x326fjf54FL/b/Xf/Q7bacdc9//zjjz/Yc1i6n/ibHv/92O/4m5j466+/5I6BgLLvYcechNj0559//vHMI+3vSgWmUvbqTVdccObeBx91/EqrNll99tlnn2PuUNb4O4Al9VnScWH/wjMdHur5xqsvT+vz9n4JSEACEpCABCQgAQlMC4Gi33SblkG8VwISkIAEJCABCUigNAIdOzx4LxEGG2621XbF3kmkw4XX3nYf9RQQLTbafOvtDz/xjPPz3c9b4TvsvvcBVfV92c33PnLPky/lddgedPRJZ1x/72Mdfwtn6xMP3H1rg+VXWAmnc25/OHMbLNdoxfT8CWdddOWN7R9/rnGTZi2XXrbh8gcdc9IZaYQGtRmOP/PCK8KX+t4d111+AQ5m6lPsc+gxJ3J/6DfzNGnRak2c2IgKC4a4gDN76QbLLc+b+Sus1Hg1HNO5cyDH//lX33IPqXDWjNQ848d+9+3qLVuvfcejz3VN025tsuV2O7aIwstLLdtwOc7B/peff5qwWvNWrZuFQ52izE1btF5r8aWWWZbf62606ZbLLtdoBcZbboWVG4dP+Q8c82lbPplToeiTQs92x3hGCEbPPNr+rkJts9cRdR6JAt2sE0Hou2+++rJZq7XWiexZS5bSTznafvv1l1/0fPO1Llu23Xl3nllun6uu3qLVvBHmAMMo4bLU5Ml//knkAntq+VhHoxVXWTW29hQFuCkUTiRO6GkL5JsjURq3PvTMS8ecft6lETjRi7+nECPWOCDqN+S2J5qHc8eEUBZ7crnnnni4PXvggvhbYp/l65+9eOlNdz+EWHL3jVde/GbXF59DuDvrsutvS9vTb2gms/8Z4triSy69zE8//jCe/UXBa6JDGiy3wr9/F9kxiKx68tV3BvP3+WtswkUXX2JJhCf+pmlXyl7lb2Pz7XbcBbGENYVwURHpAV9EOfY1hqAxT6iT5Xje9iEBCUhAAhKQgAQkIAEJSEACEpCABCQgAQnUMQI4Y6kzgChQzNJwjPPWOXny73688+u8mX/mpdfd+sbgT7479ozzL8vt49DjTzun+3tjxlWWqom3zOmLYsS59xIhwbVLb7z7ofT+6+559FkiAXLbbrbNDu1oy9vo+x9+3Cl8v+ymex6uSBMVQkK28O8ZF19zM9dx7tIPba6+48EnU0dttm+iK2ib71ruHE4+77Jr07XgaOY6ERGcO+DIE07LbY/wwLWjI3qkGPYv9BzyUftnurxVTNtS27zc+/0xN93/xPOl3Eediy7vfvApAg1CAPdG1qOF2BcDPv3xr2LqcpQyXjFt032w9yFHnVBVe+bY4eW3+xfqk+LVpLiqrB0O/oGfTfh725133zttc9/TL3fv89F3v+Wmh7qrw/Ov8bz3OuiI49K27HvO5RPAaJMWE9+u3R77pPccc9q5lxx+4plTCYREejDuKedffl2hdbGfGffhzm+8m6ZE4++Atd7y4NMvTuteRdCkPk4EW8xRaC5el4AEJCABCUhAAhKQgAQkIAEJSEACEpCABOo4Ad5sxrFZTP79Ox57risFiHE2F8Jy3lU3342jk1oFqYiAUMG5p17r/V7u/fR928PP5k3/gpBASiruJRIjey9z6Tbo42+feKXnoKzTs7JCvmdddt1tOGt5ixsB5twrbryzsrUguNCm0Fq5vs+hR59YlUM57YN0PziuSX+V2y+Fsq+4tf1juefX2bDN5vS9xfY771ZoLghFA8b8MBlxqFDbUq/Dl7lTXLzYe4kIuPepl9589MXufYkyyN5Hei8EkC59PvisXA7ryIrVCEGoqhoRzIG59Bz+5QSiPqpay1vDPhvPHi603gc7vfYOkUT52hGVw/Mjmid7nYiH/XMiLBATeo385heYZdtefst9j9IHwmG+MVLxDeGs0FwbN23ekr4oeF5VW4S6N4eMHsvfK88q25a1vtp/5JfTsle5t/2zr7xdbAH0QuvyugQkIAEJSEACEpCABGqCgCmhaoKqfUpAAhKQgAQkIIE8BHDa3vLAky+Q4ug/sxQuQk3dB+4htVNVQPc84PBjdtv34CNeevaJR8i7T358HLHbtduz4u3vXt1ffyV7P4IG6Y+GV1J4d7t4K52UQh9+MHRIbn2LA4868XQKHpPvnxQ+9MtYK6/WtPmoEcOmEkbWXG+jNqTkIXpi6KD+fa664PTjK1sLKXPoK42wqGrNpDf6+ovPP/1+7LeVvmWPmHB+vClPYe4rzj35mNz+Jv76889p/YHsNVI58XvU8KnXk9tHg+UbrYjAU0zbUv8oItvUMggQuTUXquqHiAKYX3rmCUdQ5yPbltRST0dqqai90XDN9TZsU+p8cttHRq8V7u/YtQdpy/4pUGeFubz1WpcXEMAqe75wJ+Jm6MB+71Y1N54r6cPytePv5bSLrrqJNFT33Hz1pdl+qFfyyD23Xp89t2rT5q2IYHjyoXtvT8/TBwXCqT1SGfsJsVdpX6gwPG1S0W/owL5VruvUC6+4gfWfe/xh++bWjYnMZ9O8V5lLZNlaZVSkXJvWZ+/9EpCABCQgAQlIQAISqCkCChY1RdZ+JSABCUhAAhKQQA6BC6+7vX2zNdZe98i9dtySItWFAPV+q1tX2qyz0aZbVNaWt8bPuPjqCjHgotOOPZT6DrQlVQ0OZb7nFlmmoC+pgvI5LhEM0jf6uzz3dIfsuESH7Hng4cf06Nb1JcZLr+20x74HLRG1HV585vGHs+2jvu98KzVusjqO6FVXb97q4tOPPbSyAsnc16fnm6/zufEW27QtxKb1uhtsMmRAn15Vtdt+lz33xTl/29UXn0sB7Ny2c88z33y//z5pUu755SLf/x9x/otPR39caB7UBqBNtiB0oXuKvZ5Gyswx5xxTREpUdf/u+x1y5KB+vXuOfP+9wfnavRO1JDjfpMUaaxY7j3ztcPLfFimnqLFw6O7btUnFq6r67PXW68l+bpN3P7eO+iLcX+i5rtasxRpEdLw38H8F07NHu70OOJRnfvu1l56X75nnto99tPHfUXC6dzI3rh9+0hnnI0RQML2y9UQx7m78rW28xbZF7NUNNxn33TdfI5xV1h/1Orbavt3unaJ+BsW7p96r88Ze/X2a9ipRG6S4qom9Oi17yXslIAEJSEACEpCABCSQJaBg4X6QgAQkIAEJSEAC04EANSFwoF9yxvGHvz9kYL9ihvzmqy8+J4og6lO3ztcecYFUUJMmTfrtnOMO2YdixbTjjf8jklz6OFWz4gLXm7ZYYy0+Q7CYyjG68577HZxGGCBMZMfdbJu27UgJ9cQDd/2b/miDTbfclrRPLzzd4aF+vd6eIq3OylGEmAgBHMgUPR7z8aiRVa27W5fOHaPO9Y843atqRxqiijoTfXv3rKrdgUefeDr8Xn2x01O57XDeYhN+GP997rXlIrwktIpRRKoUek60pc2Yjz4cUahtqddjauO4Z4EoXF7MvQgcpN6qan9RfJu+5o8HWUyflbU56dxLr+G5nnjwf3fKxzDffYP69OrB+SbNWuXdz0Q1jB839jsiG6qaGyIdIsOwwf375rajDgXz6fr8s08Us75WkdJp9McfjkgjGkg1dtjxp5/75EP33E7EUmV98Lf5bo83X9t82x12oWZIVWOxrkJ79YAjjz81gq7+8/Ddt+Stc4EgOM17NYkcqom9Wgxr20hAAhKQgAQkIAEJSKAYAgoWxVCyjQQkIAEJSEACEphGAkeefNaFvNnctfMzRTlS0+GIxFhuhZUrnOK5x94HH3n8KiEKXHvhGSfGy9ufpNd32+fgIxo2WnFl3jD/8vNPRyMCZO9dadUmq/NG/GehIGTPk2oHZy3nuCc3CmT9Nlts/f247759t2f31xEuTrngiutvfeiZl/q98/YbCDG582NunCOq4sE7brq6EELm+8SDd99GQex1N95sy8rat1p7vQ25Nqjv/xzg+Q76IJLk2Q4P3INzO7cNYgrnPvlw6kgXoiZGjxo5vNB8uU40Bk72NEVQMfcU24bohd8mTvx1+RX+F8VR6IhMRnNRm2KW/5tllsraEjnCtcnxUAr1V9l1Ujrtus9Bh3d++tEHi4lCSfshwoBnnApiuf3zXIkOKTQvBIsPI13XxF9//SXbtvkaa627wiqrNun89P67FjIAACAASURBVGMP5qbDqqxPalB8NPKDYUQDUZD6tAuvuvHuG6+8+KrzTvu3AHdl9z54503XEHWEyFFZG4SGpRs0XH5gFXsV4ZH6Fn3i7+qzEMpy++KZkqItdJWporJK2qsrrFKxjz4pcm8Xeg5el4AEJCABCUhAAhKQQE0QULCoCar2KQEJSEACEpCABDIEVl61aTNSIz3/xCP3lwpmXNRoIP0OYkL2XlK7HHXKuRcPHzpkIA7a9Fpkelrw6FPPuZiaCl998emYj/Kkl2EuX4wZ/XFueqad9tz3oEUWW2wJ0tdQuyJNL5X2TcqeYYMG9D38hDPOi8LNnyKY3H3jVRefcPCeO6bRHdk5sm5+d3/1ped5I72YtT9y963X46g/5JiTz6qsffPW66wXTSbgaK6szUabb1NR96Pby88/m6/NehtvvhXnc6MRiE6hLsWn4dUtZr44jMcU2baY/nLbkB6JtEXF3IsYQM0Fap6wjnz3LBOL4/w3X37xWTF95muzxXY77sp+fC7SF5XaB4IXdRpy71tw4UUWRWQb0u/ddwr12WKNddaLuihTtdts2x134d5XX+g4VURNvj55dtRjmWuueeZ5+vU+Q4kWOmbfdtvcdcOVFxWaA9dJtTawzztv//fAI45F8Mh3DxEvnB/Sv/J1tWy9zvowqWyvItDw34By7FXEu1JEpmI42EYCEpCABCQgAQlIQALlJKBgUU6a9iUBCUhAAhKQgATyEEiL7r7/3qD+pQKKF7jnITXR3+FpzN574FEnnEZKo5uvvODMrLBw9KnnXkyKmjuvv+LCRis1Xi1fpAC1LXKjK3iLm+iKZx594G6cx7kFghFIIhPTim222m7Hw084/bzur77ceZc2a652z01XXZIvgoG5Uoibz6ygUmj9RHY89dC9d1C3Y5UmzVrka0/BcAoo5woq2bYtw8k79tuvv6osDRWFoomKGJJTBwE2OOMLpSVKx8Lp/VmBFEaF1lzV9aiV8MZiSyy1dOr4LtTXqy92fIq38Umbla/teptsViHU9O/do3uhviq7TsFzBKrQi4aU2gf7OV+9C54pfQ2uwrHPdVgQsTA4j7CxbuwZ9s8HRf6drRGpmuiTPf3D9+PG7rrZ2k1J81TKmtrfet0VRBvt/N/9D6lsrxIlUxUrBAnu5Vnn64O9yvke3V55MXu9OnuVKJdi6o2UwsC2EpCABCQgAQlIQAISKCcBBYty0rQvCUhAAhKQgAQkkIfAwvEWN6fHx9vlpQKKGgkr43jP1lPgbe7d9j3kSJz2fXr8r1A1BxEQe0XUA2+Yj/9+7HfUNCAlVO6Yi0eamq9z3rDfbb+Dj0So6PFG15cQL94b2O/d7H2RBagBv8nrv8NGLVY678TD98+mocq3rsZNm7fEgdyr+/+Khxd7dLj/rlsQQdrlcQJTbLlx02Yt89UvyPbfaOXGq40Y9t6gfGMSYUL6oDe7vvhcbpRJmq6oUL0N+sX5TnqkYtoWu/bcdvBGHNj3sGNOKqaPGy4977R927ZZO99b9ERdsG8QK/KlHiqmf9qwn6mnUJlQVVk/FHpfOEIaYjt/kdsGQQZH+sj3h+YtFp62b7nWuhvwPTdiAZGJfTEw6mQUU3uk4u8lESwQ9YhwILKnWAZpu15vdetK6rR8e5U2rGv40EEDqmLFXiW91edjPvkod3zSRe24+94H8Lc2YtiQKfZzKXuVfmlfk3u1VHa2l4AEJCABCUhAAhKQQD4CChbuCwlIQAISkIAEJFDDBCbFK9YMscii/xMuij1IV9M4Km4jTGTv2Xy7nXZFtHjmsfvvTs/zlvclN9714Ldfffn5ZWedeGRaP+Krzz8dk72XnPtEZnz/3bffpOdxJFOku8P9d9y81NLLNuR8rvM06j4vyvkuzz/9eDHphHjDHycwhbvzpYuqigEpqXjTfZMtt90ht92KUaMA5/QH7w0eUFUfiy+x5NL0k69NWtT7mUfa35V7nYgJIjfGRMGAQs+J2iIUFc+t9VHovlKuUyT75U5PPbZV2132oN5CoXt/j7xQlUUY7HfYsSfjtL7p8vPPKNRPVdfZz4hbCGKl9LNe1CXhntz9TB+xz1t8PHL4+4VqTxA5Q3qx3BRjyzRcrhH7Ivb7VAJdZXNE/GC8e2+55jLSURUbxZLb34vPPP4w4hyF4HOv8XdYeK8utfT3kfotX8TQplttvxNRJdO6V5kXe7sm92ope8G2EpCABCQgAQlIQAISqIxASf/IEKMEJCABCUhAAhKQQOkE0rRMaWqXYnvY66AjjuMN65c6Pvlo9p6NN9+mLW+RvxVpmTjPm/NX3/nQk4gNZx138N5ENaRvX4e/e4raEWmu/YkTf/m3YPERJ515/t///P13FMa+ZsXGqzWlz9y34BcIxYLz8RL878XMf7VmLdeg3TtvvtqlmPa5bUj502D5FVZCYMleC8GiYn5VOV4REWaPCtSk4sntd6llGjRst9cBhw7p36dXbk0A2q6w8qpNvo3wk19/+eXnQvOmLW2KLdBdqL/Krt961cXn/BTpqy656e6HQgOqeA6lHhtvsU3bE8666Mr7wjmfb92l9Md6EQciBVOlhdHz9UdxaqIoSFuVe50C6VEKZKqi0rntWq657gbU9cg9Txo0zo2tRKTKbb/QIosuxt8ItVpefbHTU0QikU6tFA5p2zQ9VZoCLT1PwW1qyhQSCSJoaO7fIsQid2z+rg8/8Yzzib7o9PhD9+VeL2WvktINUbOm92p1+HmPBCQgAQlIQAISkIAEsgQULNwPEpCABCQgAQlIoIYJ9O319hs4wfc6+KjjSf9SzHCrrt6i1YFHn3QGRbVzc9c3bdl6LVL6hC7xA875sy+97rb1N9l86+svPefU9O31eNu7IlKC4tTZ8eYM7yi/f5806Tc+ERb2PfSYk24LpzgpcciLT20H3tTP3jcxLvIb52px82/einb9evV4s1B7nKm8/Z1tN0u8iZ+U7piidkdaNJo30tP2rIGixOlv3lSnJgERKrljn3L+5deTyumWKy/MW9SbCI5ia1KsuErjJjjgqQtQaI3Tcp1IkYtOO+YQns09T774Bs72YvsjomH/w4875cb7Hn+uy3NPdyi2oHRV/RPxwbM5+bzLroVlMXPZff9DjyJl2dMPt7+TwuC591CXIvtMifohaiHbjlRlqzVv2TpfhAZ/B7SdO898qOnBHsv2ldbMGPBuz7dIC3bzFRecyd9QGn2TbUsaMiIwODdHCGFpTZq0DXuV79HNn9n7iPrgd3ZdRB7lRmJE9rZv8+3V3SN9F/8dePDOm67hbz2XWWl79X/iWrG1WYp5praRgAQkIAEJSEACEpCABCQgAQlIQAISkIAEZlICG7TZYpsBY36Y/Pqgj75Ze4NNNqtqGau3bL12t0Eff9tr5De/4LDMbdtz+JcTHuj4ak+ctOdffcs9gz7/6Z9zr7jxzmy7G9s//hznSf+UPc8b+pzfbd+Dj+D7828P+rDDy2/3Tx2+dz/e+fWnXu01VTFlnL7cd/Cxp0zh6MeJfsbF19ycGz1yw30dOr0+cFTelEy567n+3sc6vjlk9L8CAylwXuk7/PP7O3btkdv2yJPPvpB5pA7otrv+d7+Bn034e6PNt94+2/b2Rzp2eWPwJ99lHeo777nfwdx73lU3/5tKK7d/uMO0mG129R0PPgm/YtqWo80OUcuAPdS134gvtth+592q6pPnyZ57+PluveFz4jmXXF1qCqeq+j/m9PMuhSX9U4y9qrZwZ94d3+j3AUJEblvmxfVzr7ypIkUXbdiTj77YvW+2bau119uQMfOlbmI/cO2+p1/unr0HkeTdUd9OPOS4U8/Onj/61HMupv26kaYqPX/5Lfc92n/0+D+32Wn3vbJt2XPvjPi6QrDb+5CjToDnOhu22ZzfCBi3Pfzsy/yt5q5tzfU2asMYaX+kh3pr2GfjTzr30muy/R98zMln0q5pizXWSs/TljGfeq33e4yRj28pe3WP/Q87mjGouVKOvWgfEpCABCQgAQlIQAISkIAEJCABCUhAAhKQwExOAKc+jnkch7wp/98Djzi2ReTkJ/URggBO94uuv+N+nLc4K/PVcABBpzf7D8ex+kLPIR/RF+IA6WOmcIKGsMC1Wx965qWswxNHdvehn37/ZNd3BuNsx9FKEer0XuaVTyjgeoeXewzo/t6Ycdu122OfzbbZoR1z7fvJuN/pL/dt+Bd7Df3kunsefbaYR7bjHvscyFxxaLOWt9///IfeH377az7H9LY77743ba+87f4Op1141Y2wuuXBp19MBZd0vC3bttuddjiT4YiDfcCnP/7V/pkub+WmmUrvIWVOPlGmsjXA8PZHO71SzBrL1YY91OXdDz5lnp26Dxhx3BkXXM7zwIFO2ifEAcSrdG/QJmpHbFWu8bP9HHb86ef2G/39H+yBq26//3HEI6JdiCLA4b79LnvuiwDGXF94572PqxI2nntr4EjEvEOPP+2cJ17pOYg+c2t2EP1AX/zdINrkpsfiWXD9rMuuuw2xhr4QK+gXESw795vuf7IzeydNkcY1IjjYS/SBGLX5tjvu0na3vfbvOfyrnx7v0mMgbYi04G+Pv+Nr7nzoKfY57Ul3lcsYcQBx4+HOb7x7xElnXYCA9nLv98ek6avS9swNjp17DB619Y677rnL3gcext8Zgh//bcj37Erdq6dfdPVNfT767rfcv5Oa2Bf2KQEJSEACEpCABCQgAQlIQAISkIAEJCABCcwkBHA0HnXK2RfhuMTRmWs4WHGEErlQ2ZJwpPJ2NQ7QE86++CrqCeS2JbKAKAOclLnpZriHcXt88MWPOHaz96ZvmeeL7OBtdQSOdM44cs+89Lpbc9PtENWBoxZxoZjHghP1zEuuvYV7cNzi5E6Lhufez1of7PTaO8yB9jjK86Ulos/Lbr73kXSuiBUXXHPrvZWJFYzTfI211qU9YkehedM/ogrO8UJty32d9RIxwNv3+fYQjniEJ/jnClnlngt1IIhIYS/lmwt7NNJwXZcVBvLNgYiRPh+PnUQfrw348Kt89V422HTLbbmOYHDKBVdcn9sPacUQMrLzIAIkreeSbY+Q89hLb/XL7QPRgmgU/m7SfvhbTeuV0J5Il/TvgGikqvYLa0/7QfCrTIAgZRbPLW3b/tlX3iZNVmXPq5S9Sh/8t+CZbn2Glfv5258EJCABCUhAAhKQgAQkIAEJSEACEpCABCRQRwggSvBWPG9xb7XDLnvwRnkhx26pS6dod+49pOBBkMiXnoc5EOWw6GJLLJlvrAUXXmRRHMet19lg42zdiGxbRIVd9zno8FLf5kboKHb9iDC56a7yzRfhA8ZVOX/T+9I3+CsTS7L9pymy9jr4yONLfSblbL/Usg2WI8UY4gQRDXyn0HM5xyimL4SRVZo0a4GYRsTMplu33ZkUR6UIJtSKQPyqKnXVWutvvGlVaY3Yk4zN31STqHdR2dzpp6p6MvxtrLPRpluw1/OJXAgb/C0Uw4bnUUzdEWpbsFdzo5XyjVHKXuV+ojWKjXgqZk22kYAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQggRokQA0FIjFwnBcahroEvA1PoeZCbb0ugXITKGWvpvU9jj/zwivKPQ/7k4AEJCABCUhAAhKQQLkJ/KfcHdqfBCQgAQlIQAISkIAEZkYCTZq3av35mE8++uP3SZMKzT99e3/UiA+GFmrrdQmUm0D19ur77tVyPwj7k4AEJCABCUhAAhIoOwEFi7IjtUMJSEACEpCABCQggZmNAFl7mjRr2frDD4YOKWbu62y46RY/fD9u7Ljvvvm6mPa2kUC5CJS8VyO1FWN/+MGwovZ2ueZpPxKQgAQkIAEJSEACEqgOAQWL6lDzHglIQAISkIAEJCCBOkVg3Y0325J6C4P69e5ZaGELL7rY4qs1a7FGMW0L9eV1CZRKoJS9St8btNlimwk/jP9+9Ecjh5c6lu0lIAEJSEACEpCABCQwvQkoWExv4o4nAQlIQAISkIAEJFDrCGyyxbY7MKm+Pd/qVmhyG2++TVsKihfTtlBfXpdAqQRK2avLNlx+hZUaN1m9X6+33/wnjlLHsr0EJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlMRwJETPT56Lvfnntr4Mhihu3wco8BFOdeYqllli2mvW0kUC4Cpe7VUy644nqKw2+78+57l2sO9iMBCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAI1ROCIk866AKfuQUefdEahIVqvu+EmtL3t4WdfLtTW6xIoN4FS9uq88803f8/hX07oPvTT7+eYc665yj0X+5OABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIIEyElh08SWXemvYZ+Pffv/zH6Lu9sJVdf2fOB7s9No7CBZrrb/xpmWchl1JoCCBUvYqnZ1w1kVXslePOuXsiwp2bgMJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKYcQRmm2322e9+vPPrOHX3O/zYkwvN5OhTz7mYtjfd/8Tzhdp6XQLlJFDqXl1v48226j96/J+v9B3+OZEW5ZyLfUlAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkEARBBAV7u/YtUejlRuvVlVznLiPvPBmXwSIJ17pOYjoicraU2A7TcXzav+RXy62xFJLFzEVm0igSgKl7NW7EmGtc4/Bo0Jnm72qjjfZctsd3hnx9c8IFuts2GZzH4MEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQnMAAIUFx4w5ofJfT4eO+nEcy65utFKq6yanQaFsvc66IjjuvYb8QViRb9w6vJ57V0PP91izXXW5032tD2ixpZt2+3+6IvdK4SNboM+/naVJs1a1MSyov//S2y2+Fwg87smhrPPWkCg1L3aa+TXv7APKfreZqvtd8pGTsw622yzrbneRm2uuuOBJwZ+NuFvxIrtd9lz31qwTKcgAQlIQAISkIAEJCCBkgjMUlJrG0tAAhKQgAQkIAEJSKCWE2jWas11TrngiuvXWHv9jZjqH79PmvTzzz9NmGee+eabe5555uXcpN9+m9ih/R03P9vhwXuOOfXcS7Zrt8c+/5l11lknT/7zz58nTPiRt9jnj6IWtP0njje6dO541fmnHz/uu2++ronlI1DEgVjSNGzxsEFh33NyjYYL1MSQ9lkLCJSyVx+448ar9z3s2JP2P+L4UxEr/o7jl9jXf02ePHnBhRdZNI0SGj50yMArzjnp6GGDB/StBUt0ChKQgAQkIAEJSEACEiiJgIJFSbhsLAEJSEACEpCABCQwsxBo0rxl640222b7lVZr0mz+BRZaaNJvEyeG3vDlsMH9+779WpcXwtf7Y7qWpZZp0HDTbdq2a9p8jTUXWWzxJcIHPPmH8ePGjhw2ZFCPbl1f+vLzT0fX5LpDsOD/yxEqGoehULwX9gVjKljUJPna0Xcpe3Xe+eZfoM1W2+3Yau31Nlxy6QYNESpiK//wyagRH/Tt2b3b0EH9+9SOVTkLCUhAAhKQgAQkIAEJlE5AwaJ0Zt4hAQlIQAISkIAEJCCBshIIwYLIj0XDlko6RrCYpGBRVsx2JgEJSEACEpCABCQgAQnUcgKVFhes5fN2ehKQgAQkIAEJSEACEqgTBJLoCsQK6mMsEjY2FSvqxAJdhAQkIAEJSEACEpCABCQggSIJKFgUCcpmEpCABCQgAQlIQAISqCECcyRCxfLx+U/YV+k4poOqIeJ2KwEJSEACEpCABCQgAQnUSgKz1cpZOSkJSEACEpCABCQgAQnUcQJJoe1ZY5nNw1YM+ytsSNjvdXzpLk8CEpCABCQgAQlIQAISkEBeAgoWbgwJSEACEpCABCQgAQlMZwKJWEE9uYZhrcL+CJsYNj6ditEV0/mhOJwEJCABCUhAAhKQgAQkMMMJKFjM8EfgBCQgAQlIQAISkIAE6imBOWPdbcLGhc0eRioohAsPCUhAAhKQgAQkIAEJSEAC9ZKANSzq5WN30RKQgAQkIAEJSEACM4pAEl3B8IuFEWWxQFiDsFHpnIyumFFPx3ElIAEJSEACEpCABCQggRlJwAiLGUnfsSUgAQlIQAISkIAE6iuBVKhYJgBQu6J72Nj6CsN1S0ACEpCABCQgAQlIQAISgIARFu4DCUhAAhKQgAQkIAEJTH8CpIBaLmy+sB/CRob9wzSMrpj+D8MRJSABCUhAAhKQgAQkIIHaQUDBonY8B2chAQlIQAISkIAEJFB/CBBdsVTYWmHzh40O+7n+LN+VSkACEpCABCQgAQlIQAISyE9AwcKdIQEJSEACEpCABCQggelEIKlfwf+Dk5r1y7C5w8aH/T2dpuAwEpCABCQgAQlIQAISkIAEai0BBYta+2icmAQkIAEJSEACEpBAHSUwV6xru0S0+Ck+f03XaTqoOvrEXZYEJCABCUhAAhKQgAQkUBQBi24XhclGEpCABCQgAQlIQAISKBuBeaOntcN+CSM91I8hVFTUr/CQgAQkIAEJSEACEpCABCRQnwkYYVGfn75rl4AEJCABCUhAAhKYEQSoW7Fo2AJh1K5AuPCQgAQkIAEJSEACEpCABCRQ7wkYYVHvt4AAJCABCUhAAhKQgASmIwEiKhYL+y2MYttfhf0+Hcd3KAlIQAISkIAEJCABCUhAArWWgBEWtfbRODEJSEACEpCABCQggbpEICm4zZJICTU2bNawH8P+qkvrdC0SkIAEJCABCUhAAhKQgASqS0DBorrkvE8CEpCABCQgAQlIQAKlEyDCYr7MbaPiu/UrSufoHRKQgAQkIAEJSEACEpBAHSSgYFEHH6pLkoAEJCABCUhAAhKotQSIqlg+bOOwZmGTLLhda5+VE5OABCQgAQlIQAISkIAEpjMBBYvpDNzhJCABCUhAAhKQgATqNYE5E6GCWnKkhbLgdr3eDi5eAhKQgAQkIAEJSEACEsgSULBwP0hAAhKQgAQkIAEJSGD6EZg7hqLoNsLF7GHjpt/QjiQBCUhAAhKQgAQkIAEJSKB2E1CwqN3Px9lJQAISkIAEJCABCdQtAhTYXiiMuhXfhP1dt5bnaiQgAQlIQAISkIAEJCABCVSfgIJF9dl5pwQkIAEJSEACEpCABEolME/csHjY12ETwuYotQPbS0ACEpCABCQgAQlIQAISqKsEFCzq6pN1XRKQgAQkIAEJSEACtZHAHzGpMWHLhrVQsKiNj8g5SUACEpCABCQgAQlIQAIzioCCxYwi77gSkIAEJCABCUhAAvWRwA+x6AFhs4S9HzapPkJwzRKQgAQkIAEJSEACEpCABPIRULBwX0hAAhKQgAQkIAEJSGD6ESAF1J9h84ftnHxOv9EdSQISkIAEJCABCUhAAhKQQC0moGBRix+OU5OABCQgAQlIQAISqHMEKLI9exjCxVphS9a5FbogCUhAAhKQgAQkIAEJSEAC1SQwWzXv8zYJSEACEpCABCQgAQlIoHQCRFcsH/ZN2MdhvkBUOkPvkIAEJCABCUhAAhKQgATqKAH/gVRHH6zLkoAEJCABCUhAAhKolQSIsPg2jKLbrcJWG/T5T9Sz8JCABCQgAQlIQAISkIAEJFDvCShY1PstIAAJSEACEpCABCQggelIAMHi7rCeyZhN43PW6Ti+Q0lAAhKQgAQkIAEJSEACEqi1BBQsau2jcWISkIAEJCABCUhAAnWUwJeZdR0T3xeoo+t0WRKQgAQkIAEJSEACEpCABEoioGBREi4bS0ACEpCABCQgAQlIoHoE1mj4ry5BlMWPSS8U4J6nej16lwQkIAEJSEACEpCABCQggbpFQMGibj1PVyMBCUhAAhKQgAQkUPsJIFh0T6Y5X3xuGXUsZg37P8xDAhKQgAQkIAEJSEACEpBAfSWgYFFfn7zrloAEJCABCUhAAhKYUQT+iYGHZAY/Lb7POaMm47gSkIAEJCABCUhAAhKQgARqCwEFi9ryJJyHBCQgAQlIQAISkEB9IjAsFotxrB62ULp4oyzq0zZwrRKQgAQkIAEJSEACEpBAloCChftBAhKQgAQkIAEJSEAC05/ArzFkh8yw+8b32ab/NBxRAhKQgAQkIAEJSEACEpBA7SGgYFF7noUzkYAEJCABCUhAAhKo4wRyCm+/Fsv9PlnyYfG5eB1fvsuTgAQkIAEJSEACEpCABCRQJQEFCzeIBCQgAQlIQAISkIAEpj8B6liMDJuQDN04PtdIp2FaqOn/QBxRAhKQgAQkIAEJSEACEpjxBGaZ8VNwBhKQgAQkIAEJSEACEqhfBBJBgpeHLgy7IFn9B/G5btgv/M5EY8xwOMl8+bcDQgsH3//9HXP9J9rMwicXs9+LmXyOQJM7Dn2m/25Jr/07j3TMYsaxjQQkIAEJSEACEpCABCRQuwkoWNTu5+PsJCABCUhAAhKQgATqIIGMg36lWN5LYasmyyTSYlS65NogWsRc06js2WNec4b9Gcb3+cOoxTExjH9XcA1DTPgrufZ3fHI/vznPd85xpN+5d9bkPOfmTX5z/vfEuHee5NrPmTlwnflwpP0mP//3URsYTjEhf0hAAhKQgAQkIAEJSEAClRKwsJ+bQwISkIAEJCABCUhAAjOOwGcx9HVh9yZTOCs+jwjDwT/djkwEBf8+wFJxAtEAQeCPsJXDVgxDVCAKZMEwokLGha0QhtCwUNgcYcPDfghbIPlNrY60X9pzULODfieHLZp8/yk+Fw5rkvz+MT4RRUaHLRbWNIw0WvOFIVB8EvZRMgZzRthIRQz6xdJojGRYPyQgAQlIQAISkIAEJCCB2krACIva+mSclwQkIAEJSEACEpBAvSAQYsFmsdA3MotdLr5/nv6uyQgBUjfFOAgMRDggOCwZNj75RDRAiEB4QCRYKwxBAoHgy7CNwogOaRa2ZtjgpE3r+Hwi7P2w7cMQHbi/Udg3yf0sDwFkqbAxYYgf9P1yd27p6QAAIABJREFU2Ophe4UNDOsf1ipsQNiwsLZhPcOWTe6nb9pwP0IHwgZiybdhiySfCB4IQH+YPgrsHhKQgAQkIAEJSEACEqi9BBQsau+zcWYSkIAEJCABCUhAAvWAQIgGpDq6JGyfsKXDDgt7IKwixVFNCBZJmiciHnD0MyYREEQ5bJ583zQ+ESGIaiDqAfs4jHRMGCIF9Ta6hyEerJPcx78vEAp+C3s7bBvWEAeRDpVFd2evdY12m4TNHYZwQnQE8+obhkiyaVifMMQLUlJhpNUikgMjegNxo3tyH0JQurav4zvCyeRgmjd9VDJXPyQgAQlIQAISkIAEJCCBGURAwWIGgXdYCUhAAhKQgAQkIAEJQCCJctg1vj6TEMFJT7QBIkHZBItknLTWBJENiAKNwhAfqEOB6EA0Aw5+hAqEB9I/fZXMiznxmygM7uVAmEAEoD8OIhu4Xo4j2xeRGYgr2XG5jvBAlAXHMslvhA6EC4QOoj4QOxCFEDnGJHOmP1JH/WPURTkelX1IQAISkIAEJCABCUigPASsYVEejvYiAQlIQAISkIAEJCCBahHAYR5iwltxM6mXSGuEqEBaKBzs03wk0RTUd0BwwOlPVMIqYTjscfi3CGsYRkooRABECMQK2lJEm3RKzG35MFJHUb9ibBg1KOYKQ+BID/ou15HtiygMxuJg7FRsYW6ILXBDZGFNiBVEgXAPNS+YNym2RoZR3Jw1UdicNhOCD4LHn0ZdlOux2Y8EJCABCUhAAhKQgASqT0DBovrsvFMCEpCABCQgAQlIQALlIkCUwoVht4Tx9j9pkT4Moyh1SUciUHAPtSmILCBlE/UnVkt+E8HBOYQJhAhSO30XhmBBBAXjklaJOTUOQ6SgODhRFPz7AWc/52iLEILoQVsEDsYr15H2Rd+MgcBAAXDEB4QKRBdECeaGWIFwwtypscG9DcIQNhAxWGMqCHGO9FIIQ4gdI8L6BzfO8buCuQJGuR6j/UhAAhKQgAQkIAEJSKB4AqaEKp6VLSUgAQlIQAISkIAEJFAjBMJZTr840p8Nw/GP4/zEMApIIzDkO/h/+fT/5/nk/vQc0QjNw6jvQPFsUj3h3KdvnP/0j2iBM59UShSmni+M+3DY9w4bGrZDcs9z8UmqJQpqE8EwKYyaEQgFfE/FBPpYMQwhg3MIJXzPHmmBceplZA/ECOpT0AeCxJgwojm4n2gL5sbYwOI7Y1OYm2iQdmEIGy+Gse71wxBsmBt9IMaQ2oroCoQJBA0EF+5BhCF1FKyp08G6uQ/uGMJO+gzSc3Hqf0dN1Bj5t3O/SEACEpCABCQgAQlIoJ4RMMKinj1wlysBCUhAAhKQgAQkUGsJ4CR/OezsMCIYTgk7Jiw3yiKNbECgoE4DTvS0EHaj+I4IQRuc+AgYOP9Ji4RQwT20fz/5pD3naUeEAo59xAt+U6T6lTCEgTfDOBiHefYPw/lPyiWEgZXDcPrznZRN9Ik4grOflEv8u4N+uadH0hcRD6wtFUkQJeiX/hEhiJagnzXC+iVtP4hP1ocQwn2fJH1xL2IGcybFFXNI10I7xm8UhmiBMEL0RVogHFa0Jw0XbBBnGJe5jglLC3ynjFgTfVi4O4HvhwQkIAEJSEACEpCABMpFwAiLcpG0HwlIQAISkIAEJCABCUwjgYi0QAAYEpa+WLRZfMfBjyMdEYPzONIRHvhcIYwICYQEoim2D8NBj3CASPFF0o6oB9rgmE+jK+iDqItUUEhTLxHBgOO/UzIuwkLq6EdIoBYGv1MhZIn43iiMVEyMwXf+nYHQQRvGRGTgOo7+7MGaSDXFJ/cipHAP96YRGqSlGhNG2qpPk7asmXkT9UEEBr/T+h+7xPelw4gAQYxAOGGdzBt+CA5plAV1OBA7ED6YI0IGYyCkpAISURe0Yc2jk3b0QXv6Zb4W7w4IHhKQgAQkIAEJSEACEphWAgoW00rQ+yUgAQlIQAISkIAEJFAmAiFYIDQ8FbZz0iVO8UZhvM2PEVGBMx/HOuIGYgGiBSIDzvgdw3D0c+DAp4g2/89PCiSc7TjvERCWDCP1EumPMMZFsOgbhoCAw/6lMJzxREbgmKcNxjkEhvRgTkQzMFf6RBDhOuIGjv1UtEgLeiMiZFMrIThwP20Zh3Wm9TcQHhBmmEO2uHc6B+aJsXb6YNy2yf3UAlknjDXThlRRGCmimAtiBWuGH3NmTnBBoOFApHghmRPiB/wQTYjyQAgiooM5sR7EjV8jPRTz8pCABCQgAQlIQAISkIAEqklAwaKa4LxNAhKQgAQkIAEJSEACNUEgRAtSIFGbIT2ujS8PhuEMxwF/eBiOfIQFoiQoGo0IQa0KHO4cOOBx9BOBgPH//QgCiAhECpC+iagEojneSc4jCpB6CQd8mhIKJz4CAp/ZfzukogPX+J4eiAYYDvxUeOAzjUZAOKioB5Gt/ZDU8OB0tiZHOibn0nmkc8umY0rbpddgk7ZfO5kPDDYMa5msn5oerJ/zaZos2GDMNS34jbBBbQvEDYqWwxAhhAiUe8MQeJgfa0Y0oj3s/4r1VVZ7hHV6SEACEpCABCQgAQlIQAJ5CChYuC0kIAEJSEACEpCABCQwgwmEw57/L8fhTjonohQuDjsymRZOcOpa7BVGtMC6yXlSFeF0x1FORAIRFRxEKfDmP+mXcL4jSuCIJ0UUwgaFrQeFEUFAhEFaU4K2pFni8+9wuOet0ZARFxhrllzHPGtJzyXrQpyo0nmf22eyjqmEjeR8lR/RFxwxBBvSQPHJsXEY/IhAQRSCI0IEKaAQLhAzaEvEB1EjaVqutNYGURaIPaTe4oAj/BAueH6rho0Jo+bF52GINhXCTaH1J/35IQEJSEACEpCABCQggXpPQMGi3m8BAUhAAhKQgAQkIAEJ1DSBHId8drhUqEhrU5DmafUwoh3uC+PNfY6uYTi/ESkoxs2BuIBDnsgLogAahZHuKI2IwLmOdQnDCb9sGOIE0QGIGggTtCfNUZqiKZuqKRmm0mgIrldEWkyrQ74SPhWRFdlIjH8nlPOlivvpIzXSZyEGIUrAm0gMRAzqWRD5Qf0PBCAsfS60HxNG9ArpplLmzOCGMNJJkSoKsYM6IdeHUauDlF3U40iLhKeprqYSbopZX2Xr9rwEJCABCUhAAhKQgATqGoH0raG6ti7XIwEJSEACEpCABCQggdpMIHWiIyQQGdEwDOd/s7A9w0jT9GbYDskitolPIi1IR5QeiBGkKEprQxA5wJv9fFJjAWECgQOnOREYb4V9ltxTUSg6sYIREFmQOQ72v9MoimmBXYnTvuiUSlXcX9FHMkd4pNwRHyi0PSYsrUGBqLBKGEIGggMRKDwXeFLnI61vgUjEgZhEyilEC1JI0X65MKIzNgqjFkmamornQqQGUS95RaGkTz8kIAEJSEACEpCABCRQrwkYYVGvH7+Ll4AEJCABCUhAAhKYHgRyajTw/+CkfkJEIOoBR3fjsBZhOMA3qWJOCBCkJMK5PiYM0YI3+YkeILKCVE+kKcIZT6oonO1pYWiiKX6qLNXT9OBQm8ZIUkelkRSIFtQE4XmQ+oloCdJHkTqKa0ShEPlC9EWjMF78IpJi5SrW9HZcoybIe2EfJs8ijeYgWqZCuDDCojbtCuciAQlIQAISkIAEJDCjCRhhMaOfgONLQAISkIAEJCABCdQXAqlQgUMcZzh1Jfjkzfv9w7YMQ4hIj/7xhbaIGemBwzt1epPSiTf2SWdEnQqEC4ppt0nO41AnQoAIAGo0jFOs+P8gUxYhXKS1OhB/KJiNcETkyithI8MQKoiagCEC0JgwxCaiXVLBYlR8J40Xz2+tZJQN4hPx6fWwc8PSqA36QVRCUEqFi/8/Mb9JQAISkIAEJCABCUigHhNQsKjHD9+lS0ACEpCABCQgAQnUPIFMQW3+35vIClIJkQaqeRiFsBEYSCHEQY0EnNjUWcApTlFo0jiRaoiDlFG9wkhvhFMdsWJMGM5zvnPvu2GkIOI3TnNSHJFiCoHDI4dApkB4WqycYtqIF7CEISm1iL5AHOKZzB2GkETkBKITKaKIwkAYgjuFzWHNs14sDCGK76TkosA39zEWfZNSq9L6FkzVCAy3rAQkIAEJSEACEpBAfSKgYFGfnrZrlYAEJCABCUhAAhKYbgQSoYKoCuolkPYJ5zbGW/cUe946DEd29sDBzUGNCQQJHOA4zEn5RFvuR+C4NYw39XGqI2DgROc7aZ/GheFc5//1iRCgz9+ntTB2zjzr1M8kZVdaW4JICVJvwRvhgk9SbHHwHTGJqBfSQyEEcQ5RCN6IFzwjnnn2QJDCeEavhlH8nJRRPMM0cmOKuiJ1CrCLkYAEJCABCUhAAhKQQJEEFCyKBGUzCUhAAhKQgAQkIAEJlEgApzXObNIy4azGIT5f2DlhvIGPsECaoGwEBW/dk/IJEYL0Q9w7OuyRsMOT8RE/eKO/Wxhv8+NgxxHOm/p/ZSIGcKIzDtc9iifAc+I5IPoQDZFGxlDHgtRQpJCiGDpFuHlWRMxwjms8N54PkS3UwyAigyN9xjzzdcIQrHheCEyIWj3DEKfS51j8bG0pAQlIQAISkIAEJCCBOkRAwaIOPUyXIgEJSEACEpCABCRQOwgk0RU4svn/7XnCqIvwRdhqYaSDIqUTb9nvHEY9A5zXtL03DAc2NRG4D2GCWhZ8J4piv2SFp8dnhzAEi8nZ2hRJtABiCWPhMKfoNm/xe1RCoJK0SwgXPJfJwRQBA+EHQ5ggBRfPhmfybRiCBOcRHaiDwTPl/mOTPvjNeZ75pmHsgZZhI8IQrQaGEbnBc6O2Bfd6SEACEpCABCQgAQlIoN4RULCod4/cBUtAAhKQgAQkIAEJ1ASBTAooHNlEVrQKoygzb9+vGbZ5GEW2OYh+oC4CDm6c4o+G8WY+9RPSSAzexuc66Yh4W//ZMASIPcNwbF8fhkOc9EW5R5qmiAgN+uENfo/qE+AZYggPREUgKsCWGiP8m4pICxinz653fEd44hkTKYM4wbPkN8+eY6swoi3oE8GC/UKh9AFhRFowXpqmqvoz904JSEACEpCABCQgAQnMRAQULGaih+VUJSABCUhAAhKQgARqJ4FErEAkoIYBb9oTXYFDmogIalEQ7ZB7IGJ0DiP6gSgKHNS8wU8KKPohBRGOa0SKIWFESuDYRrDgoP+uYZuG8YZ/9uDNf6IC0ggN+vFICMTzgguizz8RXYFgVOyRRl0gAvHc+PcUogXPG8GCPUC9EYqnU4S7U/IMEDiobbFTZiBEKIyDiAueGcIVz4p9wPP+MeY6yfojxT4e20lAAhKQgAQkIAEJzOwEeOvHQwISkIAEJCABCUhAAhKoJoHE+Y2jepWwtcKobUD6pwvCVkq65TcOa/7/G8c0x31hpH5CkEgd1LPH935hONQ5eJuf9FETM7UpeFt/cGa6pJE6Ka6TcqjiiDkxh9Zhq4Y9GfZtNm1U5t5p/pqsH8f93yU6//8dO0ljlf6mLzhh1OSgGHXZjhiLZ5Wm26LftAbIFGmYKkkTNdU8ErGK/oicoEYJB+LT2mHUwUgFLAQk9shhSRuELMZE+CAtFAfRMpckv0k1hZDFHkkjLqYav9h5lg2gHUlAAhKQgAQkIAEJSKAGCRhhUYNw7VoCEpCABCQgAQlIoG4TyERWkB6IKAqKa/M2Pc7rVKwAAg5pzj8fxtv3OMnHJJ845PmN4IDDG2GDKAtSCf0cDuk/cehnnPpD4/w2YURXcFCMu2FcPzjafhOf/D/+JmHrhlEXgbGpuVC2IzMXxiI6gCiDueI8UQFfVle4iHsRb0ibhZEia2z0OTb6o3j4NB+Z2iIIBbBBTCCSBYEI/iXXjkiEpF+j70+TOTNvoitggeDE8yYCg4gO0j8RncFvomioYZKKFayPPYPQgeCBuMH9iBWkk0oFjmnmYAcSkIAEJCABCUhAAhKorQQULGrrk3FeEpCABCQgAQlIQAIzAwHerG8a1iSMt+mJCmgWhrM69+CN+ZfCECNIB8Xb9IgYvPHPNRzTOMzTOgkVNQwQB3iLPiMScJ70Q/TVNhlk2/i8J9rslfymdgZz4u39CTWYUghHP+smoqNx2JgwnPfjqxnRgWDB+og0QQQiGgXBhuLinK84piGqgOeTikIIQ8ydfxMhDjF3flfrSISlH+AdhkiB6MJ4PF/48HwXCIMZdSoQNdZLzmXHpG1awJu2CE/c90EYwpaHBCQgAQlIQAISkIAE6iwBBYs6+2hdmAQkIAEJSEACEpBATRHIpIEi5RK1JIioaBFGZAMpnN7NGfur+P1KGA5tnOM9whAriK7gzXvO8wZ9sYWWiQZAnLg17KBkrB3j8+qwa8JwePN2/uNhpKOqOKahdkPOcqb4WZEOKoxaEKQ9qrbTP+kVpzwCDmIQ3Dj4zvmSIyDyTBzOiArMm0gHRAHEBZ7DNM09EYb+Cs48W54zfSO6MCbPmkgXjO88c/YEc1gmM0/mhdhEkXZEjffCiMLgnhFhlaaHyrNWT0lAAhKQgAQkIAEJSGCmIqBgMVM9LicrAQlIQAISkIAEJDAjCSQOf97+XywMUYC0PYgUpGhKC1sTJUB0QHoQ5XBpWOqsph0ObfrBaY0jGqvSGZ8TZUHfCBKnh5HaaO9ksOPik9REvJH/fhhiBSJCejAGb/0vFmtJx+WTKADmhWMdp/2/0QzcWCCigUgF5sB6GBcR58MwogxKPZgr/TAPRBnSTTEfzlUrZVN2AkR9xLoRKxATOBAp4MX8y3YkwgWsGY/nxHoYi/UgaMGJ/fBGGJETl4fBkYO9wx7iWCeM/UX6LyJyEIWI3iGt1FTPqWwLsCMJSEACEpCABCQgAQnMIAIKFjMIvMNKQAISkIAEJCABCcyUBHDsE01B2ic+NwvbOFkJ1zhwfo8JowA39SbeCUO04BNnOW/dIxIgCkwhDOQjkhUL8ggH48IhfmzS53+T+0kh1CsMBzlO8GzRasQKnP84zpdK5sP1NO0Qc0NswJmOIx1nexr1kW969Md13vznICKA/nCuV+fAIU+f/DsFhzziB8yGhZUjuoI5IYqkhc8ZL60twfeyH4l4Qd+Tk9RWMCZa5MswxAv20FNhG4Y1DxsTRj0UjnRPscfg8GZyDzwqirGXfcJ2KAEJSEACEpCABCQggRlIgH8MeEhAAhKQgAQkIAEJSEACVRBIijXjRKdQMvUhsLvDUsd37t03xQmc0rxZ3y+sb9hPyRv+/D849+G4Jh1QWgOCwtIIG0Q64FSnHfZXoRoUMT/6uS2MtFCMhxN+YFj7uHdU7uSSwtykIUoNoWG5ZC7LxmejMNIxvRr2VhhRCJPyzSP6Yi0IIPRFwWmiOj6NttnIjtwpTPE7U5+D88w9jTAgigUeaSRKxX3TUMOi4v7keSLcMA4CC3OdQpiZ1jGyC8xZX/YSe4BoCyIpKLYNS57lSZUAYz8dGfZRYkSxTC60P6qE70UJSEACEpCABCQgAQnUIgIKFrXoYTgVCUhAAhKQgAQkIIHaSSAczjjiG4XxFjyRCbz5nxa4zk6at955E/7EMBz+RCrwFvxvWady9EdNBiIxSE3EJ8WXVwrDWU0RbxzSpHTCec85vqfpgLgHJ/6/kRNJuijexj8lDMc3Kat4C//iuMYc8h4Zxz1iDELFlmEHJPPJ3kMtjOPDEA6mShcV/eD8Z558/hpjlvTmfyUOfZz5FUc1C3hXtuxadT55BggV7An2FsLPzWHU1SCKJ/d4Ik6MDOO5ErUzJvikKa5q1dqcjAQkIAEJSEACEpCABEolYEqoUonZXgISkIAEJCABCUigzhLI4zjnBR8c5zjicdSvHnZgGMJE9qAwMlEIpEYiHRJFoz8LI6XSP4gVOX1n6zHgoG4bRh0K3vhPaxnk44yT+rkwohhwUhNFMTr65k17UiaNCds5+SSyIq2rMVVfST0O/j2Qplri7X3u576WYdnoEebG2okc6Rw2hXAR6yNKpDo1KyrmVUk0Q8F0WfkAzWznkr0B+zSyBpEKzghYpIZaPoyC7unROr6wXx4Ko3j77PEsuSdv6q5yRorMbGydrwQkIAEJSEACEpDAzEdAwWLme2bOWAISkIAEJCABCUigzASqSNmDUDFfGBELB4dRLwIRI7dIMw7l/mGkFkKM+Dzs52xURR7HMU5q0hMhfgwKoy4GURKkB6qsCDRv4B+VZ/mD49yTYRuFITZQ6wBn9lR1GRLnNhEjRFQgljAWb/MjliC2dEvu5176OyIZjzXen/S5Q3y+Hpatj5FnWp4qkgCiEYYIxd6BNXtpbBhpvrJHo+RZsRdJI3ZPchFxrOg0XEXOy2YSkIAEJCABCUhAAhKYrgRMCTVdcTuYBCQgAQlIQAISkEBtJFCJYIEjf/EwnMdEGOyXmftP8Z3aAxxEUiAOIBIQYYEA8UWJNRzSWgZENSAUrBm2dRjCAvUhdkv6TosxF8L4fDRAYKGOxt8xFwo+8//+vIlPHY7twkhrheBARAWOcV5mooZGmqYKQYWxtwk7P8+ACCf3J9EVhebj9SoI5Ow/hKMGYaSD4nmnhd2pMcKR3Xv8fjSMlF1E+fAcETH+PYywcOtJQAISkIAEJCABCcxMBBQsZqan5VwlIAEJSEACEpCABGqEQB7BgnoCFKLeIGzfsDbJwDiDETK+DOseRsQDkRXDw0aHkRaKtE1/lFIIOTN++v/niAdpOirGI00UogYCxhphiA2MhWMbEYKaGURn8JY+0RZ3hhENQZqgNKUVKZ1wdiOErBVGCifaIrAQFUJKIr5/l9zDuNSlSGtJUN/iwbDsQR2P52KtUzjJc9rUm5+IQqU89xRMzv7juSNasLdIB8U+bJI8M/bWpmFEx6R7kW4ojP5YWK8w9uG/NUQULOrN9nOhEpCABCQgAQlIoE4QMCVUnXiMLkICEpCABCQgAQlIoIwEEAAQLHDg88Y6TuP0SFM14TAmBc/DYdRzGBpGdMJEohlKnUvGqZzWk6AmRHpMCoc2hbzTY0h8SUUEHNsIFaSDIhUU8yCtE4JJRbqmJLJin/iKMTfWhOObOht9wigOPkX6qmQgHOI/Jffz7wbe4qd97zCiNDgoAH1htLmxvhd+DgYwmjM+4UZUS3VrcLAH6ANRjL1FBA9764MwBDT2Hkc2bRh7lOfKnmXvcr/puhJQfkhAAhKQgAQkIAEJzDwEFCxmnmflTCUgAQlIQAISkIAEap4ATmDqVVC3gpQ8pIJKHcTZ0XEkjwsjygGRAEEBJ3UqOJR1pjlvyTNG6owmbdNvSdHtwbnjx3lqcJBKaJcw1oYYQ5ooUli9zbyLmDN9wID6CAgp54ZRP6FpssiL43ORGOv0+poeKilgnvKtKIDNuWJFC55vnigfxCXSc/G8iIxpHtY4jL1Hqq7swfNhrxI1UyGchLE/jXzJAeVPCUhAAhKQgAQkIIHaTcCUULX7+Tg7CUhAAhKQgAQkIIHpQCCJIsAxv0QY0QNLhrULo5bE+jlTINXSu2G88f5+GNEJtept9sT5TRTGtmGkf+L/+3F848B+KYzCzv9GgmRFi4RFRQQH64rf1NVoHYajfOUwanoQ1YEIkooWONTXjPYfTYfHVeuGSKIriHZJxQIiHeA7qQhBqOB6MoXSSesF8/XCDsm5kciXAWHPhRE9g3hBeq8/yzGHgpO0gQQkIAEJSEACEpCABMpAwAiLMkC0CwlIQAISkIAEJCCBmZ4ADn0MRzPHDmHHJd9x8o8J4611aj5QJ4DoBCIOiHCobuqfGoGWeVOfGghpJARRIMPCOiVrIUqDfwtQG2OuuAcHNw52GCC+ZNeEeIFowdv+FBonhdRKYdRM2D+MwtCcfy362SI+R+eJ9GCt9D1VBEodqbEAL1IxsUfgB7NyRtvQP3vtizBECH7z7FqFsT8bhSGsYTzH9mHs5XRfl3MuPEsPCUhAAhKQgAQkIAEJ1AiBNPdtjXRupxKQgAQkIAEJSEACEqjtBJKIAopLk1Zn0zCcvrtm5o0TmsgCoipeDCMNVFoHoqTi2tORBY5q6hpQrDlNLYTA8F4Y/wYgGmDFMN7WR3BgfRWpjML+QXDIiA4IM6mTnE/6I1qDCJMLaJ+sq1F8XheGuPHvkfDlHA52hA3GqVNHkvqJtGBwQbBADCrnOmHMc6D2CHuPPcheZE/y7LL1LNi77OFNw9jT8ybPoE4xdzESkIAEJCABCUhAAnWTgBEWdfO5uioJSEACEpCABCQggeIJ4OxtEIbjHmfvOmHUfeD4Ooy0TxSXxjlMW4oh/4STOk/dgeJHLbJlUh+BFEw4wNM6ElNEdeSJUkCAIX0QNSdI5cQaRkW7PzLpr2hDtAR9LRNGmqiJYf9Em3/fyKcuRfzGQU57eJAyC0Y4578P2ybs1WQ5pInaOoy0ROmBQMLcES0WDMOhT1RAycXJM7wRZPi3TEU9j9qQ8ijhRBQKYhBrK/e80mLcPNO0yDt78vWwvcJ43tRdYe+eGdY3YT0iPkeHpdFDmUfjVwlIQAISkIAEJCABCdQuAgoWtet5OBsJSEACEpCABCQggelIIKk9sHgMSSQCdQEoXIxjeFTYKmGDwp4Nw+lPuw/DxhdbTLm6S8lxzCMUrBCGwx9ndRrdwffKjvnjAvchDBAV8UJyb9qeNX6WrAkxhJodOLsRLbiGcJE9cMTjhEewQaigVgJiBWmKaI9ggVDB8UDM/81gRMQBB//mQKjgE7GCWiF8p5+SRYu4B7GCOROxgRP+l0SEmcIhPyNSTSW1TGBSkwcC0/gwRCCKcPP98bDdwniG7F2iLkjbRQopeMHo65hfdXjX5FrsWwISkIAEJCABCUhAAlMQMCWUG0ICEpCABCQgAQlIoN4RwMEdhvN9sTDS51CLYdMEBA5exAoOClYjFOD8r0jHw5v00xEYTmmc0KT24f/dEU5w1i8cxjzzHZznLXtEmDFhvGk/Mo1CSD5xXONYhwERhNtcAAAgAElEQVRFtBmDFFGMg5gwRd+JQIOIgQiBYEJxbeZCHwgFR2UmQgQGxcuzB3OeL4yUUAgNzB/hojpHWpcBx/2iyRoQRIhsqC9HVrhib7JH2asc7N30+W0a39nb7PHF2POmh6ovW8R1SkACEpCABCQggZmTgBEWM+dzc9YSkIAEJCABCUhAAtUkkDhscaDj1MfhjRMeR3rDTJdj4jsRBKTeIZpgeNivM+ANdaIXmCuREjj5cfqTkooDMSPfG/Oc3yls37CulWBKC0MjPryWcCAqg3HyFhFPhA7um+oIpqSWuiSMmhYcreLcR8k9ONcp6p0KFekY0yL8wAWBAjY46xE/KHpNyqw6dxAtkif9GPwQjkjThTj1cljz5Fk2SiCwp4mOYY8jSLGnP4u+JtWGNFp17kG5IAlIQAISkIAEJCCBaSagYDHNCO1AAhKQgAQkIAEJSGAmJMBb6TjmSUtEKp3Nw7LOfxzB14Th/MchPCPECrAyRyIZ0rfmmTdpm35J5pZPsEjvQdzgzXpEi3xCA5ER9Me/CXB+p8b5f2tYFPlsEQrezrQ9Ob53DyMihVofiBS0wRjzx2qMkXafCir0xVz5jUM+r9BS5PxrfbNKUlxNDrbsYfbok2Edws4Ia5QsiAgi9vbgsIcTRvC3nkWtf+JOUAISkIAEJCABCdRPAgoW9fO5u2oJSEACEpCABCRQnwmQLoeURauG8ZZ+0wRG9v+Nyf3fM4z0RqQ9qizqoEY4ZpzTFMDmrXgEFESKpcLSAtyVRSgw15FhiA6sE3Eg3/xJB0UKKPrDif1xGGNRLPrfdSURKWmKIfqcQsygLW/rRzuKO6cHQsnWca5DJsqCWhqILxwILdMiMCCA0FdaiJpnVFmKrMy06uTXVLAZkjzrfTKrTPc0e5yi8og87A3qXpQqStVJeC5KAhKQgAQkIAEJSKB2EVCwqF3Pw9lIQAISkIAEJCABCdQggUw6qOVjmFZhvGmOQz/36BgnEARw4E/lpK/BKebrGmf86DAiJnBOE/XBnPKmZ0o6oN4EDnz+f59i4p3CstEY1MMgldIaYdR/IGUTa/0pjGiFitRKCS/aUnCcdqQXoh3Xcx3enH83GY/bGfcJ5pkIIMwdoaEcB30xB8ZMhY+qeFQ5ZpJuibRSGHP8t69yFO/Ok87p3zocZeif50CUBc8cFuzdg3IWzB4nJRTiFHt+TMzpN9NClWMr2ocEJCABCUhAAhKQQDkJKFiUk6Z9SUACEpCABCQgAQnUdgI4iql1QEQBzumjw7KRAcz/+DBqOyAMVDjuZ6RjN4leQCjAIU1UAfOuNOojeQCIDumxd3y5OAwxIj1YG4IMzmuECHisHIY48W04s7+McXHa0446H42Sa0sm9yB+5AoE9JfW12AcalZwf7WFhMx8K77mOPdxzk9LlEa2e+ZJjRBSKI0LQ7RgPXAuZyRCGgWSRrUQmfLTtBRyT/ZHKkYRMcTeZQ/fmlkgkTRbhN0XxrPmb6A6qb9yH4m/JSABCUhAAhKQgAQkUFYCChZlxWlnEpCABCQgAQlIQAK1lUASLYBjGof/CmGHh+GgJnogPd6JL6RfSgWBf8rwBvw0I0kEE5zSGHMrdLCGbmE4qZcOI7VVVrDgfhzXw8I+DeMNfaIVaEfaKZz2CCQ460kdhRBBhAephYicIP0QdROyggFtGTc9KPhc69M0ZaJuWB/7gmLs7BPSgiFmlSsqBC7sPcZBMEiLnJPqa1qPVFThebA/eA7s5Q2TjjdOPtnz1Gbh2qyxdvZ3OQWZaV2H90tAAhKQgAQkIAEJ1HMCvEHlIQEJSEACEpCABCQggfpAgJd1cBiTDurgMMSK3OODOIHD95OwfAWtZxZORGQgRqTHieGczr6sRPRAmv4JQYP6BhiO9G/C/sgIPERY8OY+/3YgtRD3UhsDx3tWkOA7QkZ6lNPRX5PcmTcRD8wXEQaR4r0wIhAQa8p58AzgDcPPko6XC9bzwJvUUXnSR5UyPnuWvcseZi/nHux59j5/A/wt+AJbKXRtKwEJSEACEpCABCRQ4wQULGocsQNIQAISkIAEJCABCcxoAuEE5v97eaN9pbCdw0h/lD0Gxw8c1dRgoChxGl0wo6de3fFJw9Q+LE0NdQrrTkSINMUVTm2c9DjsiawgIgInPYJFmsaJN/aJviAKhTfx+STCgigEnPxZwYLf22UmjEO+bOmgqgui0H0RYcAaWTcpoVgDtT1IBVZZUfNCXVZ1HR6IBFQ1RwxBIGod1iCMqI5pPXhG7F32MHuZPc3ezh7sff4G+FuYP/nbmNZxvV8CEpCABCQgAQlIQAJlIeAbNWXBaCcSkIAEJCABCUhAArWVQOKkxzlMqqN1wrYO4+3y7MEb9T3DiErAQV+u2ggzEsvwGJw6Buclk3gmPqll8BW/w1E/OdggTryQnMfZ/V2y9jRNEA52CnI3CiO9EJ9pO8SOinYJYwSPdpkFD4jvtV6wSOaLQIGAQ+RIkzBSKiFilDvKhv6oQ4IwglBBnQ8Y/ssyw6+6X1ORib18Q9hGYRSYTw/2Pn8DrLE3647nl7eeRW1Ih1ZdCN4nAQlIQAISkIAEJDBzElCwmDmfm7OWgAQkIAEJSEACEiieQJryB2d9yzAcxbnH23GCN9Fx2OO8LelI3lJPow3+riV1AXCO3xm2X1ijZEHnxVxPjflV1MEguiB+80Y+zmvmnyvU4EwnvdSoMFJAUdcBZ3taBDwVNkgZRYQCUSwc1MMYWhLEGds4TdHEulgf6bKIyqkoul7GAwGHtFPUD4E147HnSLVVbZEMYSEnlRR7mHEYj34PyFkDfwP8LRAFQ7tyCiZlxGVXEpCABCQgAQlIQAL1jYCCRX174q5XAhKQgAQkIAEJ1D8CpNqhbsC6YftXsnyc60QbpDUaiqaUKdqMo5uxJsW5X5NUQ0X3U66GOc5rnNEnhj2f9H90fD4X8+sV7SqKPSdv0SM8VFZ8GVFjTFwnMoN/P5AyCUf75GQshI7GYaQZSo/X48uHtUS4KRYtogXFxjkQK1hXTUSIpPVD4E+0Bb+J6ilX8Wv6oc/xYYgVlQlH/C0gllBQnblUWzApFrDtJCABCUhAAhKQgAQkUIiAgkUhQl6XgAQkIAEJSEACEpgpCFRSrDitXUGxYdJBUash9xiYOGuJSCjpjfpErOBteYoYM1bq9KafGVZ0OpPK55+Y40sxl0PC7k8W3ik+b4/zt8XnF8UIKwgP0Z41pamT/knOseZVws4O2zsD9t74jsN8pjgyvFKnfU077+kfG1+Dog7Pij3NOOzx3Mgi/hb4myC6KBXrplg3f1OmhZoptrCTlIAEJCABCUhAAnWGgIJFnXmULkQCEpCABCQgAQlIIA8BHOoYkQ9tkutj45Pi0RwIDN3CcO6SBqg6NQvSt/CJPCAVDwWVKxz8NeiMLvphxxz+irk8ETdQx+CEMAo9n57YBnGNWhOpY3uqfv8fe+cBH1d1bf07XV2yZLn3ggs2NmB67wEChNAhlAAJCYSPUAMkhPIISSgBktASSgqEEFrovYReDKbYFGODjbstN3Vp2rf+o3vFaDyyiiVb2Pu8tzMzt5yyzjn85L3O3iud/HBvcoLfr/fQQiCt0GWyA9JehCD5Qu91h2h1u8fdkx5ci9O/q6Iqsg2XOWVNs7ZZ4xNlnnaLtwfYE9czn651N1HTk6bF+mIIGAKGgCFgCBgChoAh0AMR4A9TK4aAIWAIGAKGgCFgCBgChsDGiAApfSARxsuOk0EkUDyygu/oVrwl44R5VuHhtQHjEhJEUuAA9qIq0HKgDUiSHlFczQpICvQs0ssb+vFHGWLZw2Q4tOk3B5tSmhycsnejV/i3A9fRqZgiO1p2oyydrEDEmXbm9YiBb9qdgAxhTbO2WeOsda94e4A9wd5gj7BXPB2WTRs5G70hYAgYAoaAIWAIGAKGwAZDwCIsNhj01rAhYAgYAoaAIWAIGAKGQDcjwN+6I2RjZNu7bSE2jWPWK1P1ZbYMTYYWp907kArHe69UdZAeCoc+juIedThI42l0Iy3QtbhUtqsLwmn6xCjvuPalPj91jbGQUmusOybSCJ2XhqH39U/68i/ZrJ4QWZKlfxv1pVbWK5E+rG3WOGt9mzQQvL3A3nhbtlr2icwiYzbqlWKDMwQMAUPAEDAEDAFDoGcjYIRFz54f650hYAgYAoaAIWAIGAKGQOcRCOtVoh1ek/2fW006WYEwNGLUc2Wd1ptwtRwQT54l48Q64tToN3QmvVTW0Wboc0CENKfu6QCxgh4B6aFe1vuctr9W9sOMBiEjsI6Wu1yMV1sqqI5C1+3Ps7ZZ46x19Eb2ztgLkFHskb4y9owRFt0+JdaAIWAIGAKGgCFgCBgChkBrCBhhYWvDEDAEDAFDwBAwBAwBQ+Bbj0AWwW1S25DaCAKhj+uMTR8nug0QFhWyallnoytSdeKkVx/m6yt/X1NXvD1i1h0EnrpJ5YPhVMYJXdvBOuhrSuxZ/T1Vn9fIvis7Szawg3VByKB/8KTsc7DcUJEV7vwz555eSbMmR0cInQ6Ov8Xj6oPXNtcjzJHa7jQRti59yXiX9cgaZ62z5iHxtk57BqICfQsiadgz4Nid2hpdODSryhAwBAwBQ8AQMAQMAUNgY0PACIuNbUZtPIaAIWAIGAKGgCFgCBgCIIDzmPRMpGkikiCzPKQL02Qph3JXONpdIgAdi+4ojGeIbKQMh/Mg2XQZKZxWdaZBt7+fytE+U+/f4mK1iz5rZFfLOI1PJMZQt02c2LT5lGy57DMXw4VEbnSmD134jkdQUSVzzm90RbosymVtfXXJCtYbRpQCaci+1PUFwgYiYIMVNwKI9lnrrHlIiXTCgns3y0jzRf+Z/w09nxsML2vYEDAEDAFDwBAwBAwBQ2DDImCExYbF31o3BAwBQ8AQMAQMAUPAEOgeBPg7t0Q2SZaXpQmc/l/Jlsqa0yt1T1e6pFZvPIwJ7QEIDPQI5sopXr8uTnE3TRQn8LF7ZTj7n5UVy2iX6zi5ierAcMDzDLgl11cEQxso0p8Ct2/0D5IFjIgqWB9RDrRF+6Qco31SgvWToRsyvysIsXVcRcwVQuhgsU+Wutgj7BW0LOi7ERbrCLi9bggYAoaAIWAIGAKGgCHQOQSMsOgcbvaWIWAIGAKGgCFgCBgChkDPRQDndX/Z92UHy3Ai42gPuV0mHdSbMsiKmm5I3dQdyOBwRjx5iQwhcUqObIBswbo2mEY6eOQNqaY6nG5qXfvR3vfTUoAx154xzzje6TeEFOLnAT07bz0QBjj40TEhBRkRFswTqZYGyyBNIJmaSxZNEk+XhM8WUSFdQQixxtUmkROsedY+e8CLsmBvgB17hb7eIyPdmKWFau+CtOcMAUPAEDAEDAFDwBAwBLoMASMsugxKq8gQMAQMAUPAEDAEDAFDoAcggPMa5+tw2QSZ59z3yIp3de1vMlIa4ZDFkZut2ziOKYmucBh3AS44sTkdDxGDSPInsq9lkBjrJe1RF4yhy6pIm5Okm46J+VotIwKFAjakhgKz9aXJ4Dn4ISlI00VfIAkglloQFmlA0G+IDYgW3qHPfHZHlEMqIkbG2r9Txm+idLy9wV5hz7B3IDbos5EWaZNlXw0BQ8AQMAQMAUPAEDAEuh8B7x9i3d+StWAIGAKGgCFgCBgChoAhYAh0PwKelgEnxD1tB06Qe45XHMI4+XFotxZdwaGeMhmO5Bw5xMOuU7z7e7/2Fjj9vljG6f3ZMlL8LJJtcoRFOkyufgYRDl66KgSvScs0S4amSLf/m8eN4KD9he7aYr0R6eGlYWptZukbURmQG8NkpLJCO4T1RxquLituJBEEikd0sRco9JW+U9gz7B1PfLvL2reKDAFDwBAwBAwBQ8AQMAQMgfYgYBEW7UHJnjEEDAFDwBAwBAwBQ8AQ+LYgQDqecbIdZD9xO+2dIOcnDmyc20tbEYrGgYzzeKAMhy4nzXHiLne1IjbkiXMc4KTzgaTA8czf8ogkQ8Bs6sVLZUVUAAQOpAXRFczXetFjcAmBKq0THP6sHdYa87Q2DQ36zZpjLr9w1xoEBoSFl2aq3RorbrSQl14qtSbSI4RcvRLWNHV7AvGQfN4eYc8gps46+0i2QQXDN/VFbeM3BAwBQ8AQMAQMAUNgU0TACItNcdZtzIaAIWAIGAKGgCFgCGycCOB4xVG9rey4Vob4X13H4d+aExvCg5Q+pF1CNBlCAAcvTucGHMLrQQ9hbbODk3mmDKd0KnJA/VkvERZZUmeBd6psYEy8buDYx8HOXEFcMMcbIqUXc8SaSaUcawc2EFGQZPQX8okUUqxjiAsEzzsqGu5perRGrtEOe4C9ALmXWdg7PPO52/aGJOmydM8uGQKGgCFgCBgChoAhYAhszAgYYbExz66NzRAwBAwBQ8AQMAQMgU0LAS+9Dg5bcvFnlk9dJyypglo7tY7zH/0Az/mNA5z0OAUyNBJw5K6XE/vpnc+io0H/2n3yvouXgZd2C1w8HZB4OxzzXdyNb6pL17Tw+tRtjbVRsRtpsda5SRc5FxFEii8iHCAoIMhYX0RmIK7Cv9c6QlgwNynh8VYiiOg9fWMPDJGxJzJJC/YO9XiEyXpf7xtq7qxdQ8AQMAQMAUPAEDAEDIENj4ARFht+DqwHhoAhYAgYAoaAIWAIGAJdgwBOX4gFHKwIb2cWUu5wkp2/gVtzwuLM5VQ75Ad1cdIdJzJ1cxIeHYl2FTmicfp6+gl8pk78Z77cEVHvjCgHjzhIr7v5NHxH6m3XgL55iPaKXVzAGef6CvWtbkOSFh0cQ495XJjVC7s57nqDnIA089ZKZ6JnWBfFqnOVS55kjpW62QPsBfZEJmHBnPIM6591b4RFj1kt1hFDwBAwBAwBQ8AQMAQ2fgS6XYBu44fQRmgIGAKGgCFgCBgChoAh0AMQwElLKp3tZLvJPBHh9K79Tz9ekKFJ0ZpjH0JhpWyZWwfOWoSuMdroSHocyA4cw6SX2kyGg7irhJQ93QHSVg2S9ZKla3V055TQdh/ZVrKtZbvIRoK/S9J0Z9sba90QE6xLCDHSWXlprTydiTbH7ZJZzE2hjOiJvCxpvKiHNUxb7AX2RGZh77CH2Es2p20ibw8YAoaAIWAIGAKGgCFgCHQlAkZYdCWaVpchYAgYAoaAIWAIGAKGwIZCgL9rETqeJEOHYoYsUzDYcwJXt3Ly3Ou7F2XxsS58KOMUOpoEpIRqF2EhRzH9oR+cVodM6C+DUOHUelf8DQ4RQpSDR1Lwm3a6ihBpbR5xiBNxQroghMm/lM13x4lQdLOuxYZaCN/ydll7HmEBidGu9ZY2Zt6HjCBKiNRQa6wHd+1z32snHTL2DHuHtcteYk91xXr9lk+Ldd8QMAQMAUPAEDAEDAFDYH0hYCmh1hfS1o4hYAgYAoaAIWAIGAKGQHcigKMcB+xC2fdkRB14f+t+re/PuE7Y5XLYrhF90Ur6JOpz3KgBHLnJDqQ88jQAcOxDJOB45tQ7zmRSS62r/gT1YZAoXtqebGmwuhpz2iQFFETFRBlRI0QBDHX7YoRFJxDPsv46SlSkt8q6JUIIsoEIoeWZXWIPaF1zHWLir7L93PUJqYaGBfP6hoy6bE47Maf2iiFgCBgChoAhYAgYAoZA5xAwwqJzuNlbhoAhYAgYAoaAIWAIGAI9BAE3moHT5KQl2kM2LKNrRARAWhAxgbO9Q8UlKTrqQIaQ4B3SQUFaQCxwDXKBv8GzpazqSL+8+jlBj1Oa0/ie9kZ3aw54UQAQLzizSaFFtAfjzerc3nrnH6SPzdPe4BPzyBvvJL9HxqTG+N5rd3cU+47guNE8C+nhpoDy8NxWg/tA16p0L1tqKfYCe4L9gXmF9TlMxl56U1ajOlhbLUi2btRI2WjmxAZiCBgChoAhYAgYAoaAIdBxBIyw6Dhm9oYhYAgYAoaAIWAIGAKGQM9CgL9pISs4Gb5/lq69omuvyd6XdUbEuMOjheSQkxc9AvQEOMkOsQCpgpO4KxzwXuofTsSjlYFDGof/ukZutGestEF6LdJlcYofsmKuO84W7Yuo8FJjecQEn6TFQnuDqBVwwSA90MWABIHMoc4lsirVwdhaTY8kQqM9fd7UngFb5uZQ2Ytai+9miQ4C03dcbNEj4dn0wl56VMaaJU1UC9IDcsRIi01tWdl4DQFDwBAwBAwBQ8AQ6H4ELLy3+zG2FgwBQ8AQMAQMAUPAEDAEuhEBOU5JhTRFRvQCQsLpBac3ztgVXJSDNVPXoht7lkon5WlY0DeMlFA455ujIDri9M0iogwhkB6Z0Kl62wJBpIHX/4QIghSG6kuKhGlsbMyPNkZr3ntnWv0nH3+WmPrW+xBIHhFBhAlEDX2EiKB/EBMQOZ/IIFww5mmsbJSMVFN8f14G0YSjnFRfkCR8p/0UMUL0hfrmsyiMb2YwTXx7X10lSgKi7mmts8pvnmr6pmfBngK5wXN9M57ZS7+Zt6myVIq09NKRtZv5rv02BAwBQ8AQMAQMAUPAEDAEsiFghIWtC0PAEDAEDAFDwBAwBAyBbzUCcrpyYv8k2WTZKRmDIaUN96pkRDpEO6BD0SW4uBoY6X93f2tS60AGCARPzJt+Y15EROLgww/0vfrSG5GaqppSv9/fUF9fzz0Ih3IZxMVgGSf5IWqILJklI0UWGiPYoY7PF1MjiWQyOVq/PQc62ENOPCTj+j9ln7n1QFwg9O2l94IMgcSgrx5h0xzFsqlFYKSRWkSxnCSDaICMgPyhpEfiQEQhlg6B9DfZDu4z3scd+vKBe4+0UC2KERaZiNhvQ8AQMAQMAUPAEDAEDIF1RcBSQq0rgva+IWAIGAKGgCFgCBgChsB6Q6CVCAOiGLaUnZylIzhkibBAQDi+vskK+tNJDYz1hmkbDXHiHuc/RIUXOYHDGyd33aMPPAFBMUC2m+wj2XDZCBkkA8LNEBCc7EcE2i9yYnOfz7enPif6fHo1GXd8gZATCIacWGO9k0ykZCs+0ycRFghCH+32b3N9PiWDrKDN92RfyTj9z28IC0iROTJScUF2rI/0WG73euQHmBPNs1TWX0a0iyfSThoxL9LH2yN8ZhYIwDtl98m6Qiy+RwJlnTIEDAFDwBAwBAwBQ8AQ6DkIGGHRc+bCemIIGAKGgCFgCBgChoAh0DEEOFHvneL30iJl1vAfXeBUf4WIg+4Wo+5Y73v404qugAiArAA3PomMIGKCFE9ErBDZwsn8SbKdREJAUIzQp+NLJifqhYDfH4gnnWSurkzy+QMj/IGA5sznBMJhJxSRzrOeDYRCTiIed+pWVegT/sEnBkMNJmIpAiOZipVIQnykayxsr99ok0Bq8ATOdqIu/ub2D2c8BEar2hc9HP5Ody9DfPs5VdQ0L46zs+xpFzNw87EnXK0V9gh7hdRqmYW9xbxDdjBBXaHB0unx2YuGgCFgCBgChoAhYAgYAhs3AkZYbNzza6MzBAwBQ8AQMAQMAUNgY0YAwgJH9deyOVkGigP2Hhmpg9bIv78xA9NFY4MkIFIBAWxxCz4iWbZ1fP7++v5mMpnYRq5r7i2QD7uXLxDcOhjO+UKfdfFo4wS/zz85GMnJgZQQcVHlDwQhPoKxxgYnnF/ohHJEWKgkErrc2Ji6Fgzp8UBgpN534tEGERgxJ67IC36nnmtiLyg40BGFJk3Uy7KhMrQxdpKRuoh+f0rfRLyQCiy+IXUuMiKDvPRgqcF0Y1ol6kcMHTH6bV1MXmcOmE7X6AJ74wsZOiEQFke6GHsfc/SFPcZe2+QIoAws7KchYAgYAoaAIWAIGAKGQDcjYIRFNwNs1RsChoAhYAgYAoaAIWAIdA0CWdJB8bcsJ/w57Y/OQmYhFRHXV26IVFBdM+r1X4sc/JyoJ4piiKxBhMNmPr8TFOmg74HvBILhIYqW6C0SYT9/wJ/rD4TuE5kQ8gdDY8I5BTWJWOMOoUjuKP0W9xASx6DMTD5foX47fqWBihTIV+4PNHnM/f4UERFUxIXfX5T6HQjnKrIinjIIi/qqlY4/FHViDXXKIOVFXeCLTyIUvaMMQoK+shZ2lUFU4FgnIuBd2TOyLzSu+g1JWrgzmRIqd7+TYqlbon7SSBAiKGaqHSJSZsjQtYDAI6UXUSj0ATAheNAUWUOYW9fYQ5Aa4EuEBc+mCnuyGwkXrxn7NAQMAUPAEDAEDAFDwBDYhBAwwmITmmwbqiFgCBgChoAhYAgYAhsRAvi7SWuDAxZn9YFZxoZzGE0FTplbWQsCLkkBUUFUBSmExigwYrNgxLdKn/sqsGEbfyBZFMwNDXYSfpEJTt9AKK9AZIUTj0WP9yeTYb8eFFkxQZEU4jWCIiEiIhrCIibIAqX/FeuR8o3re4rEUK4oER8+kRtNPfM++R5g6kgLJY0LPtUBvkcbGpyGmpWpqIsEehdNERfMPeQEmhU0MkeG4x2nPLoNhHKg2YCjvVMEQRpZRnc80eqORkjwHoMlKsUFI0UEdKpPTaC1q4AH0RMQD8wtBB99wCAsKN5eaQK+ZQHff8nAj+gVSwvVLtjtIUPAEDAEDAFDwBAwBAyBziBghEVnULN3DAFDwBAwBAwBQ8AQMAR6AgI4jBF8Plg2KkuH3tc1Ttsj1NxmyRLBkUrds7FGZ4ik8FITQfygR4FGBXiGxSmMF1NwYDDsm5hb7BtQJzrAJ/mJ8qFJRUAkYrWrAnlVFYJfhIEiLsK+cI6CJpo0m4O5+U3REyIo/H7+uZFU5IRLQIh5UDop7qWnJGp1bngvlFeot5JiKOLhYCQvIFbEiYsIaayrUaqolO8cMe9iT+xCF/aSIciNhgUEDGmi6MCHGnOdoiyIvuhMYTCebgcNE9nBZ3sLJAUkAXXg+Af3XK27Fd2sr8L6f0eGEDpC3PSBaImBskVu53mGvcKe+WHGgNhbCNo/KiN1lBVDwBAwBAwBQ8AQMAQMAUOg2xAwwqLboO7MNqcAACAASURBVLWKDQFDwBAwBAwBQ8AQMAS6EQHP4e05jrM1hWO2syfYcSanihzKCTmUO+vk7kYIOl+1G1EBPkQeQFRw8h+H+ljZsEDI/6u8Xkmn14CktCUCy5QNqjQUSdRFCpKxhtrckliDL5WiKRhSJIVkKoJK40TKJ0gDPomgSCYUFaFPkRNgl/p3h6IkqhR9QXsdKZAcyhUVjKqDPn8k4k+oXje6oymhUVKkxTcFPYv+MoSkMSIEDpI9IntTY/9En5UdTA/FegMjnPxEJeDghwTpCGFBBAjvgrmnD0Lv6Xt3RlnQ98UyiL1xMkgHfldpbacCWNz22SspvZIsxSNnvH1nwtutAGWXDQFDwBAwBAwBQ8AQMATWDQEjLNYNP3vbEDAEDAFDwBAwBAwBQ2D9I+CJbZPu5weyE7J0Ae0CnMPk6++oc5X6cSrjRMY4BV8v0qIjzun1j0obLboRFYyNfwOQHohIhAaRAVFFMHDqn5P1eytLk1PUL+z0HRV3ivpGkwpo6CVyIJDfq66gobbeCefGlLEpmOIIahXDEK2PyWqdnMKSVCRFIh4XmSCNim+SCzX/m0MaFe2KdskYCg595kOuffEW/lAy4W/0hfMKUoRITOmh0sS4m171+cK6tpm+kRYKZ/t4GfoWL8rulEFeEOXQ3uI59nHqs568z6DWRrydUTgQFqRjoqBjQR3dKmKtvjHPjJsoCUgcL0XWk277HlnCmNgr7Bn2zjYZwFys32hcQHYQlUF6qI7uq/Zibc8ZAoaAIWAIGAKGgCFgCGzCCBhhsQlPvg3dEDAEDAFDwBAwBAyBbwsCWdI1EQHBaXdS22SWu3ThPdnnsrp2OpPT68CJS34jCAoMRzORFr5O1NUjIHbJCsaEUDXO/4Fy6o/y+/0DxDJs7Usmpjg+/M8Jp6RfwikfhhA2uhEJXzCcCCbiASevhHRQTk3lEqemodbpk1Poc0Lhamf10qT0JJoyMpHpSQSIpyXRcuzJ5EdycZem8kV1shBoEc4vjEonwxeLNgQUreGPKjVUtA7ugf5LR0PC3BIIJ5ojKCIGBz2khVeI7iDiokaYPMv6aGekBZXzbyfPwU+EBA58HPdopLQ3AgcCDKICjNKtk4hkf01rFboIguIQ2b7uU8MYtwywtpZBnkDmeKQe/frYHdN0fWamhvLSSPFOs/B2l3Z8I64sJzc379BjTjz13jtv/eNGPMz1MrRAMBgUnPnVVZVo11gxBAwBQ8AQMAQMgY0MgfTQ6Y1saDYcQ8AQMAQMAUPAEDAEDIGNFAFc3jihcaCmO6O94ZLuhmdWylJkQwcL7xAJgBPaS4HTnSl7Oti9jj3upn+CrMB5v6cMoXJSNfWRJsQOkfziKeG8YiecF5ybUxBwBk6IO303q3UKyxudfKWFKhta7/Qa1NAYyvXVFPVJVhX3i6+qrghJI6Ih1mtQldN7aLUTyhFUPoVWUK/f9w1WyeT/dAk9CRrcQhEWOPnX6WS+ojhqApHIywr6eDfg91eEc8I14TxSUonDkj5G05Sl2uN/cdwr3MOHgx0h7smyY2TnySAvAi4+bYFKnxXKkSItiEZBvJrUU02RH+0vXj2QBRAEjSLBOrNGW21RZAWpqyAkICpGyqbJ5sggIdgTEBT8OxBs0vtPP7jvpZDKbCN9z60D7dR+sDamJ0/8yc/Pv+Dyq28cPW7CFhvTuDbEWH5w6hlnvzBt1uLS3uV9NkT71qYhYAgYAoaAIWAIdC8CFmHRvfha7YaAIWAIGAKGgCFgCBgC3YMAzlNOgJPuJrO8pAs4qHGUt0o0uKfQceTjqI2lOY6Tugdhwd/K3G86ut/DT5XL8Z4NaRzTpAWCrEC/4ABFQExXZMIu+jwglJPnBCO5Eq9WqqecwNDew+XBFmkRCMWU+inRkN8r4SssjwWTiaiiGZJBcQA5uUWxsrxesarqZU5NMJIM5pfGYoFQ8quqivCAaEOodyLurPA5yaUiCRS94byh0Ive+t7klE8mY4rbqFPbwhbjUnKufhMxM6yNpeJFbszTCevKQDC/IVCS8PvUMX+wdtLqxXmRWEPIaaiuJDJEk6b/E4eitFEKIElQf7Muib5PUp/2000IFQguyIi2CmviaxnC5JBZpEZaKGuTzNLayqy7S0kKKnfXc199nSDbWwYx8YIMoe3vyYgEYby7yTw9Dkgc0kAxfsbBnoGQITrpooxOs9fA6moXh7bwsvtpCOyy134H1tbUVM/+/BOIIyvrgMDELadsFwyGQrU11R1J67YOLdqrhoAhYAgYAoaAIbA+ETDCYn2ibW0ZAoaAIWAIGAKGgCFgCHQFAjjhIRG+UUn4plYcyTNlPOPpDKzRZprYsHfaPwxJ4aV8QmQ7LQ0VzuX26hR0xfg6XEcWsgKCxdN+wInNifvBIgaOIxIhlJvflDopEBJhkSdyIk9ERdDJLalwqpaVJQPBmprifrWrcwrjxT5/MqxMTM0F+evcokQ0FHFmi7CI5az2KfVSPJ5fumrZ8rn+FTWr8vP1MGmDlDbJd4hIC7QkmmqAmEgkG0QirIzHojjFld0pVCvBC9I0tVXUfV6IjwtG4uVKYbW4oCwR9znx2pyC6DN5xaFdl8+LlASCZU591eqUtgUvJJNZgwFCunqRHkC/47/Cj7XEPLeI/lC6qPQ+edoVOP6pdImMCIl1ihhpa9Dtua+1SrTRJNn2MggL0kGVy0bLnpC9IXtb5kWZEB0CaUFh7HM1jpWqhz0DKZMi8WSZ/17kWU8ovMtJl/aM9dv4TJ9+AwaOmzh56w+mvvV6QuXbOIae1GeiVGbP/HRGfV0dZJsVQ8AQMAQMAUPAENjIEDDCYiObUBuOIWAIGAKGgCFgCBgCGzkCOL49weJsp+JxIiMwvMB1uLYGh+fQ5+9hz1GNgHKzsDakRRt19FSovbERHULqIk7GKw2Sb9cmgiJX+hQRRSFIlzrle06KL4jId1/iNNaEKuOx8PLckmhOQVktmhUx3a6Te54HwZ1S5/cnKyTOfZ+kIkblFidCuaudpbWrgoNzixsqGmoj+8Uag6R+6i1iot59X5EQfogMpYzy58ejjcvEVIyWOLc0NXztEuIW96BgikS9X/EePl+yLhiOB/OKG4NSrViSX+afJtokHMmv3G7lwmCv5XNzUoLcjsiKZGOd4w9prPITQ9K4JSKiYoxq/LM/GILYeFJ9qmxNzyItQgIceoz4utYr+4HoGdJcKT4mFUVDqZAR1gFxBIH3SWqim0iID2SIkDOfRCJBdCAsP1ufpIRq0jhpImT4TC/sOUgN3uV0uznfMwDK9nP/7x1xrPRi/J98OG1qOx63R9aCQG5eXv6gocNHPvbAv/5uQBkChoAhYAgYAobAxomAERYb57zaqAwBQ8AQMAQMAUPAENhYEcAZj4Mbh+yRGYN8V785/Y4zlXQ9axNCph5OmOOc9YQPVmwEoDEWiApO3CMMfYCMU/e7+AN+6TwEnUQsKsd9WKRFbirSIiBnvoiDZKwx4GusSxTkldQ6sYZwYzwaqvY5jZWiM2rk9ocE8kSic/1Bp284mDyYeVAERn3JgJphNasLo6sWFQ31B5Ke0xxoGxKxhkqloAo5fl+9iAH6FNfPQa7GBHPENS/t1hpT0CRLkaz0BxJOKBJ7RbOVHwzHysoGr2zIK6kL1KzMy0smQ8P12LTSIfWj+4xqqJ47NVRc8XWgqK5SAR1xvyr3i6iJpKIuGH9zSSZ7SZz7el8gFBeR87Cuf2vEpEUwsHaJpthcdqgMQggRYj5J7YS4M+mH+E20BeQFBNYXMsiJITJSqwEIJ9V5DjKCvUNkxpsyIjG2SZsU9tzZMvag6VikAbO2rwcfedxJ3J8/9ytwt7IOCGw2fuIkyJ8ZH7zPf++tGAKGgCFgCBgChsBGiIARFhvhpNqQDAFDwBAwBAwBQ8AQ2MgR4OT4XjIc815BS+A9GY5UTpyvjazgHZzvOKebQgyaUt98a0+Lk7rIFY/G+Y/GAk5sTsjvJDtR0Q0S1S5yU0HFiXJIkRfBcE5MItk6pS/aQSjUrsr1KzoiqCsrFcEQF0kQDudFK8J5jTi8cWqTxmmijNP1YL1UXmvaHBPJa+hfUFYzWCyHE20IKqKBkAhfJBCKlKHwrYgGvZNEnZuQBjBHePpFWdZ0UHqDXn0QyW+IRPKiNapvSSi3cUYkv3FzpYQqDIWjoWBOtJ+iPUK5RQ1z+o2unKAEUYr8iIcjBb6K2HPhSeHcfL+0LZyGmjonHmtsYqY0uFT0hVsUedEn4UR/EArlvb7T/mcuev2pP7WpSdH88gb44kZVoEsyRXaIDMIB3Qn2A2TEZzLSQC2VDXON9c1zRGGwV9gfzCmQ/FsGIUW0xisy5pY9RJQSxCBRFqwpCm2w99DG2BgIPndY3fexw6577jti9FgiWpzFC+fP676WNo2ax02YtBUj/eSj9y1aZdOYchulIWAIGAKGwCaIgBEWm+Ck25ANAUPAEDAEDAFDwBD4liKAQxUn6+GyKzPGgEP1O7KnZDgFcci2qi3g6g40yPkLaeFFWHQJYeHqY6Tn+scB7hEjLbqdRYy5U1PjkhVElhBZMUa2vwxH83eJZCDtkcgJJ5SjiAqlg0o57ROJShEKGrOv2GsUvYfG2lDeygUlQ2MNwa/ye9UuUceLA+HY0kAwJVyN05tT+JANDYpeqIxHA4GGmvCixtrwAH1vTMZTZEQqfZSiF6rVTqPaL1VbONVTl10jQmBbWTrxlAq8SJEVvmS1PufoZ60Ik0hJv8pVodzozLrKHL8iLXJEYAQbaiKKnIguEMkS1nsDw7mxhZrNioKy5Ijh2zS+2FATHzbvw7xRlUuU2yoWdKJ1SiAVS4i8UJRJKtKkmdfaTZgcpnfvEJY1raWG6tTkdOFLWltgBekwUnasbAsZKZ4gKFjHiG6gR8HahkhCcJuoC+6xHnifeXxNRoTFYBkgPC0j+oLneYY9RGQFe8ojK7yR3Kovv5I9IIMU6ZJ941W+sX0ed+oZP/fGtGTRAiMs1nGCx06cvFU02tj4xaczPlrHqux1Q8AQMAQMAUPAEOihCBhh0UMnxrplCBgChoAhYAgYAoaAIbAGAjhScbDiMG92sqc9RbqVf8lmyNqlM+ASF10mmuySFfQT0WMc9BipeDitTv7/LmvLG7dLVpDOByc2KX5wTHMKWQ5nRTlIaCIQCjmJRCwVWQFZoVITjzbM1D2//l+n631EraQKpEW0PuisWlTcuHR2778U9688WkRESNETMaV7iopImC4iYaUIg8ba1blDVy8u7FddURAT0RGuWZGXW18t/QhFV1BUfwHtf1M3ERZOrcgL0nF54ukQOs0PKTuTSIiYI7JkuaIrkjmFDYtKSf9UXDdF7W2zeGb5slBOrCG/tHZY0B+vrqvOKYvHA7m9+q9O6N2h6l+O+JlefUbFG0SYzCsdEquY+15k+4aaXKd6RdiRMLjICqdFm+pjRBoWmyca4tupL9NkPS56QGuLNb+brJ8MsoE1RrQE0Q4Y66tSa9pb+5BxREtwHXzRsvB0SLhOuigIj11kH8tq3HnifaKVeA/B9GHNE9j0hX6wB9mLaF60S4Mko45N4ue4iZO22mmPffaf/sF770yYvPW2FmGx7tM+XuLlsz77dHpjY4Otu3WH02owBAwBQ8AQMAR6JAJGWPTIabFOGQKGgCFgCBgChoAhYAhkQYAT+TjiydufreCAxTGLM3VDnfrGCQ9h0UfGSXi+j5V9KMNhTN86RVqImMg2ZpgBcIGoOEgUwf6KNNhBTIGIhVRKJscXDCuqIlcpoQpT5IVKtUiLhdKvKNBdOa59nPrGAU50RnNReqWBCz7pN2b5vF5fhXOjJQM3XzQ9lBP9ShEO5cFQ/L1wfmPdos/6/lDRFX1qV+UVSgNDUQ8iA+KtSxuoO3KG+8CAU/5gA3HAXHmERVRtJEROBAp6V9eLtCgpHbSqn67107ulIFc6eNXE+qrIUKWvKlA6qJL62gjkBumvlirioyDgj4N9XSDgROJJR5EhSX9h72hOyYDoyF51vsKcvJAzf3okkEgGJI2RaCJwpEAej8V/JLaG1Eh3CetHwUmRFhs8PZRLgkE0HC/bWvapDIKKaAhPUBvioF5kRfO657ve5TcRFswtY4GoAGvICEgK9gyRFWE97+l38B5zxHPcJwVUZpmsC/xbkhRh5jjOAhCXTjv7okvnzfly1rR333xt1JjxE1atWE6KLSudRCAcyckhvdbD//7HHZ2swl4zBAwBQ8AQMAQMgW8BAkZYfAsmybpoCBgChoAhYAgYAoaAIZA6jU+KG06XIyKdreCQ5ZT4hiIr6BNOXk6+QyAMk6H7sErG390QCziCu6rADOD45zMqzztxDTuQ/kmpn0L+gAS244JEF4OhiKIsIov8gVCuSIxKRVrwHv3BSLPlnbxP71uBCICj61bnzJIlqyryeWaKoizGSNsix+dPzBOJEGisC4X1XKmiKrLV4daXrBXZIBEJH+3hbGcuKRAllBSJo+iImD+YAKs5iupYUFBaG1S9A+oqcyOhSFSJn+JDCntXF+m5goq5pVVKW1UlkqSyoTr8rgS/64v6Vo3PCSb66r7yXjmBQMiZnFeSrBkwPt6o7E/zGmp8iUTUKatc6u+/YkHYSSLIjXgHzfP/ydTaQrj9HdkiNz3UBiMtRBwwT5AUe8ogDsALPYQ5MnL4IxT+tSzqRgu5cDZ/eLojpbri6bTU6tmY6oZsuAnYISv0O/1d9hB7qbWxgxPO9xy9V51OlGR2YFP9PX6LLafsts8BB19y9mkn7qwoC6WDmr+pYtFV4x47YYstA8FgcMaHJrjdVZhaPYaAIWAIGAKGQE9EwAiLnjgr1idDwBAwBAwBQ8AQMAQMgUwE+LsVZz8CwaTFySykgrpNRk79tgS3uxNdTysARzOpoEh9hJN+nIxT8Gg/dFX/wKSvjGiKKfL2741GRaSg2BEx4SjlUyoVFP74QDgcDQTDhf5AoEAXSHcEuUBfvT4S7UA/M8sKpYj6Uhe3EYGwgz6D8ahO5Pucvd3nVV8qFVUbRWEMvlREBUQFJ/lxiKdyU6ngFKdP9GWggh6SSkPlFwkSkDaFiAZ/xEn6+pJyCmJEBElUREWeNDOiui+R6aRP6av2lTB3fWF59cImPe+UaDRfImhihHKTqwMx5xNpWLxSs9xXk1sSvTI5L9k/gTC4/i/pEhZ6BQxIk0TUAdEIPpEW6z3Swo2qIJ0YOhWIkpPmCwKBdE2kgbpf9jbfRRa0Sqi4JEaNGzEB3gmPXIC00G9SlWUr3JslY09BEtKP9MI6Zi+yJ1mHXnRGK9VtepfPuviK33/91ewvnnz4P/ccevQJp3SEsOjdp5/WZjy+omIZ/z2z4iJAOii+zlCKrY6Cov9G+i75/R//MmHLKdudecLhB6TPR2FRccmFV17356WLFy648apf/6KjddvzhoAhYAgYAoaAIdC1CBhh0bV4Wm2GgCFgCBgChoAhYAgYAt2HAI5ZHHhEL2QWohg4ud8tOhEdGBJ95OQ6UQscWUe4mJRQOL9xyONs7jBhkSUdFM5nnOuTZMuU6unEYE7e7rlFZSlxbZ/yIYVy8pxYQx2RFfFAKBxV5EWT6LXPR6oqHM2cvici5DMZQt2QKzjq0wukBif5ISUgOfj3Q5H8+zixGRPEQHsKYwYP6kg5zmU4uT1tBSIAZokciUbrw71FSlQX962ardRPEDLbi3QpQFujZmWeE86JzmusD+XombJ4Y2An+SEVTZKs8AUSs8J5Uer1Ik+omzGtEmmxUAEnyUhBsn7YNrFBirSYkWh0Fiz4NDglHm2RoYu+kXbsLdmfZc/JXhH+OOjXIAaUMqo9Y2/3M2mC7aRw2kOG6DVED+2LnHEekt0nI81TXStRFWu055IUHYk8AhT2EnuKvZVZ2IPsxQ0WfdJuUDfAgzvuttd+2+60254XnnHyMeId4qW9+/T99OMP0AVps+BYv/PBp195+pH777352t/8us0XNqEHNp+09Tb1dXW1s7/47JOODnucyI5DjznxVN7b/3tHHPu3W2642qvjl7+74db9DjrsqLlfzppphEVHkbXnDQFDwBAwBAyBrkfACIuux9RqNAQMAUPAEDAEDAFDwBDoegRwPuP4/66ME/BewemOE3yijGfc/D5Nt+Wo7fqerL1GHLikysHxDVnBJyLFj8mIVOA+DvUO6VikO8ZdkW2c2JAAo0VAnCtSYrecwl4O6aAwtCqSScSrc6b6g+GRgYBfKaOa0j7J+U/7OK85rc/nVzJO8PMdBz99I+JhgIz0ViNkc2TgD6HRy32WaAn60VZhzDjYP3DrHaZPyA5S5NAubRGBcoDMLy0MZ9lXZf2rlhWMVSRFoLhfpSItAo7SQjkiKBRB0rCgvjoyOFqnlE7JVJ9XBKKBr3KL6qcFgnHGyKR7Ggw43LlWTIqoSH7ykHBusjIe9c2ddHD03foa351LZwd+qvusn8zyM7fPRDZ4JEuH5q0tYLLcB1vSLY12jUeYE0+4HQIF7Yp4e8mK9vaBvZKWFsrbR+wpDxtvr1Ele/BM2eMyNDWsuAhAOJx54WW/JW3Rs489CLnk9Cot691e/YqJW22z/eBhI0Z9PuNj9ouVNAQ2n7TVNp9O/+B9SKCOAlNTXZXKebZyecWyZ9x58erIzc3nvxPOf/7x15s7Wq89bwgYAoaAIWAIGAJdj4ARFl2PqdVoCBgChoAhYAgYAoaAIdCFCKSdOidq4fKMqnFG/1eGUxmHKk74DVZwIqu/HmmBvgAOfk6okw4Kw8G+rk5vT9ibqARIkd2IqghKWFsERULaFW6qJfmaA6Gxji9RGS5oeCsYTu6mtEplsQY4hmS9IhY4tQ954WlYgB9RD5zuh6yg0H90ExBfJjKDVFdehAjO9fYU+sOJfASt+feHp+tBR4j68IidVF3SrHAaayKKDgkqKVQiKtHvuL4XKSVV6n7t6lw0JhB9BsenlAIqR0RFTOmiqBcShTFBkFAgi3BGQoggLh5XcqqGQDg5p7hv0r/TiQ21T1+Xe2ldpe+hVmZlH73zoox1RZ0QLc3zR+RLV0RZaM2AEcTQZTJSb0F60RZOVsZL+iXS4KzoaqLCxSnbB2MGUzQy2GPfy3iIvUhaqpns0fXYr7V0ecPfOuDQI48bO2HSlqceccDu0kdJrZUC5RyqqlyVLVJljQ5vv8uerDnn/XfeeHXDj6bn9CC/oKBw6MjRY1674+YbOtMroieuuODMH7396kvPL5o/jz3VXC4846SjR43dfOLH779LZJUVQ8AQMAQMAUPAENjACBhhsYEnwJo3BAwBQ8AQMAQMAUPAEGgTAZy5OM4PaeVJTtS/JOPEfrvS3rgkCPV6J+ezEgmdidBwSQucvRACOHyfkeGs5He7+tcaInKQ44zHCY/DfidFVxzt9/sVVREkBVRSYtqeLkSqCp/fV6CMULOKymtXkGYpktdYumpxEaINBfqfeqVKavD5k0tFEnwuPYdKfUJIQFikF0gh7xrOa9JBDW5j1jzHPmmFmB+IBNJOgQERFRAYWIv+enXKzZsUQfGkbKiuLZERdeClAiPSg4iD5er7q+Hc6PiBmy9aXDpImZ/8SU8zxBsHnxT6j5OSdF2TNe7BojVyJchdNn6v6KtfvB68sXal/yzpc6Q0P9wyR5/DZNfK0HpAJ2WqCIoUYeOuIc3FzbRJO/PXpifRXGvaF7cO3oesOFpGjn5P5wMMP5ahVzFjfQhbZ6z3hPpHCjNSgh2Urf+6xp6cISOipcOn3lup81t7OZKTm0t0xf+ee+qx99567X8MJByORBCKrq2pYT7bLKPGjJuwcP7Xc4gEaOvhvv0HDuqINkZb9a3LfcY+euz4iXW1tTWzZ37KmshahgwfOVqSEb2md1CHgnRQ+s+bf8a0jutXeB15+N6/356tU/R5bWRFvhgnL0KjIxgRbSPdoEA8FutwGsCOtGPPGgKGgCFgCBgCGxsCRlhsbDNq4zEEDAFDwBAwBAwBQ2DjQwCthvEytAWyFciK52UtHIJtkA04yjl5jzO9QYYj3RODXmcE3dPmMTfaAie/5wbvdHSFS1bw9zuO/1Nkk/xK/RTOKxRZkS9ywg+Z0bJIgDqR9DcEQvHk4FHLluQW1yXqq3IWLfikX3Uy7v9M6ZZyc4vrv65enr945fzifKVdGi3iIiHiAoIFRzq2mQySAuKC/uOcxznN92z/niCS4UP3OS/VFM8SIkGkBjjv5XaUqAWceR4ZcY++E3lByqHdZW/KiCRJpbNSNEW1iIaPFB3SEAgkVuSX1kSGbjl/Xp+RFQWKxoDUQlcBkog6iBwheoPCfNMH1gi6GH1kywVfw6gdY+HeQxNLZ78dfHbB9MC29dW+Egl/U3hmkGw7GXg8IuuleagQaUFdrB+IFNbmFNkLmu8H9bm6PdEGblQF2O4og4SiHogVoiogKkghRruMxZeWrmmNVGfp91I9bype6rGspJBHgHjREfpkfhgT8wHRROH7CzIiYfZMq9v7yp6k35BQ4L5JlxNO+3/n9S7v2y9dByEUDqVIs7i81tnAwal93qW/u36YogcaGxsattxmh52V8Sh+7W3/fCA1AXrv8+kfTbvr5ut/n/7+ZuMnTrr3qVffP+nQfXbynO041k8756JL9/3uoUeKIwne/sdrfvPvv/0FLRYHZ//3JP597Ck/PQtR7z9ccfG5j95/z99amzBIFjQf9jngkMPL+vTtN/OT6R9ef+Wvzl+2ZBEkVouyw6577vvbm+66VzwEe9X54rMZH5/34x8chuh45rN/uP1fDwfkxT90jynj6NORJ5x6Ov0qKCoufvf1/714zWW/+Hk2cod0UNT18bR3iepJldHjJmyBoDlE7QP/vOPWtREl6f0IBkOhI0445ae773vgIcsWL1rw21+d+7PWCAkIlvuff+vjc0499tDXR9CGHQAAIABJREFUX3ruKQiIH5x6xtl7H3DIYczN32+58Zr/Pffko+n1gwOi6/sdfPjRwVAw9Ncbrv6/2/90zW826c1hgzcEDAFDwBAwBDqAgBEWHQDLHjUEDAFDwBAwBAwBQ8AQ6H4EMpyvOF35mxWHKWmfshU0GHB8t4sMcB2zOMDRZ4AMwSnPCXFO0eN4bVc97UHCdVx3WX1um9QHwRKSPkVFMJLbO5ST68hhL9JCoQlKqYThrg7lRBGpdoZtPa+0oLRmgBz9vqK+VaMLymrer1ud+0Fx/9W7B4KJ7URS1NZX5sz/8t2hy6oq8jdvqM4pTcSb+Y9haovT3pABOPw9DQzwy1YgH8ASXNE/IGIApy3Y8okDHtKC+4tlOLo9wuI4fb9LNkRjyfP7k1tqXPXBSGyeIh8qJK69PL+0dmoi5l9YOmhlcf+xSwvDuY0RPYvDH1KFaAyc/F5kxr36jjYGfSbN1QT3OZ7n2XfDOcmC3sPjg3OLk7VlgxMvzXwtuP+qhf4ctZciSdwCGXKujNRM/xVp4eHAeEiNRYTEMBlOfxzNjLXVojUIMQCZc6QMQmS2jKgRyC00IYgEYU1DWjDXQS96A4JBBoYY/WINQ7pBTHii5p6GB+QHxAuF+eMZhNIrVIcX/VKm77RB8UTU39d3yBNPr2SOez/zgz3J3gxu6mmhyvv2H3DST39+wX1//+tNX836vFnXQ2fsU4SR95kJoAIT8sZtMXnr2urqKsiLYgleKMDiy/6DhgwNhUJh0kpVLFmyKPO9CZO33haHf1QsB/dKe5f3+ct9j784crNxmxO9MFyhGudffvWNU9987WVIhmv/cveDW0gf46VnHv8vxMbFV/3h5icf/s89sVh0jTR6JdLc+NPfH3iCNubP/Wr24oXz50GC4Lw//qA9tvNSXdEu/f+/G277O1EEt13/28shUvbY77vfu/DK6/58+nHf2y+z35Aln0//cBqkwTW3/eN+SAMIjk8+fH8qxMWqlSuWZxO+3lx9WVGxbCnRJ9R51Ik/PuP8y353AwQCuO1/yOHHHLzL5NGVq1eReq/VkiJrRJpM3HIK+y5VPlIqqNb0K0YrVRRRMoyZsd54138eQ1CdORKPM+CI40/5STph0affgIG33//ky7Tz2AP3/H3chMlb/fS8X17xxMP/vjszFdXa+mn3DAFDwBAwBAyBTRkBIyw25dm3sRsChoAhYAgYAoaAIdADEciIjEATAgf9LBmn7xEjxjGNsxanMSk+ICxwgLe38DcwDnLS73DqGQcXTl3ve1cTDO3tV6vPudEVOMOJbCDdCumNapXaaHQi1ugEwn4np6DBySupc2pW5jnxmN/J71Xr5BQ2fF1YXl0vgmKKohMGicrA8Vmi3zvo/gJdK5MrfwxqF8Gymq2GbjnPqZhTVr14Zp9QfVUkKoIDZzQOVzDDoQ5uxB94J/Cz9RmnOSmrcJrjAPeEuSE4ID5whg+TEb1AtAhOb8Y0UsYYRysiZJnG41f0x5e9hy1/X2RKXiAcj/QasDomMqYsEI7NKOxdUywyg8gGHPs44zeXMY8QFjjyIU28CBr6wn2u40yGwKCtRfo2WZEWhQVliarykc7ycF7yjrf+Fd4+2uBjfaSX/fUDxz5aEpwch2h5TQbZwHgZK31hTESGrFFcsgwy5UeyYTJvLROVQl1gQV1cp36IDbAnWsfTieDarjKIINr05gTdC9YF9fKdMdI3tEPA9hW3TogSdEloA20P8OB5+sVeSMcH3HCIQ5ygHXCqjDWBkxuyiT3J3ky2J6pEz2205ZxLfnNtY0N9PU779EEmpBDN70gkh/lao5CO6OTv77cLN4iu2G2fAw6+5tILznrl+acRNG+1jBozHvLNwYkPcfG7m+769/CRm4296GcnH/v0Iw/c+/8uuvx3Pzz97F/s8Z2DDt3v4O8fBaFw2F7bTYCAOPtXV15DNAi6EPLvtyDXiKz4o5zy4yZM2uqqi885/YG777gVZ/3xPz7zXMY4buLkrT/5aBppwlJlx9323q9MUSUXn3nKcU/9937Spjmny0EfjcbWIEL6Dxo8lOiDj6a9+9a5l/72D5AV//zLn6674TeXXJBQua1X6Qs77b73d7IRFpAtH0+bmoquOPiI40668Mpr/8w4f//r8/8fuiHnX/b7G4houP+ft9/SGmik0Prrf554CVFzIk/+fssNV19/x72PHH3Sj38GDs88+gCEZIuy1XY77RoVK/Th1LdeF8b3Ttl+592uvfzCs/91xy03QmAkFI/mvQAJc91f73motHefvicftt8un4mYgfD4z3NvfgRxYYTFRrv9bWCGgCFgCBgCXYyAERZdDKhVZwgYAoaAIWAIGAKGgCGwbghkibDAQbuz7AhZunYCjlNS0uCU/Sy91TbSQeFAxPHsnTjH+eylw+FznXQm1m30rb4NaUBEAqfeweFX/E4m404oz+8UlleKsPBLf8Gn71VOtD7k9B+7pKqwrOYjOf1niphAyJniRUWEFJXwXf0mzz4kQr5+9ykqr25oqI4slLD1AIlYJxtrw56mA07x3V1sIBdwrHMNQiBbgVhiTiCBPMKCMeCMx9ILEQIQIJ/IBquv+SX9K+9VuqrCwt7VfYr7VY1TREUglBvtJSIDDHCeL9VzOORxvBMFgFgunxBXGI53L3IDMoC5pq/0ByKDfwexljhljVN+lcS4Y4XlicWNNb5opNCJRxtShFZmISqDqIq8U485vfr2e29eqbW2Qmv2Jl07R8aa7EO6p3TNCVerghRVpID6voyUWBAD03heRgotfkPCQbjQNql3eIc1SX1xN40UfWY+GS+YeqQM+8CbF5zZEA2Ml1Q6W7r1QMZBvEBQzJSBJzhCfOBgBiu0YGJqb5nbb9phn2GMj8Kcgt/xMhzxS/Vs9aZKWuDU/o5O+F954VmnZZ7wj7mO+7z8fA87F8I1P4i04OqMD78hBFp7eKS0LiBIKpYtWXz4D075yTY77rrHdVdcdA5OfN6R7zy173501vm/mvXZJx//+Kjv7lVdVZkSo+83YNAQnPCZZAX3Tj/3l1dMFDlw6Tk//WF6yqipb776MvcRFE8nLAYOHjqc64sXzCc6KFVuvvY3v87W7/ETt0yNTxrkJURIPPHQfXf/4f9+eZ737Lw5X84aMXoMJFqL0m/goCFEsHw87a83QdT88nc33Mo4IUkgUz6c+vYbvAAh0hpekAs33PnvRwcOGTbikrNPO/HxB+79B8/W19XVMqbJU7bbMRthsd0uu+9N/d897NgTdt17/4No08MYsim9vRN+8v/OIyrlgp+eeCRkBfdol8/WUoK11l+7bggYAoaAIWAIbMoIGGGxKc++jd0QMAQMAUPAEDAEDIGejwAOWRymnKTfPUt3n9W1d2UdyZ8PYUGqHBzk6Bng3MZZi4Ovx0VXuGMGB07EcxL7bFmuHOxOKNKYiqQoG7LaScSL61YtKM0tGbgqkVPQWKXoiqpwXuMIRSHgkMZhT0RDeukjgmOLeNR/t9JCjRBhsac/mCiReHVVIuGP6qVeFXN7ObHGFv9kgAzA0Q3BgLOOk/7ZCqQP5EpW/YS0F+boO/NLFAD6FNPVj9mlg1d+Uj58+WClgspTSqvxuh5TdMhcfeK8p0M4PknrRBuQMAfLmD+c/Dj9IUFwytNfnPGkg2KecdCDIfPNyXLqgrzC6Z8bDDmjc0uSr5YPjzdWLw/O1WrIdICeqecgAhBSf02khRdpwolziIZjZR/InpOl1qQc+RAc9AESB2csfaGvOHjnyCAq3pOxJll/EEikhKJvPAPB4gla4/yE8ICw8NKkQTCwlmmPFFxoStAW7zPnHpFDv1kHkBJPyCDqeA4ShsgMom/qs5AO1MseA+/M+d5d14hwQkeGfm9ywtucqr/oN9fdhBM/m6gzuhQKsogXufoOwqjVMmHylG05hb9cJMTanuMejvsvRESIByk844JLrnxH+g/33H4zUTCpMkyefz6rKytX//zkow/xyAqujdhs7PgFc+dA/LUoI6SafZKiMp597KH/ZOpb1ErkgYc9nQrvRY/0gFRIrZK1lLETJ6V0iL5zyBHHzJn9xedXXfzzn6Y/nitWp7qqin3QokzccptU+qYZH7z37hXX3/o3+n75+Wec6qWmCoXDKZ2Q9DFm1nH5dbfcBTFxxQVn/sgjK0hxtcXW26bI3Ndffu7pzHdIjUWKLdJFnXnhpVf9TREZHlmR+Sy4nHzGuRehc/Hc4w/f790fozb5/sWnM9ClsWIIGAKGgCFgCBgC7UDACIt2gGSPGAKGgCFgCBgChoAhYAhsMARweOPgxVmfreCUQ+gYB3S7yAYcsnIic/Kck/U4tnHE4mAnXRDpbbKK424oBNx0UPSRaAKczmVKBeXkFiWd3sPoapUTyfWtzOu1slqp3Ot7DagMBHOiyUheoz+UEwspKgHnPvgwNhzznqZBUumVeou0ODbaECwWaRH3B+NV/lBikZD0Ke3SsMLymsjqxYUR3Uk5BFVwJhLxso9bV2uweKf2wXdtZRg3RapURQoa7s0rqp+dW1IXKh+2PCqB8JUa52xFUuBUx2mPUx4xbvqPZgTzR3omHP5Ee9Am7XEfsoKT3zj4GTN9xuGK8x0MOWkOucG7fOLYz1MNc4TrtNE7xQYvnR24pGaFL3UKO6OQFgmCAdLBIyzAhWgV+oXbdozWmCc8jhAxpAHkCtEI9AHHPv3lWRyZDR5R4GpLQFh40T5xd83SDfpJtFG6bgXjgiwgkoKxz5GBF2N8XcZ9yCV+Q+BApkDe0AfaJpqiRVRRWpQTe4q146W6og+Zhb3JHmV9fasICzeCBBHzdv23I9vgT/7ZuRfh6D/xkL12IK1Rtmfkg1+N8zvbvfRrW223467T3nnz1baeoy40K9Cj4FQ/0RtXXXz2Tz0HPmmdJm+z/U7Uc9Uvzzl96eKFrIdU6VXWuxwn/CP/uRutmBYFDQ5SWN1w1SUXZN7zIkQaFNWRfk9EyQu0u8te3znQSwnVWv/TIyxOO/qgvTLFtRlTZUaKKuoi4gNsx2y+xeQx4ydOPkFYExnhtUPUBN+ziXxznfRX+x70/SPv/utN16eTSswd6bRIl/XeW6+xf1sUoiW4QGTF8mVLl9x63VWXtja2w35w8mmk2Lr52iubo0siCq84Qam03n/79Vc87Y225tbuGwKGgCFgCBgChkDTqRsrhoAhYAgYAoaAIWAIGAKGQE9FwBN4zowO8PrLdRy7nXE44vCaI8Mhi+HUTQnY9rACaQNh4J3QLcDVLa0Fp2xoQuITiWRx/0Q0r6TeV9in5mvdKgqG430VqZArZz+OZsZFpADOVJz+NYqaWFa3OqdQ9RRE64N99GxAmhHJnIJEjt+fqOkzsiKnZMBq3+olhdF4bHCyammBxH9TItw4xCEQWksF5UGHUzOb8xpHOc775iIhbUeaGoleA1fvqOiOOrXb6PMnGvy+pF/9ox36D5l0uIwoBqIEiC7gZD+6DKRN2lkrYIh4FmXJ8n3QWB96JpwbPVnXc1RXWMQH7UIwgOF0Gtd4nhNhM1UYbabx49RnXOWhJhHuYdsf0zDvpdtyliTiisJpubroC5oQ6f+WYv3QFyIoOEVOpAP9g0iBpOA6pAZpmxgTRAtRGnMzyQLXeQ52LfAjzZlLJDAOCBhSbv1VBjHCWsbAnXnmXaJJ+ITYQf8iGxGXVfslPaWaqyHDHlvbHqTNZpV2fe/RxSUqIJAgW1bqN+sqpbnQWjo5UhKdfMY5FyrSgIP8q/gfHPWnnHnuxR++9/Yb0rEu3nbn3fdKyrGOA1z+9Fqc6vX1tbU44XtL52FtoChL0zA0FkRYoGWy1uLpV8ye+emM08/71RX3/+OOW+Z+OYvIp1TZatsddyHtEo7y55/4LyLwzWWHXffcF5Fq7qVfRyx6/0OPOPaZRx+6L5vWAvd5frVEsdPfQ5D7rVdfem7P73z3UMiQlcsrIM+yljETtkhFG9Cnz2d8RCRSiyKd6oGkhcq8PlH5mhZI5Pr4H//snP/8845bZnz4fotYjs3GTYDIdGZ+8jF7oUUBVzQ1SNH0x99eeqF3c9DQ4SO/+/2jSWnmzPr8k+mZ6Z24joA4n0qhNfj8n5xwBNEyrY0NXY2PJd7tpcsiFdQ1t/7zfvQ9zv3RcURFWTEEDAFDwBAwBAyBdiJghEU7gbLHDAFDwBAwBAwBQ8AQMAQ2CAIeGdGargRO2w5rTrhO4QY5KkmHk+5o7Qzx0d3AQFZwoh47jsZIBxXJTzqFvZPSrkguyilMrJCjXU70+Cg518GMUXmpr0gvg5OcaINnEwnf6lWLiqjrwGhdaIQvkIg01kScqmUFtf02W5oIhBJFSg1VFMlvTErYul7khb9uda50MZr/6YCzvq3iiVpnPteCrBBR4IRzGxtyi+oDigQZXLsqJ6l0ULkiTXJi0aCIhWR/ETJLRSzUp9JC+ZI4DN+CjHHx4DdEwxAREI3xWKCwenl+ztz3B5UPGL94Zk5+43iNJRrKiU6XkQJqqYiauQ21kZFLv+xduPzrXmMHT1w4pO/opYNEcOBQxnGtNp1JfUYmxpf0T/xu5Xz/9RmLAgKFNFSQBhBCCTcCgnchPnCekr+eSAja5BnwJ3UTz0BafKV3IBI6Wliv1Mn4aZ86IBIgR/gOmcFEMb9gTdfpb1BrfZ7a7Ig4fXrf2GPstT2ydJh7tNO07npwcYkKyC6ib3DA03cwIY3YGiLR6UMZL32JAw87+niICRz+6fcQy77lX4+Qnq7Vgr7Cfc+8/sHsmZ/NuPz8n53aIDYj/WEvImLaO2+0GWGx2fgJKUf6iFFjxpGS6o4/XXtVel3oafD7zpv+8LvMDu11wCGHEa3w2ovPPpl+b7+DDzuauloTrR4l8Wie/1J5qDLrJFUSRMixp/z0rJuu/j/0ddYoEB5lEqOG5Ln9T9f+JvMB2iZF0wtPPkLEXHMhWmScUkmFlPcJfZCbr/m/SzLfHS3CAsIBQfHMexdccfWN/kAgcNGZpxyLbod3/8xfXJrCjGufTv/w/Wx9RjCb66SvyuxX+vPM7dARozb73a/O+xnXt91ptz1/+dsbbhXHNYh0XF98ZumgWt0YdsMQMAQMAUPAEMiCgBEWtiwMAUPAEDAEDAFDwBAwBHoyAvy9yslxcuynnHQZhdPrLfzJbQhut3jdJS7aTVJkppDhxHt72vPeU+Oeo5M2m9tNr0MpoNL7yPNgQEooTuujueEk5Watr/Y5qxb5nf5j4qFgOMnJehzGRE2gUUDdiCLzDtoEOPJwYiecpK80EIzvLGHtgUtn947EpVERym106itz8/JK6uLSxKgTeRDTc45Et4PxaED1x5xYQ9AT4G5rvXhphEiFtNYiMsJR6qeIL5AMi7SQ8HWyvwS2p/rCycKVC4qTEgCvLum/esWK+b3mJuK+irIhK/PiMf9c6XPME6HiF4FBtMUeIjRWK2pkUV1lzrAF0/tvtWpR8S5KY/VQ2dAV9RpDbigSHVE2ZNViBWCs+mrq0PKlX5Wd6Es6Y5JJp+rLd4b+TZ/v9R+zpJdSaJE6B1IgGQgli0dsG5s5bXH4pXi0haMesmA/GY7be2QpIWMVyBM0JzhFDnGAlgRpZiA3wAJnKaQF6znhpV1qz/pJA5EoDVJYse6ZV9qAHNnc/Y6oN6mH5shwwrJ+cNCn0hGpzS87mf6IOaXNbIW9yZh67L8t3f3n6eGAFd/ZM95/X9qMrPrfc089tuvmg3vh/C4UaXHWxVf8/pAjf/DDi8889bjFCknw+/z8v9akz6edlE+EQ2FRSUlhcXHJnt856NDxW2w5RYEXUfns+wcC/jXInYlbbbs9URuc9m8F5+bLWyhFEpEMO++53wH3/f0vNy2vWMqaTRXSEJH+aMmiBfPfePn5FroMpHXaafe9v0NESGYkxM577nvAsiWLFn703jtvZmt/+1322AeR71mffbpG/9557eUXiNhASPsukSSZqZ6ob9zEJkHxt197+fkvPp3+UWYb6GpAWkz/4D2ij5qLsldtwZi4cItSMhHdkvkuz8wSKZCZkosx7bbPAQeTCmrOrJkQbqkCOQRGiGzvd/DhR/NutjEjbM71+/5225+9dFvZnkN0net1GvgdDz79ChEujPG4A3ffhiiYbO/YNUPAEDAEDAFDwBBoHYEe+0elTZohYAgYAoaAIWAIGAKGgCEgBDgBTYQAJ6AzC05U/p4lJRBpRDocadFehOXwxMHp6TEE9BsHJyl22k126FlO2ZOGxkvZw0n5tZ7qdsfHafAjZTjqhhJdEc5NOuXDE86gibElRX2Ttf5gKuUTzntSH0FYvCDjlDWkBZEVOOIhO4bIua86kr0rlxYWRetDjiIS0JBIubZXfN0rIMKgtwiBmAS7E8FINKp7SUUnNNZXR8KQGO0o9JNohbb0K1LtIhqudFTK5eT4Q+EYY60Qqv5QJDZswYz+gcplBYPVz11FnBRUzC1d2lATqR2xzVynz6hlC/1+p1SRFbMV/RGpWZFfrs+GmlW5E6XJUbZ6SdGJtZW5gyL5DY4iLfo21ofn63pt9fK8PVT/JBEaDCUn2uA7aems8ocKSmtHSLC8zO9PQgqsFh7FfUfHJ+QUJj+sXenbQ/3zCi8iEs7aC4lg8r/32t3MqadNwbghNCAnwBwHMOmfELlm3WQlqtqBK4/wLif5r5SRZoooGvQ0aItUVUTjkLJnX9nR7r1/6xOBZS/qpaMaLYyXPcZ4aT9zEbA32aPdtv/aiU3qsTT9DX5CHEHaNZF1TaQRRE96GrhVHSFxENBGS+F7R59wyh1/vvaqZx578L62+oezG8LirB8edXDF0sW0v0aBhIAsWJtj3Htpi6222wGRZ6ID/nnbn65Lr2yv/Q/6PlEgj9x3912ZdaHFgPM/M1oAHQcEv//33JOPZmtfut5Fk6ZstyMESHqUQnq7RHncdPfDTx9y1PEn33vnrX/MHCCC11x76uH//Cvb+Lfbabe9uJ5JWEyY3CS4TaqoB/91118y3yUNFWmXXnrmiUcy75EuCxLo9j9d0xzRAeF0weVX38j1VxVlAmHx1Refo2XTokCeDB+12VjG25Y2x+QpTXohl//hlrvmK3XVpef89IePP/Tvf7JW2lobdt8QMAQMAUPAEDAE1kTACAtbFYaAIWAIGAKGgCFgCBgCPRkB/l5F0BdHfLaCI7jVnOldMTD3dDany0mxg8MZhy0RD/SJtC5rJS3c9yENcPpCIEBa4NSHWOBEfrNTKyO6gu5zshjnOKf0cYIP1NnsWH6vZLCoPOEU9E5WSQNitXqAI/Yd9Yw2cJLjuCa1DCd/Od1P2qQ4zn0RD1+JsOgrEiKALgWOe5EBDkluRAg4uu4oWiGY0xhQJIc/rPRM3E+qDRzd7fn3Q4u0T1nmgHqa0iT5kiGiLII5sXqRFtXhvGi9SIxiEQuVCz/rG1fKpkb1a6kiPoYqlVVNMu7/TBEWu3368mj0NWYNnzKvl0iKWHVFfrDi69Iyfa6sWZn3pEiZ43V9EFEhDVURJ15a00uTtGvtytyQxl/kES8pEiLpKxcpcpTGPqewvDriz4mCN+TCnGDYWaRoluJWJph5BGcwAX8c4hAHOD85Tc78Pip7W9aCqACTDkZWpGBE70LrCcLiMhlrisgJtAAgFViL7AVvjTL3u8hYN6SFItXOP/R+RaZuRqrytRfqZa+1CP9xX2EfsEe9SJO26uqW+1mICki8yTLWI6QK80RfIe8g95YKh7YIwzX6ip7BVX+6/Z4Pp779xq1/+O1l7RlMxZImkqKgqKg4G2ERjuTkkObpzj9f99u26sM5Twoinvvv3f+8Mz26gmtEffCZLYWR0j4dlbr31KMPpbfTR6mLiL5A5yFb+9897JjjScn0XIYeRvqzb/zvhWdIF/W9VggLL8Li9ZeeeypbG0RDTHv3zddWVCxjbprLhC2bhK//+serr0QbJPNdT2dCfW+R1mnr7XfejTbBNF1345Qzzr2I61ddfM7pzCX1LZg3l5RqLYoX8UHqLGWiglxutaA9smrF8oorLzzrNITQWxNfb2tu7b4hYAgYAoaAIWAINCGQOlZkxRAwBAwBQ8AQMAQMAUPAEOihCJA6BWf7jln6B3FAWhdKd57u5m9m0urQF3QDRsiIBOBEOye421MgHjCICt7BgdoaCePVR7u8gy4C3xFzLpEIdLB6uU/kgl+6E76chipflZz65SIrttd9nNg8i6PaE+umDgiXhBz5zyrNEo69eH5JXUgplZr7jvNeaaKcRTP7Ootnlju1K/OcyqUFzvJ5vRylWlIERLuiK9rCAqf25zIc+9PijYF5dVU5C1VztfrmKHVTjciKJUtmlfuXzi4vF5lSKYKiqLEuNF7kw2TICr0XFoEySdEXQ2a9MXz1zNdGVnz13pA3ld5qcdXygtF6J5X+qKkkRQgll4mAgbjwSS+jIpwTjeWX1ogkiSJYLj0QcTEJ34e1q3JniuRI6jun8UuF6eq8kkTRpAMbF4UiSVI7ZZZf68JYMJezPBVtIUP4mDQ8kBScBscBjFOce1hzKiAc7BlO9rVil/Y8zu/nXQyJnKiX4x0nL23fLXtC9h8ZKasgMYjsIVUUzupbZJeprvGycFqqsrW17e0t9lq2RcDeZI9uMA0Ldxy0zz6lL6TKGiPzxMjZbxUyyKQZwmtBZ8gKUj1df8e9jxCF8IvTTzoqmwM9G5AVy5YQgeLodfq3RhkxukmL4pOPPiBaZq1l0tbb7sADOMVJdZT+MDoRU3bcdY+lixcu+GDqW6+n34OQ2HG3vfZDFHrxgvkQpc2lXGrX/Ggt+uOw4076MU7/5x7/7/1r69zjD9z7DwgEHPiZz42V4DbRB5kEC88NHDx0+DbSfeD9zPcQ3CYa4plHHiRSaI2y2djNU4Lbn378QQvC4qAjjj2R6w/e801UBkTFj8/+xa9ffvaZtxEeAAAgAElEQVSJR9DqGD12/ETmMpvIuKpNRYS8+PRjD7c1Jwp2KWNsEEFGVrSFlt03BAwBQ8AQMATaRqA9J6TarsWeMAQMAUPAEDAEDAFDwBAwBLoHAU6u42hsLYqBU+Sc/uZEfHcV2uZkL6l2ICs4VY8jFAd0LzlLl7XjxDrOVEgOTurirMfxC/lBgZDIljqEdyAaIEaaHYDoV8iZvnDolvFkUXnSH4wkN1NtRFF4mhE47oi0IAoEgiQmJ349kRRVy/L3ijUGwnLMr1q5sLhBItW56chCGkiU2pEYt9NYF05FX4jgINKCfraWEog26GN7ChXhvGU8S9R+48r5JaulkVGfJ+0MCWRXS+A7snxuaUD9hAzgJLmXFgz8iH7A2epX33IXfd5nZ419qMawSoTKKhEw9aJp+gjcWf5QfFQwHEeM21GaK6e+Jjxbyt7zwvmNU4rKq1NkDGMMhuKOPxifUlBW87zG79fzcZ+TpN0hgbAjvYzk+4pkWbVqga62XIWsA+YuMfXt95NTttsKpzhOfYgosCfSgf4y36wV1gzkBSRCh1PFEJHhEhy8y9qBiMA5j2P+PXcN0iZi8pygnypD94U8/PSDtQSm35dBaOHsnq5n5+rdNfqTRqawVvvIUnn6sxRQYY92VtC7lWrXvJxB8HjkCZEukFSQdaQVYu2zRvgNoUPf0Hj4vJNC56mOkBbpT/944ImhI0Zv9qMjD0iRAu3tuCQmUhEWAwYPHQZhkPmeCAsIlqyC1pnPTlTqKK69+/r/XswUmd593wMPIb3Ti0899lBmaqcddt1rXyI50OLIrNPTiEC4OvMeIt2IWpPyCQ2LtY35g3ebSJJRIgLQ0PCeLSkt6w2J8eYrL2YVJj/+tDPPVdV1zz72EERbcwHzYUrL9KzSbjU2NmTVGaFvpF5CzDz9XSI2Pp/x0QcLxSRwncgUkU3/1Vwsvuzc00/m2pDho0aj5ZGtbi+FVaYOSLbxF4mxyEbEtHd92HOGgCFgCBgChoAh0BIBIyxsRRgChoAhYAgYAoaAIWAI9GQEIAoQjEbolQiDzDJQF3Bc4hDusBO4nQPHIYuzDMc5nzijIUk41e6RDm1VhS4CaUdwLlMPwsk4+SFApskRW0MefWkhNNej9FCMCQczzuZUChhKQFeHbxtb3n9cPCKyIl8ExjM6276Nbk10+0NKKE5MY5XSfPgoHvXvoFRPQyIFjcMUbbBCkQozFKXwZGNtaIrga66b+iEplJhJ9k3wSIajPnOsbZEVOGvpC458CAvGTJRFKuJEERWPVy0rWFbUp7qXxLJH1FdFalYtLloh8gAnrucgZf4hLCjMOeTMSSIXFoqsKBJRkRuMxHyKGplb3K9yfk5hvU+aFqf6/IkcokYUnVGbV1xXXzJw9RhpVdSg21GzMtdJVPsrfJEYzu58pZ1qUB0rlAJriNtfdFEi8ZhvZtmQxLyqpX6lysocunO8rtx/6w23v6O5Y23E3WgLoh1IC8Vc4CAGI8SpqcEjfjobFeRFFkFYQEiAS4uT+UQPILCt6zjuSQ22swxnvhets7u+Mw8vyb7Us6/okz5DPhGxkfBSVukeC4E2wT1bYW7Yox3VxmilujUvpxEVrB9PSBwShTXC+vX+XUuKH9YWkS3MK5iz7xhTR/RmWnSCCIBrbrv7AXEV4846+eiDZ3z4/rvt7rweXLJwPunBnPE64f98lrRKAwYNHcb95W4kBt9xmM/98ouZmSTC1q7A89OPPHBvZh9222f/g7iWLXXTznvtdyD33nj5uRZC3E3tNol2l/YuB9PmApFx7iVXXUdKpL/feuM16ffC4UiENFbpmhOIjvMM4uLpz3ppmyQHscYOGinF7MOPO/m0m6698hIiKdLf23zSVlMQMX/rlZeeaw3v0RLcJrqhob4OIjBVSPVUJnXzl55+/L/8hvi48a77HlUgRO9Tjzhgdy/Fk0iUwZltenWM2Xzi5K+/mv1FOvHSWh/0X5SqHFcYvLVn7LohYAgYAoaAIWAItB8BSwnVfqzsSUPAEDAEDAFDwBAwBAyB9Y8AzlKcaHu20jTOSMiATjsj2xqS6+jEGYaDmXZwonvf1ziRnFmf+z7v4EAmSgNHPREGiAFTojyDfkW6uW1xWpw0SCO9eqVZIWe7f1DlEn+t0kP5JMLN3/RzqEfGKX5Ozw+TFaq3/dFgCOXEqhMJ/2KRAWFpPATqq3OqG2rDg+ONwRZkhdcGBEW6pY2po3mhOIWeSjejgpYAZA8FBzt93Fy2Y1VFQdHM10b0+fKdoZMWftZvQqw+VCa3NBijjUAaHRyWH7nveql/EJ2GXEil6ZJ4t3/0Tl/WD9tq3rA+oyrKy0dUfFg+fPnXg7dY+PnQLefPHbPr7EjfkRVlIi4gND5RlMrivJLaxvyyGhzt0xVbMU8EyLKk4/PmOqhnhg7eIjZ6yOTYZ6HcJGmeMsspuoCTnOgFrzC/RDWIDErNNY5zyAWc62gq8JvrnS3gAsFAP1l/yxGFz0wxxZqCuJBBriFIfJ4MjQQE2XkPJz9pcy537xNxcY9sX9WVL8txyRfWvEe4Zesze5M92t70aB0at5vuib6yX0g/RYQIouKsnf1lEEN8B1f+e8A8zZG9LPuEqIrOkhWBYDB42HE//PF9z77xgXzgQ08/7tD93n71JdJxdajgIK/U/2zhpnPKfJl2uJabV5BKGXXg94/6wb+efOU9dBjSnyUlFeLdRARk6lDg2J8k8We0FDLTQVHH5K232xEB6c+mf7SGTsUCOfxx3O+2zwEHp7f3y6uuvwW9jN/96tyf6TZkVnM57Ac/PO0fj7741rZK5cRFCIyTzzjnQgiW6dOmvpP+7BgxNfxGxDr9erEYhGtu/cf9EAOZ4uE8x1j5nPrmq8zlGgXc0JrIjDQhooOHVyl8okjq5Lf9+7HnqevX55z+w4+nTW3ex+pypKa6GhJvjTJq7OYTP/14Wpspunhx7pezZg4ZPnI0GHgVEenCPF567U13ZKvfrhkChoAhYAgYAoZA6whYhIWtDkPAEDAEDAFDwBAwBAyBnowAznic6mvkRHc7jdM6a174rhyUK3bM6WBOInPS3HPOcq09ZAnP4GDGAYYDGSc+p99JI5RN+Jdx4/zC0d0vfSw68S/CwvdKY61THQg6w0RY7KH7b7n1kKYIhz4WltM/KEf8aIlXvyKyYj+RFDlLZ5UPVmeOElmRJJqijeiJbDAyFogL73NtUGc7lY+zfJjM05o4Rt8PUV9EIiTLFenQJxBIfKX0UO821IRzdB0ygEiFTHIFsgJCh9PudSJl8pTaKSQh7zon4Xte9YwVOTFR1/sqmqRRvwOBYLxRPV9YmhOdI4LjC0VUFCn6gvlYLrHvvkoPNU99IFKCuolsiXBmvGxo4qXC3ol761YHyJefTjbgIIcwyRXZVKkoCy8aB4KKlESQIcwjdUIm8e8vrntkw9qwa+0ebZBaB7Ftb/0x762m63HTRXF/lgiAC/RJ6h2c/ue6/aefjBmBYyI2SOdD+jKc82/III4gBbIV9iZz83FnBsM7GREUjI/1yx5jb7MHIOHAmX1BdA3OcyJ3+A0GYIHWAH1eQ+C8o/3CCX/S6Wf/Aic00RU4zH99zk9OyqZ10N66Z8/8dMb4LZoiBjLTNRFJQT3nXfrbPxDtcMwPTzsTsedMgeoJk6dsi5P+5SefeCSTQBg8bMSo/IKCwiceeuIRUiRl9qtc+hYL5s75UsEPa/z3BgLkiYf+ffdRJ/74jHN+fdV1kDKIZ+994PcOJ7IiWzQH/SP64vc3/+2+d9945aXxioZIRaJc9oufK+AAgqu5jNl8i8m0O3DIsBHnXPKba597/OH7SfV02tkXXdpLYR2k2MrWL0gGiBQiKLLhPFQMCCRBXW1NC+KYtE9gfOQJPzr9+8ec9CMiR/5wxcXnPvPoAy10MD56/923tt9lj33ox23X/xbiLlX6DRw0BKLjAwmrt2d+n37k/nu/c8jhx/z66j/99cmH77tn6MjRY474wSk/GS5tkv/e988721OHPWMIGAKGgCFgCBgC3yBghIWtBkPAEDAEDAFDwBAwBAyBnowAjktOVuPYz0ZM4BjD4dxd6aAyscHp/KHM+zua1DntISyoh+c4zYvexhxZKoWQez2zHeonNz/t4bBtKqIJcKAP2yp2f/mIxLZuFAK44PwHKxzLXumjFhf7/cnSxTP77C7H/ygJSzsiLdSTVKCEHKeZzbb5m3mgzzjhOemP870jhXchGTiVnZ5Oq15u3PxgTmykSAZffq+6ScFIdKG0NF6VAPfuSg+1l6IfsvUW8mA72ZL66sjC5V+XxovKq+J6f2ulhqoW8SECw+kl8mOuFCjq9R2nfF+JbQ/IK6mjvrgIjRq1naf6S/SMl24IkoR1V6N35tSu9H0lLAfpewvND93HiQ9hROohhLmZUzAilz/RAMwhkSWkBGKdQgykxKm9lEsdAS/tWbAnqoG1sY/sM1lK2LmtonbRuMARC3l2q2w/GZEWzMc/ZZyGT6UPUiHlFYVImdYIEZzFkGoR1cvYUqmu0veFS0ikk1xepA6fkA6sYUg8T7ibsTG3OKrBj0gKnn3R/YQgoU+IQKNRwZ6iHx1f0e4A0z+UjmmrbXfcdc/333nj1Wsu/cXP//fck49meaxDl0gFNXzkZmPFmgUznfPPP/HIA0ef9PbPcHrjaEez4bLzzjglk9iYrAgKyIg7/nwdkTItiid0/aKEn7N1jGiDT6d/2EKYOv25W6676lINepfjf/SzczAiD66+9IKz7r3z1j9mq2/enC9nXXb+Gadc/Jvrb97nu4ce8cWn0z86/ycnHJEt5ZWyPm3x6ccfvj9n1szPjv/xmedi1ElkxE+OOWjvbLoe3IfU8NJVZesDUQxclx44a6C5IB5+101/+N1RJ532M8TCr//Nr87PJuj9+0vOO/PP/3jwyd33PeCQdMJitKIrEFRHnLs9k/zK808/zho58LCjj8d4h7Rh5512/OEvPPnIg+2pw54xBAwBQ8AQMAQMgW8Q6GhIt2FnCBgChoAhYAgYAoaAIWAIdCsCGcK6nKYmTclFss2yNPxnXeNkLKmWUs7KdXQEtzk2N0VNyiFLX9vTXsaYaMP7O7y5z6SDcovnwIUMwBlOmp7leqN3UGfO88sSVVse1Hhjcb/klwW9E8f7AymnOfXwPA7yb0rSWSZhad/XHw7stWJ+SQDtBkUbtDnGNh7gRDv9xzHdnAJF3yFjWra/ZkWeeDnzhSOaSAO0FETEJGcpPdMoCWJX5RTVKxYiMFPRIfcvnd27UeLcisDwfaRoiG1FvJACqEVR6iYnlNvYUDpoVVVJ/9W54bzo1ILSmgfzetWNFhlBFA4n8tFAwSlPlAyEBCK9XMfZT1QBURzk0If04Tpj4/tTc6YGH/zo6dDWqxf5b6erGc0TWXC17BFFWKTSy2i+mYtLZaTAek1GGqaUZoeMaIiVEAcZ9bTrp7uWqB9n6g5un9kf/6CC9qzH9Ibc9QwuzB3REkQzXCLL1CZh7rIdeIMoIF3XX2VEfvAe5AMkDXjSV9YMn7QDaYVwtPeblFqsJbAjWsbTX6Gtx2WsEQgViC5wBG9IoTnuZwtyRNe6pBDJgNO6SypTJURWkNJJwQD0PWshEgAthtbSFKEFQbqjd157GRxaFH8gENhymx12fv/t11/JJDp4EK2ICmlk4MBvrX3qEFWzg+QY8tCmyIziyPZeKBQOK5NVYWv1BoOh0BszF1U/ePddt117xUXn7K60U7379OtPVMk7b7zyYrZoEK8d+kwqrWVLFqH5k7UQvfH1V7O+yCYY3t65y5zrAYOGDBs5Ztzmr77wzBPtrYPnxkmjRNIZ/ebM/uJzCJ2OvGvPGgKGgCFgCBgChsA3CFiEha0GQ8AQMAQMAUPAEDAEDIGejADpS3COE2mQrXhpcfDCd5lzcW2ApJ8cb69zOMtzLU6Cp5EVNE0qHE6sM3aEkn2QFUr95AQiSccfdL7M65UskTZFjWgKBJ1xAmNEWXAKHoc4jvJ66TEEY42BqkTM37uhOtIVZAX9o34KYwBzHPhYW2QF7+C45nQ/AtwQAqQgckRMOL5AYlQoEnMgVRpqQ/P6jFheWzp45dZDJ8//euXC4moJc/9/9t4Dzq6ruve/vUwvGnWrWMVFlmzJvWFTTQskIRAICS8QAgkkhCSEkPJC2gsJvJcQWgiQAH9CaKGHbuKCe5Mly5ItybJ6m9H0ub38f9+rs8d3ru5o2p2i0dqfz+K2c/bZ+7vPMZr122utayReXJnoqzudxkqmqIjTA9F7FQmP9hxuOaX6FC2q13Fp79HmRxau6douAWO/+ocH0RVEOdyv8xaLyVZFZdwRiWcaFWXB30WMB36MDWGBdE+bZXWxJmXPyvgpLE0tDSISyhtrRQH2gNbR76WFwgGPY5iUWNSu+C+vX75n0GeW767odIyPOPH/QfZ5GaIKTn/WoDBeEc31793PONEHdS5iDuIDu8Kpm4KK9jwZ9xaMqv39iPDCtV/jzRcxiCLwCBDcw0RDIF4QLUENA4qAk1qL+5wIKfrmnkI44jjY4+yFPcezZp+Q8YwTycJYhwuWj/cZ1DkTarUUK7gwIsLZxAqO6e7q5D4ate3e+QTRXVUbjv9HH7iHKJ+qjZRUYwGgj60P34/ANu5GXYyziSDUmEDU2PH4Iw/BtLL2xtkuNJ4xP/3kdv4/YEqtcq2PKgcVNtFOdz3x+LhqXky0XzveCBgBI2AEjMD5RsAEi/NtxW2+RsAIGAEjYASMgBE4twjgCMXpSb76UuHWsobjEicnTvNhB+Z4p8fO8gmkcxpvt7U4Dscs0SREHlDUWbuz5a3Vv9xD4aIvGPQ9G60vXhxv8tX5A/6DEi525DKh/arfsF4ZjUgRdIVqNdTnssFUz5GW7XLyL9erLz1UHgwx4WHiSGbnfLkowbo44QUn/Hiit5/2jmtR5AO7phcomiIVjuRTqjFxsnlRvz/WmO6ONqRzrUv7lgQj+cU6bkHbBb2pUCTfluiLJ7OZUDwSz/okxPiyyYgvn1MdjoKSOckyyXDq2FOLQxItOpoWDr5In5dLnNinUXarH3ZLX6jPbaqNsU2CRUIpp14nVo3BcKFVNSyIFCCV0yoZUSs47FXowx9I9jfkUoPFNp+/0FGl6Ac7/18kow6By92PIPEfsltlOPT5TPqwCYOvPMHrg+geUiI5IY+USf9IgempXMCrdcF4EQYO6BoU92bdGfiNMiJMnGDlLoXIwfHrZIgWrPEjMiJoLpe5qArSEbnnlL9D6ZdUPtSdoH/EIiKquD4cSW2E6IPwUeI3lbnZubND4OINmxCefERszM4I7KpGwAgYASNgBIzAuUbABItzbcVsvEbACBgBI2AEjIAROL8IkD4Gh2W1NCbkvad+wTbP0TomGTlgXTFrRIGQPuMExVFa7nyfcFqdMS88xgHalT98hHbpIwLg6P2F0peSAYiuUMWJUv0KpYSKR+t82Xwu1Nx7vOECOd6Lqk1xa+OCocX+QCGXGoj1x5uTvoGuhv6jTy4OKrogllHdionWqwgET4cxlMQAn79X/8Mu/vJW7rgeLV1Q+fHs3MeZfZlMAkHxu40dg6lF605mNfYnNL5OCS6FutbEsnAs26z6EyHNnV344VA419K0qL9P3x/W3FoViXFU4sU1g10NYZ23TXMuSJxYp7F2MNdsOpQXl8fE5RKJE7cvWX/yqM59EfUslFoqL/HmJYFAYWnficbwoSeWHmhZ2rez/YKebdGGzO0SMHC07+e+U39BHRs5/MSalmh9r6Jchu7PpRNbioUzfOfciy5VVtG7H4/q/sLpPuUcXKPcPgg+pFyiIebdrOtR46FUz6UWYpz6YF271C/PCHUlKsUKLoVQs1VGtAdCAwIEYiJCBccTZYLTmu/Y5c/zTL0NmFF7gsgV1pnICleE3ouhmXiKq9M4rM0VAkqTtIW0TgeffYa1tmYEjIARMAJGwAgYgTEJmGAxJiI7wAgYASNgBIyAETACRmCWCeC8HG33/nh29ZeG74kVOKPZCU64AY5VnKaHZThQES1mtZFSSANAnsDZS47/QX3REIkXfQW5obMp/6FMwv9Yoi8STva1bM7n/RtVkyKmdEhxpU3qHeqpiwycbMjWtyeIKgjKAV8c6q7LkzpJEQZH9IrzeLQGZ3a3xxRt4FMdCBWkzgaVSqqrUPBnVD/ibGzG/LtCfXZIPLlU47hA42iua079Qn3b0AJFVhzSdaLR+kynxIIuf7C4TMfg6MYhT7qlRq1+h6IgttW3JYaWhE4eVX2L4uL1J/dIqAjp/BMSKLp337PmiOa+TH3fVMwFCgOnGvL+U8XNvceaXq76GP+0bMOx/ep3g3g2x+rTGxSREq9vTaSPPbVoRf/JxuC+h1YeUDFu/8bbdh3Q98fENfP0PWuaEj11y9JD8Q2xxkBLrLFte9/x/YpoSV1WpgARYUC0wxn3ohz+oxWqrsV9hnMfEQgxAIf/y71x4BhGaKhJAepxDJRx7JQRjUGUCveve2Z55bc7vH5gxHNWElVo4xUbxzEOO2QOErh00+arKKpdra7GHByuDckIGAEjYASMgBGYAwTG/MNiDozRhmAEjIARMAJGwAgYASNw/hJgdzrpYkgVU9lwlD4gI29/KX8/B5wl7Q5FlSkojFOe1DkUGKYQMju+SU0zk07e0VYUhy5O3vtlFFIuucGjDUVfWBJLvLl4f6wx6D/2VHvDUE9rk+o+1Cld1HLVa1AURiEtUWC56jFkUv1R/U94QKmTuvUdwkM+mwodLOZHCBak2VoiJz41JLpkCCRFRSb4iK6QQ78Ya0j3Kl3TfqVfCiX7o4pcwC8+ZqP+APUiSCNFuqQmUlpJBMg3LBgKRmLZU30nG+s0zoZ4U2pQ10pF6jKRcDS7UXPl75ONMtad2gUuAqZP41wmMaOxviUxIFGC3fhtShOV0HgjSiHVsnjdyaeSvXFNPJjT72FRvFkzi0p4WH30qUWrOlQTI1qfXhIIFdZwPYkwxZal/cELNh31qSj5+mwq9upMwV946GubvyVeJ1Xou0N9E1WgsZC+qhgRVKWo8l8moyaBA8F9VapNoUiZmUxbxLXI349QgcBzk4yUVkQjdeuZyNYiyqLs2eJZ45lD5CtvPJs8o0HvesNihHcQ45x1MXDMu9YOqDkBinhTKPw/PvOxf6p559ahETACRsAIGAEjMG8JmGAxb5fWJmYEjIARMAJGwAgYgXlBAGcn/2Zlp31lw3FKUd4nZMOCRbVZy+lKHzjPyZuPWOFy55PmqF2GAxwHfqWzdaYhIlgw15EFJ+Qbb2gv+JqXFJf4itHeRF9D3WBPnZI1+ZoUYeAKUC9HaGhoS0QSfbEFEiv88cZUQoWl746F08wxXJEa6oCOlwM/75MwEQ+FVXo2G2xSaqVSzYx8JpTNpYMnQtF8d2owcmm4Lqt6EUFFeoC6anNpoShwzUEUW8bBvU2iydKmRQN1bct79+taBxXRsFviQWtTx2AoFMsOKMXTIokVFI8mxRHnkl6JNeM9aYZWy3CMd+q4TokXfNcW9Of7Nf9SwqzlG4/WJftjnzrypBDl/RR9Jmd+UMeeUnTIJRIfEEEQqOokVvQX84EGnRusa0n6JXi0i9Ni1QJpldCxRBEriC6XyIiQ6NN3Ulri3G89SgelYudFImBco6D27XwoK7pdnVDtvyUVE88I9wsC3EUyxs79XasGX9aCZ61SrOAa3K/8PpNiTa3mZv1MI4F1F2/YGIvH63ZsfeTBabyMdW0EjIARMAJGwAjMMwImWMyzBbXpGAEjYASMgBEwAkZgnhFwW/rLHcTlUyR3/7dlREmM2sjFL9GCnef0h2OX/ihYjBOclD4H5wg3nOo4hXH6P9ckWBRyfhWZ9g2kBoKPBsKxzarx0IDAkE9oSoqSUOSCT2mVsq3LesNNiwP1SntE/QnqQBRUx2Ggc9+ChyRGbFKdiCV0rIiKeKwp2RsKFVokGtTXNab6VdA6E6kLRdKDkaQKWvekBmPPRgqZQ6or0RaO545lE+FeCRYvHoWV+9sCYcg1BKIdvkBxj8ayQsJEVoW0040LB+6XsLKhvn1olYQVFQ8vIiJxPqmVOB/hBgZ8d5WMYt8cQ9QGIkKsdJzmplciZhYqnVPdhVcfvKP7UOudql0RV5RFqZ6DXrenE5GG43s7Uqu3HNytc9p0bIsCLPzi4VcEhmqDFA9pHBdK2LhU52BELhA5wTUVvuJXhIevN5/LDvoDgfqKXEs48oluICqG1GIINzPVEOselVEQGzaIbggMTsCrRVooRDwiOCqL3rs5umdzXOE3MwXGrjP7BDZuvooaQ74dW63g9uyvho3ACBgBI2AEjMC5Q8AEi3NnrWykRsAIGAEjYASMgBE4XwmQbobd99UakQMLZERIjOUoZvc+O/Nx2NOnO486ANRLmCs7xHHOj0iBlUn5fUM98kKHfIsWrC4sL+SHVIOhsFhREb7+zgZFFAR8rct7s3UtibCiFoqIERII0oqICMgJv1aCRVzRBNco0qFYKAZL5Rd0zOX1zalDoXg2RFXtxsUDpxSFkFMdiCWKNMj5irlIuC6zXO+H4pFUdyEbSBYKwVdP4ibcKHFlh9I3PaJUTD3RukxxzbX7V+r6rRIKWvTKerAuONwRkXCO83dK5W5+1gcBhFcKPeNIR+DhXISFhnA8e3HH6lP7lOLpqKIsEKZKf+9oDisPPLa8sGBF93eVluoZzfeGfDbUrkiKFrHIt6/sLkq82OP3x1ZI4GAMLvLGTbdNokVvKBorhiJR9ZcRw+HbjSLirBlixYzdQ6RfkgiHUPce2a+UcSC1F/e37piaNBjzrPCsVWs8m1zPmhEYQWDDFVdec+zwoQOnuk4iClszAkbACBgBI2AEjMC4CJhgMS5MdpARMAJGwAgYASNgBIzALBHAKU6gRxQAACAASURBVE1kRLVUNAwJRyk78p+VnVWwkIN3UA7e7+s4imyTU58C3LziTCMFUS12o08VE/MljRJRAydlCxlVqeC2vlEKp3BjR9Kf6M0+qYiHaLQuHQpFc81NCwdyqrsQUGHqnFIu5SVSPJvPBTq7D8u/X/RLdAgulCk4oDiYL56OUFBERmesOZlS7YhDOqazmAsqXVKxSbUvehSFkNT59cFc8LJsMrxo8FT9YUUibJYIMpn5ZXTeMoklcO6RQFEv8YKd1zj3EYvYoY/ggIMd5z+CAcWbibCghgRRA6wvNS34DjGBV6IxEDuu8465Q+mfFqoYd/eRnYtPKBKE4uo42wti2KH6G23bf3TJ3qtf8/iTiqZoDoZzy6N1vgsk0jQNdDbEJOockliBEIJzfk3ZRBmnIhb8sUAo3KfUUE8HwsmL8ukRtxvnsV4zeg/pns7rnn5G1/2kx4VngecFntR2OVtNl7IpnvUtDEu1SEY5imeTa852OrXxzseOmyECV1x57Q1PbH3Y0kHNEG+7jBEwAkbACBiB+ULABIv5spI2DyNgBIyAETACRsAIzE8COIsPyBAZ2DFf2XbpCxz842py8J6SE5fUPa42BqmFBmtRnHhcAxjlINU+KP+FaBGiDHDWl6IhsoqwKMg/HooWe5o6co3hWP9uRQ3IgexvVRqoYn1rMqq0UAMqOj0gMSBeyPv3HHpi2T4V2l7TvGjg6FBPfJWiCfwSIYadzhImisn+eDIfCzYqhVJQERiDjR1D8WhDRtcLN0vgiJOYSed0FAajHYWiv0/9jkxVNb5JdyoRVKrrQNt61dB4cOWWQ10SVzZ4p8Kf9EXUqHBpn6i/gCECULyb9cUpjwCB4xwHOYIOIgbn8BmhAF7dqklx1drrn93xzAOrD2j+gxIhfknfX6sjBsVn+VN3rntw4227uiXe3CoP+9PJgVix91hTYyYZIRUU6Z0QsohScK1UtEMoAuor5A8ELxIsnwJYygtvU0OC6A/EoJkWLUh3RnQHEUTwROypdZFr1oBn7RVlXNxbnk2e0RmLLqkyBvtqjhFoaWtfsHLNuou++oXP/MscG5oNxwgYASNgBIyAEZjjBEywmOMLZMMzAkbACBgBI2AEjMB5TgDHKzvXqUfwpioscHTjhB/31n+JEziVaURVsJt/Sk3O4tK1ayh6sKN9pwwnfWmnP2KFUhz5ug8HE6mB/CmlPdqkmgqXq3h0KDUQOyBxIRJvSqWDC4aKctLvUHqj1rblPb+gyAa/oi0aESvkmFdNi+cKZqu/hYmeeFKxCkWJH6SBCoYiuUbVd2hSpIIvUpcNKfqgX5EVTbjg5azHif+0jMLO42msHcKDclYphkNpqhoWDL5JkRZ36vMBrdhL9ds1Mhz8CDREWrBTHzGC70h3tE9GyiGiKPid9E+sG0IF49kj4x7gHMb1MwkvrYvWdl0w2NWQObZ74RrNH9EDR/5BzcF3ct+C1fd/6ap7V2059LAiKwZO7O1YKD4bJcaQFuwWGczLne+MJVksFvbk0kMtKrq9QKavWPaSNoEznw9ENcyoWMHFvVYa4zSNgbnxjMG5WuPZ5BmttUgyyuXs63OBwOarr7/Jr/bYg/fdfS6M18ZoBIyAETACRsAIzB0CJljMnbWwkRgBI2AEjIARMAJGwAicSYB/r+JAJlVQtUZaIJy1s+IslViBuICRmofX7BSFCzzhOPlpI1LwEGkx2BXIJ6WP6H2DIgTqA0FfQkLFPgkM6xRh0abXnlwguCQcy12iFEiR3mPNqWR/rK7/ZKNEj+fECjrHeS9nfp9SIYUkclCkOhkIxVaEI3kFERR9wVA+mR6MSqwoXY9GUeXFE7hJOb5U4Bt/fmogukv9tSi91MpYY/ouCRcv0A8IFQgQiBPs1Eeg4D3nISAQVUPkBKIAKaNc0XSiKjiOdae2AscgYPD+qNJk+VduPkRkR6T7YOtWCTgDmh+pnlol4rx4qLtu45O3X0SEBjO7REbkCNf/ioyUU0RL0B/Oeoz3iwUmW1R+rkJeJT48KPqeiJgJiWY6vqZN9xz9TZdYAmP65lmr1ng2eUZZL2tGoERg87U33Dw40N+3Z9cO0r5ZMwJGwAgYASNgBIzAuAmYYDFuVHagETACRsAIGAEjYASMwCwQwKGNo3m0CAp278547QA4eJEVjA8lgJRAjBHBYazi32fDiGMYB/5KGSl+SIE03NJD/vbDO+LHmxb5lsebM8cVDSHRotDmDxZ7FT2xIDUYXaC0S4gRxb5jTaGTzyxIy0H/uOpQ3KKIDCc8uP72KjJjTbEQS6jeQ6OOiw1lgz7Vd/CFozkJDDGllgpUnsM8ST9ULlwQ9YBY4xz7Z8wP377EkeVKC5XI5wNNrcv6mjXuJ3UgAgQO/7u885k34gP9L5KprkYpRRN/t3Af0HjPeQgLe2VEFvCe6xN5kZNwk1eEyEHVs6hXTY+lx/d0HBOXTRJt1npFtYnMQKhg/ZgTERqsG0KI+27kPaeK3KphUfAHVbS85L8f1gcQMxA4EEuYy3QJB970Z/yF+fCM8ay9q8rV4cTawM2aESgReHLrow/t2r710YKaITECRsAIGAEjYASMwEQImGAxEVp2rBEwAkbACBgBI2AEjMBME6CQL87l+2SbKy6OI5VUPzREg9lwjHHN04WdTzu8Q16h4wmJFo/e8x/DU1M9C+Z8UEax2rXlc/b7g6nuQ4sv3Xt/pLm+NRNauKazVdEU0Xhz8oiiIpQOKlzXfaSloJoMgVwqnJRI0KlURxeF6zJKB+X35TMhRQcMixANeq+C2IGO4WCBQtCXUiSGoi5KERjPBREMj4J5kpqpvI1WjLniMH8j0R6FA207O1Z15xesOoUTnKgGl96JnfykHcLxzdqyY99FUCBckL6L6yN0tHm2TK9bZQgWNKIw+BunJRAqJFSMvF/CyEbZwqHu+mjP0eaQhItGzWuVjsHJTropeBM9wLUYC3bG30mKqEjnUolwPpNSeq4Ry7tfxz8km49iBUxdaA7PGutSKR7ybPKMWtFt7ya0F5/vR9/9OtFK1oyAETACRsAIGAEjMGECJlhMGJmdYASMgBEwAkbACBgBIzCDBPAM47hml321dpu+xLnPTvsZbaR+kjiBAxeHriv6jDMXpznpiibbnEjzU3VwvezCUkcKkQgEw8/PZ/0L+k7UZwqF8IXRhnS+ZUlfRAWjM6Fw7pRqMiw+unPxkASHiAQHhIUNqulQaFveq3MLPqVjOqLUTMF8NhRUMe1dOqZZznuOG94dr+9Oqb4F0QLVmitGzboQlYDo0C27cqzJlsSPgj+nKJDeJ3+6fvclz9/zeMvi/iXhePalkkY6ij7/LkVGbPPmS8QC6aBIDcW1ECpcjQaiLxAHXEQHQgZjYMwIEERfJNXXFYoWuaR58UBzXXOqa6in7p6BrvqYokpWqC4HUSyu7gTrRb0QRJD1MiIuKlsC9Ua1K6KnU0GdEfADB2qjDBe2GIvHOfY7kT48a9UazybP6IREunNs/jZcI2AEjIARMAJGwAgYgRkiYILFDIG2yxgBI2AEjIARMAJGwAhMigBiAA5qUvVUNpzDOEk7ZbMRXcF4XO0MogxwlCNU4Mgf0SRs4IBHGCCd0vBOdK/2wIhjFW1RUJQFIgw72okmOC1YMEnqJ+QyF+ZSvpSKSreq9kS3HPHPRmLZlNzoiZ7DLQslCCxRNEUQfUMiRbGpYzCzaG1nv5z3eaVEGlTR6SHVdigm+2J7+0407ZOIcEQ++BUSKpgD4xxPPRD+jsCYE9EP42q6RlTSjl8pqhbvvW/1nsUXncy1LO7b1dgxSBHxC+XuT6p2RlYFul1/jMUxRZSgKDfjZM0vlhHdMiRDtECwcPcJIgTfh9VfKNBQUFUO35CEirAKiz9FPQ+NBZGB/PoU/36ejPuJNaxUIxA3hnTCYD6XXYhwUUqv9dyMic7guoxlvqWDYpY8W/DmWauWmo2584zC3JoRMAJGwAgYASNgBIyAEZgSARMspoTPTjYCRsAIGAEjYASMgBGYZgI4SdnVT22Das3tah/+zUvJNM3DOt29F2WBAEFRaJzViBUjHP4aD6LLKhkpiKjP8Lh3LHUw6KPaWJ2ocaj8R39AXfn99RIu6gsik+qPt5UKYxNx4PftV2REWI74EbUEFGkwUNeS3C/xIqWUUeGO1ad6g5H8CTnti6op0am0UV8a7K6L959oXKAUUb+pvkakoRoDJPNx7RG9oS5EZcqoyi5eoTFen+iNP3Ng6/Knehc3HVS9iZ6mjoGL87ngcdXP2FPXnHxEtSceqGtN3KCTEW6oZ0G/OMVJP3RAtkGGs5x0TK/0LoJznZoaRARwPKJFjxhEw9Fssn1Fz9HBU3UJcWgRK4Sg58twtvN3Ees2sjL56U4VrVL05TKpk9lU4sKKgtv8zj3KGqQlNs1HwYI5IlTwrFVrPJs8oxZhMQog+9oIGAEjYASMgBEwAkZg/ARMsBg/KzvSCBgBI2AEjIARMAJGYOYJ4LjHWVrNkcxo2GU/2m8zMloJDnkJDzjKS5EViBjlF9bngvc7dRbYhb9FtsMdP4poQR8456nPcLqVUhLlfflsSnUockQU1JGdqJgPuILUI/5tz+GKVOiXOJEOhfMdSr3UEKnLDMh5n1S9C5zMXS1L++oVjeFXtEX/U3etC6nGw08pvq3fnBOfK1P8m3Hz/Wh/P+Dsv2qcwIliWCTRok5iSUPvkZYjGtPCnkMtCCWRQsG/O1qX6VtxxZFLwvFMLBTNp/Q7YyBlEymfmmUrICKjrzVl4+JeKKWEkpHaid9OyA4qNVbdmuue7dr9szX3DHQ2ImYgajAv1s1FjFQt7q6IimgoEisEw+H9uXRi1em0UKXWJSNqhhRVRGLM1wZXnrVqjd/gZjUs5uvq27yMgBEwAkbACBgBIzCDBEywmEHYdikjYASMgBEwAkbACBiBCRNwNSIozryxytl870SNCXdeqxMqRQqJEP6K7/bpWhfJ1slulpH3/14ZzvJq6az4DlGC+f9Y9hLGimCRy6R9cprXhcJRRUpEcc67iAacxkRX4Djn3/kqeZEnoqIooaJV4gXpnnD2E52Ao/1pCQFN/mDxCkVg7LjsJU/tP7F3weeeeXDVjyQk3KTfX+X194Bef9HrsxoyhBWuy1jGajj22amPIEKqp5hqabxZr3kJGA2xptQFze1DQyqW3aKIkI7+zsZkvDF1b7w51a2xUicB4YKxwNEJVQgPsHKNz/wGW4x75L8lOmRDEVUZT0b2ShRZ5Y23PDKgqlih4yT9gD7XmM9mVhVy0maeEyxgTfou1gnm89Fp78QIOFZrfO/quIxyiH1tBIyAETACRsAIGAEjYATGR8AEi/FxsqOMgBEwAkbACBgBI2AEZocAjnsc1exir9ae1pc44XGWc+yspeRBpND1cdwjIBB1wViGiMDQKymjvi1bLSPSAic37xn7Y7IRdS+8OhY49PmNFEdXy1pV9JnCz75cKukr1jeThqg8uoS+EAOc8zilNEjd8q13ykGfDZ4WLIgooC/SKiFEMNZGiRk3RuvTWy7YePROiRzPPH3Xug4JCUQoUJ/iMo+tXqo2xBciGsbTSOFESixSSREtAZtS7QeNMRWrTxcaFwyuyyTCIdXjCMSbk9mG9kT3kobjDweDRdJePapjX1E2b8QS6loQRQFv+NMvdSWoeUEkCf1v0nwe7dzXPjjUGye9FOPgnmmUnS0ygt9yxWJhKJ0YWJFNDiq6ZYQmgfCzX0bR9/HU/hgPo1k/hqgfr7m6HtxbPGvVGs8mz+hs1ZGZdV42ACNgBIyAETACRsAIGIHaETDBonYsrScjYASMgBEwAkbACBiB2hPACYpTmvoIOPhvrbgEkQfsuscBf0ax69oP56w98m9rnOGkIWLM5PTvl/OXHejMA+c342S8v+bNBwf7Zh3zBQkbCBTljfOflSEYkI6p1Ir5rC+bTijKIhkIRc+od00haQSLaDBUONG+sifQsrhfoRZF9+9+nOpEI1BP41ZvvK5wdq+Ei8GFF54KH9h6QW+iJ55V1APz4VjXnMDAZ/pyURUu0oBUTWMV4SaqgbXiOMQEml9yQ7j/ZGNvNhNqVmHsXGogFtC3YaW8urypo/5gw4LBjObBOU4YIGoFRlfIviz7ruxNMgQU0ktRvwKjwPZS9Xfs0I6laUWPvFhfEWWCqIHggDMesaNahAXrk1V0RVdmqK9RRbe9Q71Rn67dgBAEhzHFsjIhwHXgBCfOPeP88vomFedyHuwYHyxZl8pUZMODnOIb5ojIVYryqWh36jPPJve7CRZTBG2nGwEjYASMgBEwAkbACMxyvl9bACNgBIyAETACRsAIGAEjUEkAJ22ZlaIUZPfIviCjCLVzWBO1QAQC5hzfpe6qOIZnAjSiAo5rnOhEEOAA5xWHr2s4dXGSb5N1ytidjiBwgca8RDbs7CfKQt8TMYHgsdN1UFS3/qD0B+U4Kqul4H5GMFiodEqZ1uW9JxZe2NUVbUj3Kp2SEyzYCQ9DPuPUR5CAMVEKOPqvUFTGS9fduO9wIFz4uj6Twsk1eCO2EB1CREN5CiiiMfh8THa2tEhcl2LXiAXOwc4rKaFCuUywfqCzoU7WVMj7uwa76k+prkZU0RErNd3NOo4i2aw14g7cSA0FX8aOQ53QAMYMe0SUPvV7JDUQ7eva37ZShb5b8tkgqa7eJeOVCIuzNjFO5LPZrlw61ViWCsqdw1ojEk1ULHORC0R6uALhE6nFAm/mzD1HbQ9eR0tpNdYUR/xe5dmBt3vOuAdoPIPcRzyTPJtEEo0p2ExoIHawETACRsAIGAEjYASMwHlJYCL/KD4vAdmkjYARMAJGwAgYASNgBGaWAA7TMsMJi+Fcf6OMdErOUY6z990yIi/YaT7bDYEB5y4Oe5zoOKJLrXynvD7i5L5d9k/eK8dfKvt52Rs092aZExhwuu+W/Ux22llcLPgK2YyP9ETFPF2d0UISLNLBUP5YIFT4oaISSOWDMIKTmfHh5Kd/HPvlBaP5PS3aA61Le8MNrQkEFcQV1/jbAUHFFfkuvzAOc9Iv4TxHNBhttz1ObUSCVTLmjaOf9WVcSr3k36+i34oeCfvSg7Hl6aFIWzYVbkgOxNbpNSix4T4dx7gQTjgX4YLd/RSEhjnRIrxyP7TLwpJFgoocyQ6eqo/rfEQP59hnrDAl4mQ0Z3+hWMjtHuo5ESzkqmaO+qnOfZLxSGCaiMOe+S6TDd8j3rjH8/cZx8AbjqwF9z/zH47C0ftaNlhyDZ41njkazyDPIs8kz6bfS4lWy+taX0bACBgBI2AEjIARMALnIQFLCXUeLrpN2QgYASNgBIyAETACc5lAhXO/KEcoXnkcy664dOXwcaZulbG7fyJO41pjoI4DznocvEQQ4FDnu0yVItw49Hv1/UPeILbo9VqOleH4T+i3b+j1mbe+4R046O+S4WB/E1EVFN/OphK+vJzogdBwoINLO6XaDf7dqv/QJYf/bgkXh+vbEvTPgUtkOLxx9CNGkHLK1bVwhb6HguHCohVXHH706bvXPq2ohzUSEqKK0lD9hgARGqwD82SHf3mjH9Ijna0hDBAdwJryt0i5UMD1ERn2aYrMVTU6/MqAFcj0HGptqmtKJetaEw2qsfHU6d9KoghzcWmRiPxgnvRPxAh979eYt0sEWSbBwi/B4pqKwSEYIIJcUmU+HNqZTSYeyiYGfvW5OtvDPXxT7yiIzppNtH4F4yYVFSID3Ih04X7Z771WDLPqR86jH54N5gwP5lzLZ4D+GCfPWLXGvcD1cxZhMZ4ls2OMgBEwAkbACBgBI2AExiJggsVYhOx3I2AEjIARMAJGwAgYgdkmgCOXlEikpcGpX9lIE4QDndRJw9WCidKoED+mdR66VkHXxFGO45gIAJzJOHSTOHPdDnTvPc5mFz2yXe8REFbJcNS/wOtjg14/ftV1Wx555IHHqNeACIItQ7DIK8qioJoKRFv4g8FBpYg67PcHiFpoUAqlpr7jTUHVbXheQ/vQgVWth3ISHGBDei2c2xy3Q7Zftl6G05k0T4gYcR0bWLS2c1Uomnvy2FOLcFh3ZJLhI4NdDY+o7zX5XLBNbvHbpgAUMea1svJUXvAiagAe3RrDKxUZUacokVO+QPFgMJJXJqwCKbaINiH1FXPAYM68EHpgz1wwIi/y6oPxIyrAEAHpCRl1QYjEcEIDXCsFGPHN3Z4a7F0uhUjCxhk6AGtGH+MtOF6Oi3ET2cGYmTd9jCbIlZ/HeydM8Yqxbgg9U25V0kERUfEiGc9YtcYzybM50ZRYUx6rdWAEjIARMAJGwAgYASMwPwmYYDE/19VmZQSMgBEwAkbACBiB+USgFI0g+7bst6tMDEc8O+dJs8Tu+1kr/isxIuuJFvw7m93zjCWm75bqFcf5Mb3HmU6kAzUYiEjAac/xn5BtklFEGkfxTbI/+c3fefOfSrDAKU3B7gdkrxmOskgOyZdeVJRFKOD3+7eFYvUxvdbLt54Y6q5fGQgU22VtijDY7w8ql9RpYYTd/DjMiS7AYQ7bO2WIAYwHBzqO/jXtK7rrWpf2DSoyoSBrTA1FWnqPNn/l8I6lN6QHI7cp8kKHTqq9Umc5BYAxMV8+EznxQokVx3T9YsOCoVLRcIknJ2ONqUX6vl3XTOsVMYKx4yhHsMBhT1okWFJTASGBeS6hH/V8SOcRiYEwwLxdXRGiTigoXV6PY3hCimBpVCoozbPqHBFW7pb1TjAdFJ2xFkSrcE8wf8bthI/xREkwb0Qx5oFYw7nM4Yyq4FVHPr4vuQ+Wy3i2hoXAilN5Jrl/Zu2ZG99U7CgjYASMgBEwAkbACBiBc4WACRbnykrZOI2AETACRsAIGAEjcJ4S8CIScLCTGun9sr8qQ8EudWo/sOse5y1O2xnd7e1FTrgiykRIuNRGv6z3iA844REoLqpYQiJCKGyNCPGMDKfzf8t+KLtBxs721mAwePmLXvb8793+gzse1WecyK9x/aSH+pUWKutrWLCkrlgovERFoU8p0mKtnPOnsunQk6r94IvUZVbpM5ETMHRCCU57HPoUTib64Je8PnH+cwwCQkiFrgtKwRSUSRnx5WJNqZvqmpP3Ni/uf2jb9zZ8KpcJ/YaOw9nu0jNVTPGsH1lPogqoi8G8XP0GCQv+lcoG1ReJZ7KK8mhJ9MVzSmvVr5iUmGSXoD9YEniQEXD6U0PBFTyHNfcEznzW5GA2FXqs91jzEkWbXKXP1SIpqooVEoUy/kBgoyJZosWS1jOifVmffuQxnWg6KDpi7IyT+iKsA5EliAKs0XhSOpFSizVFhIGFSz9WS+EALjxTRLPc7I23vIA8zyJrmLd0UJW3h302AkbACBgBI2AEjIARmCwBEywmS87OMwJGwAgYASNgBIyAEZhJAjhyiZ6g5gIOeyIRaM6BSpofjnFplkpO31qlhapIlePqMOCoZ5c/qZtw3JI2hwgQUg9dKRvr39oUXcZpjUhwUnZYjl/mwLgf1wtRFQgKR1/92p8LSrDAob1YphoVvrYCBbelKARVwyKfz/oisQZSGrm0Rq2KqgjI0X/y2O6FT0Yb0vmWJf0LVYybKApEFdJCEZWAWIFjmkLcXNulOSL6A+c3c8Ap3imyCb+vGIrWZ25T1MJdDe2JfX3HG49IDCF6ZKy5Mq3yhjiBk51r07+rUeKFbBQT4WguH29KDYQiuZjSUC1LJyLZeGMqGwgVcZ7j5EfsgD3XJ8rApYgiIgBx56hc/w/m0qEWpbMSrgCCEJwPeNfmHkHsqNqUdiul2hVDhWxV/YtrrfL6m6xIwPWZNxeg+DmvVauojzZEfe/qZ9DXeISO0aZbelbKmnuOmCfPFszLxQqiSz7qjbl0z1ozAkbACBgBI2AEjIARMAK1IDDRPyxqcU3rwwgYASNgBIyAETACRsAITIYAAgEOdxz8lY1URjit2WmPE3dKztsq/XNt0vfg7F8lu0CGwxynLY16ENRFoBG9MFpDbPhX73jGShornNVZt0tdjmOc+YyfQuI4w9vi8Riv7KinDTuOES2ymaSvkNEm/6hOkYDhtdPFqJUKqftQa30mERna9LKd+xQdgQhCzQqXdgjHP6ILogFiBdECToBw4kX5nHbrwyalmQrFm5Jb+0409usaHD/RxtwRRRBOYOsiDmDK+vWGY9lTscZ0XKJFk8SLNRJbOpUK6qQM9inZfm/cXJ95YIwZngghjUWf/9L0UPSBE3s7qLnxen0HO0QLroNYdGYrFg8ph1RCkRXxRG9XoFA4Q4/gPuP6e2U9E0kHVaWmCvNmvthZ2yj1WKYsVIxyUe4P1oi5ViukzjPIs0iEy0RElrGmab8bASNgBIyAETACRsAInOcETLA4z28Am74RMAJGwAgYASNgBM4RAjhFcZzidCZ9TmX7FX2Bo/pLMnZ/j+kArjbvsl3mOGxx+pMaCZGC+ghvleGkvV5WXiyarpxY4br9pt4gMFCUmHRVjBknOSmJEA1wluNsLtUcwBlddm0ED673Cq8zoizYfY/nnLk9IiO9EQ7lUi+Z5KDqWARlka5gOJpRHQtYsWX+xYq0SKeHIp/PpsKpYlPqSjn8ieygVXJkTogI7m+EapzrFFHxbUUsyJkfj+ra+3X8ahms3K58r/sxX8p37CNcYLQIURtK5dQtC0gmigbCeb9Eiy5dAQc6a0AECqmr1siIFGGXPxEU1PmgoDcRI8rk5O8e6q7zq/7GNZF4NiIOd3p1N6jNwLpWtqFCIT+gYubJoe4TF+XSZ9TT5voflrEOzH2+Ouu5B4g+eYOMZ6uycW/wLP6LDCbWjIARMAJGwAgYASNgBIxATQiYYFETjNaJETACRsAIGAEjYASMwDQTwFnPrnZECWo+4LCvbDjcEQVcLYRxD6lCqEAIwFlLGhwc37fINo/RGcIE46KGwrdkP5XhzGYsOHTdrlA4SgAAIABJREFUTviqkR9l10cgoSYHhaCJhGDO90rQSF1506/S18MyRBlXLDqg1EVKCxXyhSJxCRZhBAfXqIFBe1hixSsPbl329MW37j2oyAXGuUVGeqnyRv9OzOD7anUpiFRYpd+agpF8t5z/P9H7S2VEPdT0b4tsKnJZ9+HWo/GmdDFSl00V8v58IOhvllSEs5waHwg78Dkoe0hGOiyEGtYKMQIR49qWZX0vTA1Fw5lEeOjUwbZEaiB6ob5nrhTu5pU1KzXVAenMJAZ2DHYeuSWfzaJ4jCSktdAX1McgNdl0RTdUXnM2PsOFZ6lSmHNj4R7iWUzp3pxsSqzZmJdd0wgYASNgBIyAETACRmCOE6jpHxVzfK42PCNgBIyAETACRsAIGIFzmwBRBggDo+1qJ8rhv2QUcSbCYiKOVBdNgeP9Etnvy3CKn60hSiAeEAGxU0bkBP3kXC2K8eL2BAucwy+WbZRR24A6DP8pI5qARgQD/34n9RFCSkAedR9poYgEIMoiHK8vBEORSsFmiVzr67Pp8BLVcfhhqOjfpigL6hK8UEaEgqt7gVCDEVbgCmFXTqFOo7hVXx6ra0k2959o2pPLBHHcw5pXxsh7l5uKuiM4+HF+IyI4QQQRh+9GbRIojik6YmvX/rYWTTOiaIsh1eHYpwLgCC2ciyCB6IBYQQFzhIxXeXOCwT6dF1bh7vaOVad2de1vf0T1MJr8/oj683MvkRqKCJdhwaKQz9YN9Zy4PJdNL4JtReO++2cZjPbLJhXFc7Y5z9ZvFfUrYMf6w7cycsgNkXuSKJMZLXA/W3zsukbACBgBI2AEjIARMAIzR8AEi5ljbVcyAkbACBgBI2AEjIARmBoBnMuIA9fKcIJTU6K84XwnfQ0pgUjDNKYzVY5aHOtENZBW6LWyX5cRMTBaI9XTt2V3y3CW43hHoJhqzQwX3fAn6o86DEQu8P5O+vcGwzW45j0yHPPDKY3SiQGfUkGphEUgEKwPp/XGpVfi1OWkQeo/0TiglEhdSq2kSIzCHokWFC6vFqkyXAijGgSlWeov5AI7VBsjKAHkN7xxwIG/LZyjm3RUCAKkwEJgoR4Haa5c3Qqc/tUiOMovuUTXuaHnaHNdMFTwLb3k+GJpCOzqZ3xEVlDcfIWMiAoc6y6NFwXQQ5JPOgq5YLe+jITj2fZgONcbiuaW1Lcn7somw8sUcfECcSG9FJEUvcV8vic92N9fyGYvryJWcNhXZURzcO+xDlNd82p458J3RO9QNP4XZTxTlY35s848izyT1oyAETACRsAIGAEjYASMQM0ImGBRM5TWkREwAkbACBgBI2AEjMA0E8DBjTP6KzLqQxDd4BrFf38oY9e7S0901uLbEiuooUDqJWpFXCMj9VNlY5c5UQL3yb4ve1BGwWFEiolEcIyFBsf5Td54ntEr9Rm4jt8VW1Zx54LSQiHCPC1DkLnCdaqaC77UYI8iLNBehmtBjLhmLhtslsgQq2tOtQRCeSIUiCQpb1wXB/Xp2hhVmsSKQ8n+2P4dP7l4cbIvdr0c/jiuiVCARa+MASAcEC3CmsAYYekFMgQWJ6Qg0CC8EMWC0xsjQoI+ECNK6arUf2suHfJ1H27xNXYMNDYuHFhUyAcSKsCNU52+iQ7hmggkx2QUwqatVsHtNh23UPU28hJrWlV8++KG9iEKeNdJuLnw1MHWSCahMhySHYq5XDo12Hs4PTTAGlRrRKQwRq6Ho76Waz/KJWflaxfFwzPE88MzhThWXlj9t/SZ6CIKyM9XDrMC3y5qBIyAETACRsAIGAEjUOM8swbUCBgBI2AEjIARMAJGwAjMAAGc0zhMcSDjuKbhUGVX+AHvt6obc7yICle3gPRLiB/VGg7q98iIEiDiAmc+kQ84dGsqVmhMOPRfI3u1zDnrcRZTayGm33dItGDOtFEdxHK5+9JDvb5AMOgLxerTKrxdHmWh+gz+aOe+BWsWrz+ZD4byaX+o8Bn193MyIlZoiCSjtX6JB189uW/BXtmNqgnxMh2IKIF4QtQE60BNCRp8mROiCLUOEJmIsmDspITiPDji/EeUQaxxIgk1KChI7hq/t0t08B3ZuaRZYsU6iQ4721f0NCg1FGJHREb6LNYJ82ucjYrM6M9lQplET7xhoKu+WCwGTsYa001KX6UC3IEFOvdUrDH1RGoAp3v4No2mMRgKbw6Gw/5c+ozACb7YJrtTtsu73nx21PPsIAiyVitl5WIFzxzPnrsfy5bK3hoBI2AEjIARMAJGwAgYgakTmHBBwqlf0nowAkbACBgBI2AEjIARMAKTJoDzGEc8TnJS9JQ3oiWul+Hwxvk+QrTwxAp28bPb/x2yamIFjliEjJfLKHCNY5p0R5yHk52d/1Fy/jubzEzKzsfR/3rZx7zr4rgnpdXtMsZCFMQmHY9j3keUhV4QAD4tI8JkRNorpTRSpEWvLz3Yd1TFuO/X79TWcC0y1Bt/iSIkWjQTUkHdJiNlk2sICeVigfseJ/VRRTp0Htm5uL37YGtU70MSBuBBmqdq4hDf3SgjZRROb6IwiLBgTlyT3flEZ1RzfBM5QRQDqbBI1VVqGrfv+J6FLRJMlug9/ZeYqJEm6iP0qzH151VTQ/Uu+vpONB4a6qkrROqzdf5AoVXFxlfGm5PtgWDxSDCUfbiu+eTRYjFzUtEpB7OpRF1qqK9Br6WaIBUNB/2dMqJsiAAh6ma+Nrjy7HAf8CzxTJU3njmX1mu+psSar2tr8zICRsAIGAEjYASMwDlBwFJCnRPLZIM0AkbACBgBI2AEjIAR8AjgsMeZirO7WuoidvKTFoiNOfxbt5Rj33P4EymxXlZNqHi/vv+eDIe0y82Pg51rkNqI3eY45/mda1OYeqqNMeL8/fWyjigq/i3ZDhnRBqQ7Ysz7ZRSWphF9wecPeOMglVWp1kA+m/al+ntIc7Q6HIsfC/gDQUVaDHdfzAc65MRvVfFqBBgc08tlMKJPUl/hhC6va4FoI/HDn1AapSYJFU8r2qF8x33Z0Ku+ZQ6Mn0HADYGF6xCNwTri/Kc/RArX2N1PwXHYUxi8FEWjMfiSfXFffWuiTsW4oyr6fUApn+iHtSCtl44rtuSzwaHUYOxUIFBc3rR4oD2XCkUSvfF4rCGdU3RGbyiSLWSTxSbVs2iLNcR2dz6by+ezWV8+k9Y18rIRwRNE1RD18qyMourzWawAM88Ma8QzxLNU2VgT1pG1m89RJlWmbl8ZASNgBIyAETACRsAIzAQBEyxmgrJdwwgYASNgBIyAETACRqCWBHCU4gCv5jzm37c4yHHAUxw4LbECJ+vNsnfLXloxkA/rM+mffiQrOaRdAW2dx/k4qrmOKzSM87zo6krQl44jMgGj8Zo+W30LoivUECtw1P+a7LqyMX1d7zfKcPSz1R8xgbRIw8WNFWWRVy0LHMa7ZURZIDoMF0fOZzO+bGrQVyi0r5VaUSpq4bVBCRkN/Scbr120pmufClGfUuFtahUwJ65FGieiSXBWu7oUKaIWsqlwUQW2e5Rm6Un9Vsmw7BJnvGWtSA3lIrsRgdbJgECUBeODLYIFYhDXRUyhIPgjsjtkCDKl9FaFvN/Xc6T5QaV0KjYv6T8Yrctc4Q8USS11i6SWYyqy/ZSiL1YnB2JLlP4prOPzSg9VbFowGAhGcwfyuWJPLpUOpAaKsVw615bs63xlerB4QSEnnQZhh4IWzzUiQRCOWBMEFFJPzefmRCUKmRO9Uu1vRZ4FjjOxYj7fCTY3I2AEjIARMAJGwAjMIgETLGYRvl3aCBgBI2AEjIARMAJGYNIEcOJ/VkaKpudV9PJ8fSYqAqc+TvD/JfuzKlf6e333Odl+WcYJFe44fc5JXOjRZ3aUU9DZRW2w677UytJMIVQgKuCQJ0KgqnPbEytw+BJZ8U7Z+8rG9Va9J8KCCAdXgJprE0XwkM4NOCHEEy0YDyLL8HhO91X05ZTaKNV3KhxoXXggGI4gEPDv/pJ4oWLZkURfvLUxnO+R4x9GXIvrIHwwbsYPv6yiGnaf2NPxqIper+070URNCKJTGPt4W2UKWuaOQ5yaEKRyukjGGiFYwA/hBGc4HBFQEC0QSX7fXVDiyas6n21/SmLF44vWnXy4qWPwVrnQsxJWIkoFtUgRIK16jaYGYulMItJb35JYlhyMDnQ+sfiphrau+kK+b3lmqHBhst+/JD2Y8wVDfl8hd4ZY8biu9wXZPhmF1uEy36MruIdXyxDMqkXR3K3veeZ49qwZASNgBIyAETACRsAIGIFpIWCCxbRgtU6NgBEwAkbACBgBI2AEppEA2+BxmuKor+Y8RcSgzsMVMgpKU0ehvFHv4N9kOKOJKBgRMeEO9MQInNQ49V0ERQEho6I/UhLhiGdc/Eah7KSOG+Hg9sQKTiXigygQCl679h29oeYEkQQICDiMGRvOeopSV4va4FoUA2cuRJBwXKmR1ig10NPqDwbz9a2Lev2BwAICCCRQDMabUjmlTYoOdtcdbF40wLxc6h/GxfXh+i0JAKvk9D+475GVjYpaWFnM+39N301ErCgNRfZcTqrn5ksEDDU0ECYolE6aKJzlRHvAjbmRsoroDCdiDIsfGv/FA10N/3vpJccp+k00SlLBEYd7jzffcXz3whszQ5F1iq4oql7FQDYZSvkC+XA+U7hM9SpaFV2xbqAz4Bs8JZUjJbFCURteI/UTYs1dMtIicX8QWcE9VjWiQMLRczM699/Bl2gV1oxnqLKVP3NWv+LcX2+bgREwAkbACBgBI2AE5iQBEyzm5LLYoIyAETACRsAIGAEjYATKCZCCqczhz084vEnZUxFdUDrrzTIECyITyhvFrD8l28rvZamfSsdU9M+/k92/lUmPM1QpQJR1jMDAMTi8cbBzXVJRcU6loxunMEWoEQcYP0W198s+LiP91FqZq5VA2qQ9MiIRRktHRFQC0Qp3yl5XPtlCLuPLDPYuCEViB6INLXF/wJdo7Bi8T4LF5ZG40kalQ3BYVX6O3uO9Z4w7FE1x/9M/W9OQ6o+9TbUvbhmZLanirNE/VhMrOBrBhggKGoxwlPPKuhLtQbtQhphCWibSdl3uLoP4Eooo11PRv0iWUWorSnVcGArn9rQs7l+gqJC+gVN1iUAg15ZJNUmvyUSTA7llJ/cGl4XCAV9SNPMZxArSTA0PnjUhqgKe1AvZJeP+ykmYmO8OepcOiuiKN8gqi20DCRbcs6yRNSNgBIyAETACRsAIGAEjMC0ETLCYFqzWqREwAkbACBgBI2AEjMA0EsB5jKOe3fBscce5/KcV16sUK0i/9DPZAYkIpSISrpXXo/C+I+oApz27/7kOjvQ6CRCDVdJGFfU9DlzSKXEcwgWpl0hxRGRGZSOCAMf7KhlCxAdlt8vY1Y/rHIEC0QMRhF3+GP1XRnX4cKKrlgXfUwMCMYZ+SbFUakUpDNlU0jfUdWxl0Ve8IxqPqXh2oVuChT/enFzeECrglMYBjXhAY/xEFRyTCNCoSIUTvcean6/aFUSq1Lo5sYJ+KYYOZ2paMB+iPBAtnIDBWo5ILYV4kklGfIr86FLh7QdVgPtFqmWxsG15769IjDnc+Wz9kVza155NpWPpobAiTrINuUz/gswgOP2+HGJFQVEZBV9c5hrprv5HhkDCPUaqqsI8i6IYbR0RLLjvuG+riRV/p+/vlPHMsVbzXcCp9f1u/RkBI2AEjIARMAJGwAiMk4AJFuMEZYcZASNgBIyAETACRsAIzC6BikLXOEwxBID2MUaGw51C0qRVOsPxX+VcBAv6RnDAeY7Awb+b+b7a+RyH+IDDFyc39S4QEaqlEaIfHPNEUdwjQyA4KXP7/PGob5chJJASyokeVR3EnmhBZMdPvX5JM/W7bk5FeeOzmaRv4PiBaKY+emrZhnzvglV9jUoNtUQRCaSQOiQjGgUBgbG1SgzYkRqIxnuONucK+QA1PHBQI5qQsorUU/tliAiIKrVqbh1ZJ2puONEI8YdIC66PIQhJgPD78tnAqVw6FEonIgslwJQKowtSJBjOxWINfYlsstiQz+QWZpKD7USbUNejkMtrYalXURq2i+Tg/b0yWDuhhHmfT4Wl4c3cuW+rNZ6xUsF5z2q17taPETACRsAIGAEjYASMgBEYQcAEC7shjIARMAJGwAgYASNgBM5VAuwKRygguuDnZa4Wg5sPv/2zbL+ECpz/422u7gIObP69TI0EHOU9RFm4TpyA4hXnRnTgGASOUmREZTSGdx59Ek2BMxwHMGJDuRjBe2piEDXC/KiZcdZxewW4cbAjKCCaDAsWpROlQBTy+RvSieRFnftyn116aXFfi6pD+IO+i71rc96VMupmJJJ98R/vvX91uv9E4xoJAwgTLnLkFm8gCAjT0WDNmMobTF26LYSjUg0NpYBS9Ei4vVDwx0UvqZoWPwgECoqcKG4KBLPPxBoze/OZ5C2FQqAdoSKfy/oK2VG1qj9WlxT3Zt1Iy4WgNOcKbFdJWQYKmGXPkq5svOvEfUt6si1VTkBE+ncZgtFoKb7Gex07zggYASNgBIyAETACRsAInJWACRZ2gxgBI2AEjIARMAJGwAiccwQQA+TAJU0QhZrZ9V/t37V36PvveY7WiczRpSVidz+OXHaXIyKM6vGmVoXG41I4+aqJFZ7wgCDhagCM1p8TMMaddscTLRgjzuXPy/5X5YSL+WL7yb2Bt++8PfzeK38hUxdrLC5XlEVYLmjEHBz1h5UKqvPUwbbtQz11axVdQbQGxZeHi3lXgYiIwHUrxaKJ8B7rWMQDojxYYyIAMhpnR2owOtB3vGF308K+kFJdLfIFiyEVsqjPpn0te+8r/JrSQS3M53KqVZEupcdSY31YT9eccEQarge83xFnRnBX2i3fZ770icoxIjYxHl4zWluEp5lqXBcVi6gIxDS/7j0iZViH4TaW0FUxWBhzD1QTaniGKP5ORA337rjvy5kCYtcxAkbACBgBI2AEjIARmD8ETLCYP2tpMzECRsAIGAEjYASMwHlBQM5ZdnlTpJlIgr/0Jl3NYYxD95QsonNSo0Q8VGPmRIXTBQ9OF7ym4PBZiw1PoP+arxNOdTVXA+Nrek8kwivKL4TPPpvyNx58PPQGZYpquOh5uf54czEZDBdPBUO+nSrKvUgRCYrUyDWSEkqiABEXl1UZLNdxxbGdqDPZOdEP61RebNtFuNAnAgJihXOmN0mc6NGqRPLp7IlnH/L3Dp2KP7P2+szxbMpXGOz2t2p+1/ceS7fmMupyZKVwJ1aQAovaITj5qcmAYMFajyeqgvsB4+8oGJO+6ojurwPMoUqR9clyOdt5RJxw/1NjhciaDTIia6i9AasJNe95KkUQyaqF8/A96aJKBcjLO5+gKDKhcdnBRsAIGAEjYASMgBEwAucnARMszs91t1kbASNgBIyAETACRuCcJCDnKv9+pSbF82V/WTaJWJUJvU7fkeqHSIudsmpFsEfjgKMcoYLoA1IE0c6FmgY43qnHAKdnZO8qnyD++0LO97zDT4R8XfuDvsaOwjckVOwY7PJnFq4pFFVgO5QeyhTy2exJfzBEPY7R6lTg4MbBj9hQHrUw0fuKfhAoiJahP17LBQs+xwr5HGvh9weCC/LZVFcuk1akhT+TGkhdtOe+QtOBrbG6YqG4gQLaKqatqAp6OSMQYLe+/bDH5mm9PiTjyJQiVMZY2+EIC1frgeLUN8pukx2UcX9R1P3oRAFM4njWdo2MQu8IJQgnCEfUPSE12UQbYgTCC88Uz0xlW6UvVshcMfKJ9m/HGwEjYASMgBEwAkbACBiBcRMwwWLcqOxAI2AEjIARMAJGwAgYgdkkILGC9DsbZX8k21Qxlm36fHmV8eGAZSf9SZ1/5Gy5/qvsFj9XCwyTpulu2X7ZMtlryrngx1cNat9Qt3JBdQd/Ub9dre96BroCJyQVtAQj/uXNS4rxcND3kio8EQ4QEXDYj+hWH3D6O8EB5zkiEoIEBb3P1ohYKBc92MWPeIEpTVWxLpdJxQuqHh6O1++UWLEgMzTgz6aGIoVC/kIV0r4wxYzLyiucqVWUBAXEBMbFK1EWRCOMQ6wYHjrjJJLh5TLqPVDLg/sQFtx/cQS1cRZ2HwPJWX926ckQ0oh+oMH+rBFA1XrUeBFgEDzWyqqJFa5vniHWxdJBTWXl7FwjYASMgBEwAkbACBiBMQmYYDEmIjvACBgBI2AEjIARMAJGYLYJyLGK41ulon2/UOFYJRXU22TUUCCa4jcqxopT+jEZr0H1QxHrOed09Qoq4+ynjRBKJpF2B+c1tR52ySgojXAwIj1U6SLPUbhAHy8gOoFWyBceUm0Lpf9RzELR168DE/5AAOGDWhC98toPKNbhEn3o1SsRHdT4cGm0cOondNzjqifRomOW6Iek3rOLH1FCYykq0sHPNV0diIol0/fFYlZ9Z5X+aU8+l+lND/TeIIFipa+3a3c+m16vEBCNjgFzuTGX89s6iJRSRFU8LsPRz32TV2TFmCeXDY6LMWac+0T5UC+E2g70/bCMaBz+vhq11knlRCf5mXsZAWa9NxcEE6JhJlRHw0sFhWBR/oxUDunfPGaIJOdChNEkkdppRsAIGAEjYASMgBEwAnOFgAkWc2UlbBxGwAgYASNgBIyAETACVQnIsYqz+yoZTndS8Lj2Ub35kAwH9BYZwkSlYMEueKIC2IkemItihTcZ53l3ogVfT8SZXsnO1X5gZzz1GqjVgGP7tWPdZoVc9p29R5/11bUsyIVj9cVgJNYmV7WCGbIpCRFtEgpOhiKxRLGQD+Vz2YFgOJIOBIIxHZBRzqYTGnawkMstz6YTJzi2kMscjja0KptTkALfEkTyhyRg9EgEWeH3Bxv1SjqjEY2LSbQopAa6b0j2dzerP52HSFHUepZjOQPRU+roYhl1KUiNRfuObJ+MdEnUNMlOUKhwY+NicCWagvoeOPoRQxAoLpUdliFizERjLi4SheshUE1IKCkrXM+zwf3Hs1LZ/tOb53jqe8zEvO0aRsAIGAEjYASMgBEwAvOcgAkW83yBbXpGwAgYASNgBIyAETjXCHjRBm7Y7GgnNdG3KuZBKqMfyNjhzzGIEtdWmSuRFx+TfUT2mPpOz2HRArHCCRfjCh1w85UDvtoyl6IeVJCb3f84synUfL/sH8e6J/KZlC/V3yNBItcWjirTkEIuMonBOn/A78tnM1viTe0+CQ0UlcjkM2lfIRgMKmVTPBCO5FQIoyfR27U6k+hfK8HiuA5aJtHhSCAU/rYEhyOFXPpKiSCL4k1t/lAkng7F6uokYJSEGmkUpdAPRVTUSfDwpQZ6JFLIV67vJJawxmeIG2VzIcKAud4pI+qDOSMoPCDjt8lEVVSiIu0SAtlWGQIFha9dEXK+n5BoMNY6lP9eEWmDcIII5dM9TTFsPk8oAqKs2DZiH7VOeFYqG1EcD3pznMhw7VgjYASMgBEwAkbACBgBIzApAiZYTAqbnWQEjIARMAJGwAgYASMwHQTKxAoc9i2ym2R/UnYtnMJvlv1UDtxSChydg5OYAtPUF0DEeFnF2J6nz0Rf8G/fu2TsjJ9rrbJexlSiK0bMTWJGUqIF6bKoJcHO/D/3uL50NAgSB3yZ1JAP0QAtQVEUKtatLE0SKQpKxSRxwidxAiEBh70vEAwRghGTuHCZ6k2cKmSzEgwkMlC0W33p3HW+dPI97noqol3qT5EZvlhzu0/ChQ7LSxQhExVHFX3Z5KCvmM+f7uV0/qrRxArWnygK7gGEj+/JELJc6iTeTzT9UzU0DIK0T4giT3g8KUpO/9yXFHWfkGhQi5twCjUzeB6ukV0n4xmpbDxLFNqG6xlCzCRSldViutaHETACRsAIGAEjYASMwDwnYILFPF9gm54RMAJGwAgYASNgBM4VAmViBXn1F8veLvvfZeM/oPevl7G7PVN2PE5inMU4Vu+QURB5ucz9Wxcn8woZrzjuyfc/F5srysDYaiZY0JlECyIt2JFPLQIc7DiivyG7UsbOenbZw+i5djqqwVf0y9LJ0wPKnR5WRmKDL+X3ylyfDgY5rTOU/pfohrM26k+UIjMkgCR7OyWIREvRFaW6FAgciqpQJMfpiIvR2336iSLapAWjjgTj5wRqVfDKfcRcC5NMAVXtyq5Wh4toILqB+irTFlkxFssp/I7ARxF792y4dWMuRI/wLPFMJSROzLgQM4V52alGwAgYASNgBIyAETAC5zAB/rqwZgSMgBEwAkbACBgBIzALBJQGx9/S1r6gsam5pb6hsamuvqEhGCq1cEAtMTg48PTO7Y8P6XUWhjfjl/QECJzMq2TUqvi4NwgKDLOD/vMyahOMyKfPTm+dy3krZb/rnU8f1DKg4LRrv6M3P5Qd1DlzMcpi2plLtODf/0QhkEaLItg420mlRfQCr6+UUVSatl3WIaPY+fQ1pZsqSR/eXyaIJC7KouKiP9Nn1pnUVtQvoag4EQ77ZcdlpIzCsc79wWspamWUdFkjuvbuPZjQv6sNcTbRyP0dBT+MljpX7ivNl7kiVBBlQ8o014haog4ITDE4H9C8rIbFiDvGPhgBI2AEjIARMAJGwAhMFwGLsJgustavETACRsAIGAEjYATKCKy/dOPln/iPb/zw+9/86hdXrF67fs36iy9duGTp8kgkitN41Palf//kRz74/vf+3nTBXLV2/cWf+MI3f/iW19x28/GjhynQPCvNcxjjSF8o+2VZefHsD+jzT2U4pYedyFVy+pOWxxVE3qD3OGXLG6wp4N2g6/XN513jZdEnMOXf/BiO+JznfM5LvKAeA872hzxW39crDmqEHjjDi4gW2gtlCyp41uYjURyltE+l7igejUBHOrBPeeNglz8CAYIERxEZgPBEAW0a4lNpbt5x445O8eo40Af3BVEm9M31jsqIRimOkvrIXYMIDuycaZoz9wQCFXOu/O8PAh/Pzm4ZzxLPlEVXnDOrawMBayZvAAAgAElEQVQ1AkbACBgBI2AEjMC5T8AEi3N/DW0GRsAIGAEjYASMwBwnQATFX3zwo59u71i0+A1v+a137dn15PZtjz50/7EjBw90d3WeHBzo7yOaIpNJp1XkOJcnH46adpoXd23f+uh0Tu+6m2590ZLlF6xU3WMctbPZcKKukpGiiLz6y7zB/H96pe4EtRdGEytKuGTsDqdAcJ3sdVUmc4u+gy3RGv2zOdkZurZzTJPy6UIZzudjclgfp+6BIg9wRKc84QJBgM+kzYI1zmwiK+DP94gZiAik3nqx99vdeqWGBVxJzfQC75XvKZROnzjzSc9FwwFOCqJSgW21L8s6Zaw357uUWHzHWNnpz3tXG4J1JS0Y40O8QKCojKAYt1jhjYEX7v1NsptlRFiQGgkRh2uVrlF27Hx46+rDIEKxdpUNoY9njmeJqJH5Nv/5sIY2ByNgBIyAETACRsAIzFsCJljM26W1iRkBI2AEjIARMAJzhcDSC1auWrP+kg3HDh868NoXX7txLqV4uuKa62/KZjOZw/ufZVf5bDYc5KSoYXc3qZ1ul31N9gM5THFQj6ex0x5HNk5ndsfTZ3lbpw/UbcAJzTHzPc0NwsAamau7sF7vccbD6YQDg3Ah0cJ9hAmiBeIPkQ6IBi59FEW7ibIg0oXfcOiTMopaEji3V3tcERbulBG9cUzG3xw4yWGOeEIEB99TvJrr8MraMyZqJxBlQb0NjN8ZvxMzeK2liMC4GBP3HBEnpJsiTRJjJ8riXKxNoWGftbm0V9Ry4ZmobDw7HMOzdF6mThsLoP1uBIyAETACRsAIGAEjMH0ETLCYPrbWsxEwAkbACBgBI2AESgR273xiWy6XzT58/913zCWxgrFdvuXa6595eteTjG+2lks7/vk3KQ7jV8hwXH9bhrDArnt22o+34cwmcgIHN0Wlr644kWLcF8kOyti5fz402F4gQ1zAIY8YESAtUHlKrIo6D/BzKZZgRMFuzsPBDTtXvwFBBI6IGkRBkFKMFEM4uxE5WA8XCcGxGCISognfI0ZwLFFEHO8c5K7/kqA0nhoUU1hI5kpqKUQSonIYB3Ni7IgX1EdJzrMoA9aBOiU8CzwTlY1nBy48S5YOago3l51qBIyAETACRsAIGAEjMHECJlhMnJmdYQSMgBEwAkbACBiBCRFYvfaiS1RTu3nrQ/ffM6ETp/lgUlQtXrZ8xX133f6jab5U1e7L6laQJujdMkQLdtv/t2y/zNUsGO/wcLKSgoh0PjjCKwUL+vl5GQ5Zfp/vDR6IDAgEOOTdv/0nPHdPNKjmvEYEcQ2BARHijFYWwcHvPTJECZdqiFcnUsxG+iHYEE3B/LaWsaLOA9EG2LS2spojZ3AYpYbGVMbD+pPui2ehWvuivuQZ4lmajfWYytzsXCNgBIyAETACRsAIGIFznIAJFuf4AtrwjYARMAJGwAgYgblPYNOV11zPKLc98iCpc+ZM23D55qsYzJPbHkMkmNFWJlaQsugmGWmEHpc9ISNd0GRrTOBA3yUjnRCph35LRvSIS0tEqh8ctgs1hoNeAeoZnfsMXgwHPBEqpG0i8oHUR7Ag7dKEWkURbyc2lASM8TjUy6IkykWK8jHMimOcyAmvCPU+DeZ+GXU6qKlBijSEPMSMcnFlQtwmcDDXIPLBpSpz4lBNuWiupXvfuw7PAs1F1BBd8knZd2VEmZSLUROYih1qBIyAETACRsAIGAEjYAQmT8AVvJt8D3amETACRsAIGAEjYASMwFkJbNpy9XX9fb09+5/ZTeqcOdMu3XRasNjx+KPspp6NhhP9WhmOU9Ly/I+MYr8IFpNtOF/Z6U+0Bs5nGo5Yt3MdB36jjNRT9Z6zerLXOhfOQ6BwqZeIIoAzIsNkUv24It5EbMDQObzPBQ5nGyP3DCmvKCy+W0Yk1E9kiF78VlPRoHIguge5N2MyRDtENiKDEBXg6+7bKTP27nUKjHPvs34u3RrX4Bmh8czw7PAMTeu8pzwh68AIGAEjYASMgBEwAkZgXhKwCIt5uaw2KSNgBIyAETACRmAuEbhs81XXIgoU1ebSuC6+7IotqWQysffpnaRImrFWFl2xVBe90bsw6Z+IqqBuxbAzfTy79ysGDmNS+DwrY17snL9QhuMepyzOYBzvfydzu9on47yfMV5TuJBzxO/3mPJvf+ZOwezJNM4nTRK8sPKIgMn0NyfO8aIscNA/LaMOB/eJ+zupOAP1K+BIMXNqZhAN4wQFxBNEplrVl+E63PMITm+RXektgHs2eFZ4Znh2eIbm1H+v5sTNYoMwAkbACBgBI2AEjIARmHYCFmEx7YjtAkbACBgBI2AEjMD5TKC+oaFxzfpLNjz5+COzFcUwKv6LL9u0eecTWx8t5POl4sYz0cpSCy3W9dhNTmN3+4MyUlNR7LnUJiFWuFNxtBKlQeHu78hwvrod5ByDo5Y0Xexin/UoC2+HfU3xw84z1pa0RqT3QRSifsSEU/14a0FfCBVujYiQCZNmSOZeaxYRUFMg4+uM+SHmwIhIFBz5M+G0dzU8mrzrE4nFM0G0Q2Mt7o+y6Aruee59J1ZAhmeDZ4RnhWeGZ2cm5j2+VbGjjIARMAJGwAgYASNgBM4rAhZhcV4tt03WCBgBI2AEjIARmGkCl27aclVAbRbTLlWdcktb+4JFS5Yt//F3v/GVmWJSJlbwb1DSzrCb/esyHMRPyoYLNk9BrHDTwalOweltsoQsXjFPrrlahtMdB/G0R1mUzZ+h4Nh3EQ8+/YazfFisKR/rVFlQp0P9lwpHTzFaAEasESwZK2NmDji8+Q0H+4CuNTDF61Qs1fR/rGDs0opN/4WfuwIiElEWiCSkgkI4gSvPSC0aG9UukBHVxL1f2XhGeFZ4Zqreh7UYhPVhBIyAETACRsAIGAEjYATGImCCxViE7HcjYASMgBEwAkbACEyBAOmgOH2uCRaXX3ntDYzryW1bH5nC9CZzqnPUkz8fxzeO2X1yGA+LFZPptMo5ONDZpc513iGrFGZ+Ud/hcC/VdPB2sQ/vKp+qSFBtDq5PXcs5+Xl1Tn/mj1N5Wmom1EJA8FInEaXhUkLxSu0FV8uiTe9xuh/WHPt1fK1SGdXolpiz3bDmCAaIFjDknkT8ITIG3lNqZREaiHObZdz7lY1nhHuQZ2baxbspTchONgJGwAgYASNgBIyAEZjXBEywmNfLa5MzAkbACBgBI2AEZpvARgkWxw4fOtDd1XlytsdSfv0rrr6uVDti5/bHZkSwKIsuIEf/FTIcs7y/W4ZjdkoNMaAigsHtkqcuxh7ZCdmisouQEoed5o/LqMvAccOCBX1Nh2jhOY/ZOU/xYwQKGGyRHfTGktYrNidT8ohJTnPAiY7whGMbsSLoceVvCxztON+zOq5AdMeUFrbs5Ir1db+UUlDVQpCp1Tgn2k+ZEERKNOpXILLxfCBg1IIfjLjHEZNeJCtPB8VweTaekPF8WLHtiS6gHW8EjIARMAJGwAgYASNQUwImWNQUp3VmBIyAETACRsAIGIGRBBAsHnvwvp/NNS6br77+pqHBgf7DB559ZgbHxr89qVuxXoazHif9Tjlsp2tHNw5fRImbZF0yHLKkRnLpoXDeImYcl1HguJQ2aQaaS8+D45gi4Js8Fl/V610yeMxU/YQJT5f1KhMPYIZo4dYQ3qQUmq41LR8vHEtptRBHvOueEaEyHcLThKGNfQLj5x4l4oj7k9RMpbnUQIwhsoIUbK+Wcc+75p4FrsszQp2dCdc3GXtqdoQRMAJGwAgYASNgBIyAERg/ARMsxs/KjjQCRsAIGAEjYASMwIQILF66/IIFCxcv2f7YQ/dP6MRpPjgSiUYv2XTFlTuVDqqoNs2Xc92zy5uoAlLOwAMnaadsOtMG4TjfJ2uWPSDbIKusZXGVvrtdRqFhUuKMiLJg8NPg8OYaOJGpKYCAQ0QFUQuMb7+MugXwmam1mcot4Ip5I1oQKUOkCmvtCjlPpe+znUv/jTIXqeKiERBMRr2nytIjMcZaiAG1nB/rzT3IXFwEy7jvgbNEoMBpjYx7vby5Z4Fn42kZz4rVr6jlilpfRsAIGAEjYASMgBEwAhMmYILFhJHZCUbACBgBI2AEjIARGB+BDVdceQ1HplOp5Jr1l2zIZNLpQj6fdyKBn6aC3KFwOJwcGho8cezI4bP1HK+rq6evgtr4RlD9qMs0LkSLvU/v3DFWP6UhBoPBfC43VUcmtQ5Ic4PzFKc2AsF07+bG2csu8p2yL8peK2uSIZSQiolGeqrrZHtl7G4fIVqMxWeiv3vpf5g3aX8QJh6T4TgmZRi76hfLcPwjWMzZVibiFL2C3oguzIv0UC7aYUr36RiT5zpE6hClwhrC839kpFWC4xnX9sQKzuMeWChL6ju4p2oQxTCltaoQxWrFDdGD5457inscTq65Z4BnkWeDZ4RnZdwCyZQmbCcbASNgBIyAETACRsAIGIFRCJhgYbeGETACRsAIGAEjYASmiQDCAF3/2Qc+/MmxLnH8yOGDL7vuUtK2jNq++pMHtv/kv7/5tY984P3v46BbX/KKV//yr7/tnc0trW3/84PvfvMzH/3Q/6k8+cJ1F1/6xre+490XbdhUclZ+4V8/+v+Wrli5mvd7n9pJ3vqqjT5/70//+h9ue9UvvT4UDoU//eEP/k21/seaF797RabX6i0pfHAWk4JpOiMryoflCkSTm590Sz8nc2IFx7FT/4Uy0jExNoSZaR2bVwfigK6DWMGau8gTBCQEk2m9/njWbCLHeM5++FK7YiYa9xG1Mni+SHFEdMpyGaLFUx7DEc73stohRLYgEK2S4ZwnTdhOT3QZUS9iGiJrZoJN+TX4W497mugX7nHuddfcM8AzwbzdczLTY7TrGQEjYASMgBEwAkbACBiBEQRMsLAbwggYASNgBIyAETAC00QAwWLXE9se+8gH/uJ94QgtGg3xJhqJhr0vuHR/X2/Pow/ci+Nw1IaAsHzFqgvdAe96319+4M3v/IP3UcxbQRqBX3/Hu9/7uX/58Adzueyws/s1b3zz2/74bz700RNHjxza+tD992y+5vqb/u5j//afB/ftpV6Db+cTWx+tdsGFi5cu+8zXvn8n6ay++19f/Pwll12x5bff82d//b1vfvk/KCA+SVw4h9mF/6TsWVnNd3KP4mCm3gKRE0QskKP/ZhnO7vJG0WtXDwHn7pQFA12T/nAQs8sdESRfvotf79M6hvoZ35ERKUB6KJhQ18PVL5gk6nl/GpxILYZAgvhGOiMc84hRpBsjaoBoj8qoIApPs7Y46BEtXic7IvsXGfcHwkctilzXfAHK0j25VFbjuQb3cqnGh4x7vLJxn/FMuNoZZ0R2zAPRZjyc7BgjYASMgBEwAkbACBiBOUTABIs5tBg2FCNgBIyAETACRmD+EEBEuGTj5iu//NlPfvSBn93xk6nObMu1Nz6PPh6+967/+bXf/J0/QKz43te//IX/86fv/u10Op1qaGhsqhQr/vzv//lfv/WVL/z7377v995OSqfGpuaWb9716FOr1q6/mPRUT+/YvrVyXCHlp/p/n/7iN9oWLFz0ltfcdvNTO7ZtXXfxho1f/cn92xEuJiNYeBEF7Hyn4RAeFitmyCHKNUlB9aDsC7LfrbIeG72x4dx1zu5JiSrebn6c49SnICUPESX79T0O9PK6CTjIEXBIBUaUBePEecz1J3Xtqd5n59D5iBWIZ6R4clExMMPpDkt+LxcscPSzJhyDYNUuWybje6Jc+LuIdSId11xtjLUkWIwxQI5hPqRgI/UV93a1xrPAM8GzMSeFmrm6EDYuI2AEjIARMAJGwAgYgekjwB9k1oyAETACRsAIGAEjYARqTGDlhesuqpeKsPXh+++pRdfX3nzrizIqYDE4ONBPqqb/+sK/ffLP3/22NyUTiSHqYhCl4a5DGqj3/vUHP8K1/+aP3/U2V39iQAfdodRRHLdr++OPIlpUju1Nv/Wu9xAZ8ld/9M7fQKzg91g8XsdrXh1Ndi6IFp7hsC8Vsp4hsYIhu2LG7KbfJiMVU2VDEGIX+hKmPNl5euexex+nOWmJ+Pc2aYfok3REw82LuOCYEzKiToiuYE1qVcNgitOY86dTA4SC0Qg8RNHcJ6PAOuwrnfp8RiDCme9Sf8EZp/6tMuo8sEb8PpdbaV5EXJQX2a5ScJu5cC9zT5fEzorGM8CzwDMxrXVb5jJMG5sRMAJGwAgYASNgBIzA3CNgERZzb01sREbACBgBI2AEjMA8ILDhii1XU1x72yMP4kSdcrvyuptueVx9vfevPvjPT2x95MG//4s/qhYlULrO+/72/36MlFMfev97fw8xo/ziA1It+PzYg/feXTko0k695Z1/+Cf33vGTH1Arw/1+0WWXb+b9nl1PjlrzYsoTnMYOvELXCAHsoCcFDvU02HVentN/kz5TE+FDMoQDduhPdtc5qXjYwb9UhmCBY53PONUzci4P9+uJFmPtmJ9GOjPTdRWHOheeSHqj8oG6SAoiU/5Ttk6GCPGIjDoWFNIekdbLuwecYAF/RCKO557gPeeQZmpONk/cG+99wj2HaHOZ7A9kCBLlDTY/lvEsMP/0bBcdn5PQbVBGwAgYASNgBIyAETACs0LABItZwW4XNQJGwAgYASNgBOY7gQ2XX3n1vj1P7VRAxJRTzNTV1zesWX/JBmV9am7vWLjodS++fpOLmqjkuOWaG26++obnPf+H3/6vL1E/o/J36lPw3SMP3HNGzYzX/Opb3k5UyCf+79/+hTsvqvCKN73td/8QgePo4YP7z9V1k0PW1bJ4RnP4tuzVskvK5lMqSq52nYxjcF7j4B6vk7gcDefhAF8gwynPdXCqIxKxJiMKQp+rTCc5bsQcUjPhUOfZGJSYUZ4ma7zdujoW1KyAKf0hCLlUUNXWDUc9dRv2ylbI7vQ+8zfRqelYFy89GGmrRi1qXeNII+43IqIuknEvk5assjF/ngHu8yzPxnih23FGwAgYASNgBIyAETACRmC6CZhgMd2ErX8jYASMgBEwAkbgvCSw4fItV29/9CGcqVNua1VDwq+2eOnyC77y+U99fP8zeygyXLX9ylvf8W5++PLn/vVj1Q64+LJNmxE7tj3ywL2Vv7/qtW/89Scee/iBndu3svO8lArqQ5/8wtfaOxYt/sPffOMvTnkis9+BS2lF7YPPyt4rQ1Qob5fqAymdKHC+UzaZAtzs4Oc8CkLjrGbXPyIFfROlwvvzseFIXyOjhgRsYLFPlpJjH17DjvNxOvERJRAo4In4wedRBSYvyoJrUJSbyIJOb504h/Nr6rj3Cq+TBoy0U0T4ME7uwemsUcLfd9y73MPcb5WNGinc+zwDMJ90mrcqfdtXRsAIGAEjYASMgBEwAkZgygRMsJgyQuvACBgBI2AEjIARMAIjCZCO6aING6/4xhc/+6lasKHoNf0gNHzuEx/+h9H6jERjsRtvffFLDx949plqqahI+UR9CwSJIRXDKO9nyfILVq68cO36v//z9/wO319z4y0v+LMPfPiTi5YsXf7ut7z+1XueOjfTQZXP0XNYOzGBmhGflr1VRkHwm71jb9QrKaPYiU9qHT/pjCaSMse7Do50HPLseMdBjmO+VVZTp3i1e6Ei/ZIr1IxwUip4PpG51OL+LesDwYLUWBSCpsbC5R4bWCEenJXNKCLGWUWKyvF7cyctF4Wmh+tVTFOUAcxJVUU0B+wRB7guokGpAHsN+bq5cM8iVnAPcy+79jO9IdriMzLufcSK/CzeCzWcunVlBIyAETACRsAIGAEjMJ8ImGAxn1bT5mIEjIARMAJGwAjMCQLrL73s8kgkGt1WqwiLiy4lF73vzh9/79vHjx6mHkLVtuWa628mKqK8/kT5gdfcdOsLidTY+tCZhcC3XHtjqTBvMjE09G9f/+HdpJbas2vH9je+4tarn9m968k5AbY2g3C78kn5hNP2n2TUryhvH9WHV8lwMlPnoigH9xkO5jGiANhFDzeKQPNvbj7jrJ7JdFA4rxEJEAcaZaRi6tRcuiiAXhucE+oFRzrRFVybcfGe6APesx6IaLV04o86uBmqHeL4I9Kw/tSSYA1IGYbVpHlpp7jHEC24Zztk3MPljeLaP5BxL8AakWhGWNdkktaJETACRsAIGAEjYASMwHlDgH9EWzMCRsAIGAEjYASMgBGoIYGNW66+rr+vt2f/M7vZuT/ltvbiS0sRFt/52hc/d7bO1l+6kR3rvkerFNTm+xe/4udfy+vjVdJBXXHVdaXd2H/1j//yWepcvP8PfvvNr3/ZzVvmmVjhIiVwHJMS53EZkQ84zisbKbAQK3A2Ux9heDf+eBbUc4hzHWpZkH6IQt68n2wh7/FctvwYxsu4qVmCIECNDkSpF8kaPCf3RPuc6vEIEhg8dsmIPEHQceLJfHSgMyfuNdafVG5OlKnlXN1ac69yz1ZL38Y9zr3OPc94UhZdMdXb2c43AkbACBgBI2AEjIARmA4CFmExHVStTyNgBIyAETACRuC8JnDF1dfdSC2IolotQCBEqHZ37313/vRHZ+tv9dr1F3PNaumg2hcsXHTLS15O1IBv5/bHSjUqytuiJcuW93af6vrb9/3e2+/40X9/q6BWi7HP0T5YF8QDIixw5lOr4qUyHOfu38fL9f4mGWl9cK6zI34EE5d6abRIi7Jd/LPFknRE1DNYKqMAM7v8KXq9R7Zd409PUyqkM5YdRroeznpECsQT3j8gIz0UfNjxP98a9xfRDNSvoJYF4gziAp/ZOFar+4K+6Jvi7ghi3LuuuXuaexwBFc49spr8t2m+LZjNxwgYASNgBIyAETACRmD2CZhgMftrYCMwAkbACBgBI2AE5hkB0il95fOf/ngtprV0+YpVTSo+8f1vfvWLuVz2rAWgW9raF/T1dJ8alLpRee3Xv+Xtv0uaKn47dvgQO6xHNJW3aD98cP++n/7gO9+oxbjPgT5wJLvoiR/rPU50ihQv9sZODYAPyKhD8a8yalpwzmykUposTpzSpIJixz1rjqOaKJy3yKjfsUNGFMi0N4kVCD841WmHZS6FEamKSJNVK+f9tM9lvBdADNK8YU4aKO41xATuIwSLCc+3ojaJGwYciaRZIvtlGdFYXMs16mUgVnCPcxzrzX1szQgYASNgBIyAETACRsAIzEkCJljMyWWxQRkBI2AEjIARMALnKoFVa9Zd1KFK1VsfvI8it1NuF192+WY6ufeOH5N//qytrr6hsavzBOl2RjQKav/qW3/n9/ly57Yzoyv4vkmKxamukyfGusZ8+N0rio3jdr8McYdUSez8pz6IEyxW6T12gYyIFAQMXp+RnVU4miOMECsQAth9j4MaxzVzuEr2NRkRIzO5y95FAVB4nIgPClHDm/s1OVORHjO9NtQKkdDAPYZIAW+iXCbMfRSxgvRPa7w1RQx6uYyIlfIGY5d6a5veI6D8/+3de7Bud1nYcSVAwsXWGVGoCJwAISQQ7sRauSOCRC6WiziCZbCOtDOtbYf+UW3ptNM6o2MZrbWOxdLx0gFrKRchgwIFQsCGBAJGJNzCwQBCKWoLhCTc+nwPa8XNzjmcfW77dj6LeXj35X3Xu9Znrcyc/Xve53lu1A5qu+8E70eAAAECBAgQILBVAQmLrUp5HgECBAgQIEBgCwJ/8xGP+f4brv/CF6668orLtvD0oz7l3Ptc0Cf/v+nyt7/1TUd78o033HD9Wbe5bS2Ovm77Z//mRTdVe1zzoQ/U3uhm23Wf/9xnz5qJ3Ud7j/3y+2XB9oYGUM85/eFElRO1TXroRAvKH5o4Z6IkRQv/LfqXzGjx99MTeyFpUfuf2gC9ZaLh1lVb1Iqpe6kEwhnNstjGxevuzQbI51vCpE/8d0xnznHcNIz8KMPM99wtuPh2fidzK1nRcO3uye7NWn11r5a0qOVXyanaT715otZbl0/s1LD1k3ne9kWAAAECBAgQILDPBQzd3ucX2OkRIECAAAEC2yvwqMc98clXXv6/Lv3iF2/sk9QnvJ1z3n3v95mpmvj0p/7sE0fbWQOyp4PU3e9xr/Pusz737zz/p/7pwx/7+Isuu/TNb+xnn/z4tQ3/vdn20clk3PXse5xT26j1l7eY7aK//cPP/pe/8Cv/+WjvvVd/3yfg59hLQJTIKXHx0omGE5esaKvC5UcmWvDveS0Q9/Ve+Hd092CfsG8Bu+qZrv1rJlrsbvviNiYr8qq6ok/412brzyeqBrj3xDrbYTms7XkoWbNDw8dP9ASz7B7sXuye7Ovu0UPVWLN173YPdy93T3dvf3q510/0vb2eAAECBAgQIECAwCkVUGFxSnntnAABAgQIEDidBM6+57nnXfiwRz32yne8/a0//g9e8NOTs7ixuRNf6n/zWBKjhy/1zU2/+9r3X57/u8UZZ5zxzbO967K3XbIOvW7g9ruvuOztW3F87ctf9lslKH7xJS971W/+2i//u/Pv/8CHPPWHn/O8aw9e86Hf+NVf/PlHPu4HnnTLW91qXaz+ul2+7lW/+9InPOXpP/LCn//lF1/8it/5r3eb1lbPePaPP//sc84975W/81sv2cr77+Hn1K6nuQo9NmuhCoR/PlHbomYDFI+eqJXSGyZaIF4rL46rxc82WVXJUIKgVkCfmWjQeBUiJb9qxdRMhS1vm9oS9en9Q1Uay36+cpTkRxUpJUw6pl7Ta5vnUCVLyYtjbpO05QM/zBPnXHr/Q+ewJC06vpuOYZdWeXS8VVJUCdWsirtNfN/EMxbT9Uxz/rmJ9dqX1OjethEgQIAAAQIECBDY9QISFrv+EjlAAgQIECBAYK8I3PeBD76whMP593vQQ+593wc86MwzzzzrjFve8pj+vXXjDddf/8TvueDsqipud/vbf0tDt//Dz/2rn9mKwQevfu9Vv/lr//4Xfuwn/+ELfvpnX/Qfe82Vl//hpS/8x89/7jXiDIEAACAASURBVCc//rE/nXnbf3m3s+95r8Pt65I3vO41b3n9xa++6GnPek7Rc977nndd/oKffM7T33jxq16+lfffq89ZZlrUVqfkQwv6fXK94eP/aDmnFnsPTtQy6qyJqhQaYt3zPzkL3rtqJsCmxfYGP5eoKDnQ8OUW6ktUdMzHPPh58WjhvMTXX5v41onaO31m3ufL32CfvVcDtvOtXdGVEyUqem1VPbWv2pZtSVCUNOmYeuy/0ZIVu7nN15qs6N4saVGy4gcnahlX0ufA4phh926VFSWlagG2nZU023INvQkBAgQIECBAgMD+FegfvjYCBAgQIECAAIGTJHDrM886q6TDursSFjMb4rbNljirIRG3vd3t5im36fsSGre69a1vfcspe/imSXRc/4Xrrrv6qve8ax1+3c+f/Mwffe4rXvobv/7V2bZ6iLWE+s673PXAtR/9yIcPfugDzTA4tD32iU952ieu/ejB91317nceaV/nXfCAB9/hO+54p4Mf/uD7q8zY6nvu9ecti9gtwtemqEX4O048deLBE9+z6fyqOGkuQAmA9058dhbqj6laYSe81nkVxzu3YkOFRUmPjFo4bwZFZn2K/88mPn+4pMWG1/b3RwmCkgVrlUMcN1U4nOrqhuVad+xds46n2Ro9trh/6Dqe6mM41us/x1xiJevavZ0/UfLseZv2U5Ki/7ZfOVELsJJUJaskLI4V3PMJECBAgAABAgR2TEDCYsfovTEBAgQIECBAgMBuEdiwoN6n/e8wcfuJWkH9vYkfmtjcSqt2O1WxvH6imQz/d+JobZF2y+ke13FsSjrUFqtKibY7T1R58taJT81i/83mtxymndTGv0O+uo2zNA4d8BxP17ljXpMuVXiUdNmxhMUmo/Uara23mvNRG6jHTfz9ieaBbNxK+Lxi4lcnShxVudJA+Rt2W/LluG4+LyJAgAABAgQIEDhtBI6pRcFpo+JECRAgQIAAAQIETleB2j/VSqcF4QZyN7j4wokDm0D6fYmNWvPUGunQIOlZdL7uNBlu/IU53/6W6NP+LZZ3/v2sZMA3b05AbFo0r1poyxVDp+hG7JhLSpW0KMFSxceOHdMRkhX5Vv1RcqhkxXrPbU5WRFS7re7VhqyXPCuhtuurfk7RtbVbAgQIECBAgACBPSxQGbaNAAECBAgQIECAAIG/Emiht0/ct5j97RPNq1i3dXhxC8QteP/YxPdOPHKieQJ37tP7S9uh/W5alcK3LVZ9qr8F9toW7foq7qVtVYv6HXdtk/r6eGd6nOzrnF+2Va50T3VvdY91r3XPde+1bRyk3T3avdo9270rWXGyr4r9ESBAgAABAgQIbIuACottYfYmBAgQIECAAAECe0ygRd9mePRp9RaI++T6sydaSG5rYf5Hl6/PmcfaIb1pooXi5g18bOJmrZH2mMGRDrdKhBbLm5fQYzMsqljofHPb9kqFpUKhD2P1903tu6qO6XhqN3XY81iSFrslSbHxGDv+khW1JOveevTEwyfuujypweVt67342/N11RV/NFFbq42JjCNdQz8nQIAAAQIECBAgsCsFJCx25WVxUAQIECBAgAABArtAoIXfPn3fgO2SFw0y/icTfQK+T7KvWwvJJS96/tkT75947Syi/8V2z2bYRrMSMy2cXzFRy6IGzZck+PIOnXPJiton1S6p61PipDkOa7unbaQ5obfq2KuiqKLi3ImSFmtibN3xeu+VGHrRxH+aaF7Fer4ndABeTIAAAQIECBAgQGAnBbSE2kl9702AAAECBAgQILArBPoU/hE+iV/lQFUWLQj/l4lfmfjsxMFNB96n22vJ0xDnFs7vMvEtk7S4xT5uD9WCeQmBkjolCBrwvFMVC1UlZN5ckRInPR6Y2JhY2hX32hEOYh2uXeVO59E91L3UPdW9tXHr3use7F7snuze7B7tXrURIECAAAECBAgQ2NMCu76/7J7WdfAECBAgQIAAAQL7QmCSDi0kH5jok+93mujT7886zMk1E6HF45+a+MREA7xbzG8g9WFbJR2pZdG+gNuGk1gSQiUm7j7Rdfr8RAv+azuvz+1Q1ceWzn45/tssx9y99Z0TvzTx1yeqsNi8vWx+UBVP99bbJg7O+ZXAsBEgQIAAAQIECBDY8wJaQu35S+gECBAgQIAAAQIEtkGgdjtXL4vE95zHD088ZaKF5o1bC8zFD0y0cF6i4vKJd0zUQmmnKhC2gWhH36K5IVk316G/cUoWtYi/K7yXGRuHA6rivSEbF048dLmfbjeP9z6CZud48UQtyoq/nKiixEaAAAECBAgQIEBgXwhIWOyLy+gkCBAgQIAAAQIETrFA1RG13CkJUQukBk03z6KByD840Sf6163kxndNPH3iquXrb53HhnL3qf8WqZsB8ZX5ZHyPthMQqHpiEgJdmxIULd5XoVBLqJy7Vju+rVU0c5wlVjquHkumVEXRPVRUvXPBxH+f6B5qlsW6VaXzmonuoRJfnVf34hdV6Oz45XUABAgQIECAAAECJ1FAwuIkYtoVAQIECBAgQIDAvhdouPTHJnr8tom/mGjR+fHLz2pN1PDtA4tEC9B3nnjPRAvS10y0sN6i860azD2PJS0KLaOO//ZplkbJoBzXxfy+b67GYV2P/62O7ZVLy6cSFEVDwUuuVFVR+6raWDW0/JnLYzvv3ukeKmHRfdY99daJ/zHxvonPTDS3wsyKY7sUnk2AAAECBAgQILAHBCQs9sBFcogECBAgQIAAAQK7RqBPxbeY3KyKkg39e/qSiQ9O3G/iERMtnl878ZDlqFuQ/hcTL5/ok/ItNNf2p6RFlQAtZLev2v20/xbYd3SRfddob/1A1gqYkhRVJ+R4xCTQ1nd7fM9ckhTrIO3ahpWo6Hi61l3zvm5exWMmnjbRPbJu3TsludpqJdbQ7e637rHaQJXE2BWtro5Px6sIECBAgAABAgQIHFlAwsLdQYAAAQIECBAgQODYBVowLvnQ8OMWoc+bePvERybuMrF5rkBtip4w0ZDk5g48eKIF6JIWfYK+Re0Wolt437joLnGxhWuztEXKaq1W2cKrTv5TlkRFLZ+qjqjypqRF1/eOy/WtsuKciXdOlMTonuje2Lh171RJ8QcTvz9xq+X77rXuORsBAgQIECBAgACBfSsgYbFvL60TI0CAAAECBAgQ2AaBFpDfO1Hi4QETLZr/8USL1pu3Fq0vmihh0fyBkh49tsjejIv21UJ3vy/xUeuoQuufbbiQJ/oWk6wosVCbp+Ls5ZpW7dF8kypqSmz1eNeJElxd8+6Jzdun5gdVVJTc6B65bKKqiypwbAQIECBAgAABAgT2tUCf+LERIECAAAECBAgQIHCcArNQXXKiT9H3yfnaQLUI3ZyLF07cY9lt39f2p39/V03R9usTVVnceqLERbMJWvS+fGJNeLTg3eJ1yQwzLo7zGp3Kly1VFSUl/sbEOii7RMNDJ0o2NeukREWtwrpH/u5yPCUguqZ/PtGQ9rYPT/zr5fsSF1dMdI8csQ2Uodun8uraNwECBAgQIECAwHYLSFhst7j3I0CAAAECBAgQ2HcCy6J1SYs+Nb8uUD9pvn72RAvT9z7MSVeV8eqJFqxbmF4rLqquaD8Nj26hek1ofHq+rl3QOufi0C4tWJ/622mu7+Y3WedTVLH+7RNrQqJ74DsmqpKpyqKfl3wqkVXC6skTVU5s3q6eH5TI+u2J35tYE1jt5/qdHhx+6oW9AwECBAgQIECAAIGvCWgJ5U4gQIAAAQIECBAgcIICLSjPonbJhT4VX2Khheui5EMJhp+YaKZBsQ5Ubo5Bn8KveqJF7FoJvWrigok+qd8sjBbGr5q450TJivZde6CGdO/YUOkT5NrLL+961Nqp+RNdn5IV/U318YkLJ6qY6NpVGdNznzJRW6/7T1SF0TV/9ALQa5pXUrx4osRGQ7VrMbZWVHxVsmIv3y6OnQABAgQIECBA4FgFJCyOVczzCRAgQIAAAQIECBxGYFlYbsH6K5O86BPy755onsWBiRaqawtVpcVzJ2rz9MmJ756oDVCVGP3bvJ+10F0boD6Rf7eJ9nXmRIvjDev+xMRbJ2oh9fl5ry/Pe5cUsZ06gZIJ6wyKKmgePtGw7BITJZG6Pg+b+OhECaiSTt0LT5tYh2iX4HjXRNe+9lGvn6iyonZQfzRxcHlu19uw9VN3Le2ZAAECBAgQIEBgFwtIWOzii+PQCBAgQIAAAQIE9qbAUnHRwnNVFi1gtyDdIvR7JqqOKCnRonefuq/qYv13eZUYffK+n/XJ/KoxaidUe6j2V5uhkhO1D2p485q06BP5LYzfrOpCy6ij30OHafnUi9Zqiq5N17H2TiUr8r/TRAmkkhXNLKkNVNeq31Up87eW79tPr+96dq275u23e6B7oYRHLcG6R26Y6DpKVhz9knkGAQIECBAgQIDAPhWQsNinF9ZpESBAgAABAgQI7LhAyYMWomvzU6uoKiaKn51o4fr7lyMs8bBuzasoKdHPSlw0w6CkRJ/wbzG7odxVafT9usD99vm6BEa/7716bNizhe/juwVKKORckqJWXD02h6QkRF9XTXGviZINJSn6WRUTVVBUWdHPqsbYuK3X+A7zwz+YqEKm61ayoig5pcXX8V0vryJAgAABAgQIENhHAoZu76OL6VQIECBAgAABAgR2n8AykLsEQx8W6lP2zT/o0/n3m6jl0yMnaifU9n8mSji0KF7roBbB1zkYJS/etLyuKdAtot84cXCiVlIlMGo51Kf5m3NRssQMhC3eEst16u+jrlHuzZZ40HItqqg4MFFCqeRQM0eqmmkeRQPSu74lmnIvedG1KJFRgqLt0om3TNQyqtdVmVGVRdfoZoPUl9ccelAhs1HD1wQIECBAgAABAvtdQMJiv19h50eAAAECBAgQILDjAkvLof7t3SJ2i90lFaq26LGF63878X0TLV6vVdBXLF/Xiuic5ST+2zy2eF6iokXxKilaBK8Ko2HNzc0oAfKnEy2Ml+Rony18q7g4zJ2wJCr6Te4lH0okVRFRguEBE/eZqBVUyaUqL0omlbgoSfTMZZfNHKllV9a18Gpbr+Ub5uufmShRVRKkiooeSzpd77oc5qL4EQECBAgQIECAwGkrIGFx2l56J06AAAECBAgQILBdAhtmJPTv7zVx0aJ37YOaeVCLoRbKHzrxiG9wXLV8qk1Ri+EHJxrAXaKiGQrNT7hyosXwayZaEK+tVAvr/a6o4sKA7qCu/X9VRXQteixKBHU9SijdfaJk0gOX3zVDpMRFg7YPTJTcWK/FfHnY7ZL56eUTJY4+MFHbp65HyaZ1VkXX40iv93MCBAgQIECAAAECp52AGRan3SV3wgQIECBAgAABAjsoUJVDUTunFq177JP3zS94/8TVE1VO1EKoyornTaxDmWsv9MaJEhb9O76F7yovWvFuPwcmqgJoYfxjE7WU6pP/LZxX2VGi4uOzUN9z13kJh6ou9vun/DdUUawJo2ZM1NqpBMU6H6REUZ61dPquiRJJtYY6OHGPiYZrVw2z/g3Vtci1Nl61kapi5iUTVVrU4qtqmKsW91pF9dp1tohql248GwECBAgQIECAAIFNAhIWbgkCBAgQIECAAAEC2y+wJi5KOqzzDGo11IJ6vyvhUGKi5EOL3e+ZaEZCi+Hr1qf9a2FUdcX7Jlpgr5VRiYkGc1d9cd5E/+Zfqzka9lwiowqNEiMNjv7fs6C/Hs/6eNOb7IUKgA0VLBuv5JqcWB9zuv1EzpmUmGj4+Vr18MT5OtNirbzo+bnmuCY51vfoWlRB0YyR+0/ULqpWXFVetM8qX7ouOX/DORUbD9rXBAgQIECAAAECBE5nAS2hTuer79wJECBAgAABAgR2hcCGwdx9Yr/ok/33nTgwUeVFiYSfmKhN0XcvB/3heWxxvdZPJSSq1GhrcbyZFn2av8Xykh19+r/qi5Ijl03UOqqF+NpHlcRo67nNvOjxK3u1ddTS6qmqiRITJXR6bCs5kV9JoFo95djw82aAVMVS0qHnlnhoZsX64a4qI0osVclSEqhqi7Yc83vxRH9XnTtxcOKPJ0oyVUFTZKmiYkHzQIAAAQIECBAgQOAbCUhYuD8IECBAgAABAgQI7LDApgqB/o3ep/lrM1QbohbK+zR/i94XTpS4qDqgmQu1NaqNVImIqgB6ftt1Ey2+txBftM9aQZW4aNG94dwlO0pmvG35+VoxsM52qBKj9zw0+2LZx7L7Q22U1t+tz1+rM9YqkUOtpkrGHG3BfknYbHyPdR9rdcTm99o4h2N93Xoc2azPbyZIrbUy+N6JkhKdf8O0O/9+nmHPz6YoYZN926cmqpIosVHVSobNBMmmRMU7Fpfeo8RRz8/+y0c752X/HggQIECAAAECBAgQ2CAgYeF2IECAAAECBAgQILDDAkdoadRRlbhoMXydQdEn/5tl0YyF8ydqc1SrqBbLqwh40kQVBG1VXLSA3r/5W4CvdVEVBiU3SmzU7qgZC0UVGlULtABfIqSKgtdONOuiREZVGz2n6Gcd17p1TB1jC/0t5Ldg3+tLIHRMJQT6WRUfbevfIGvVQRUNHV/JgLV1Uu/Tz0o+lHjpGKoaWbf1GHqfovfpGDquiyZ6fYmFEjydc8+5YInaYOVSEqJzzq/j63jWORW9TxUov7ccU0mj/Bq+/ScTtexqdkXHtM7A+PwkKTouGwECBAgQIECAAAECxykgYXGccF5GgAABAgQIECBAYDsEluqDteqihfkW8EsC9Nhie5UCJSlqVdQchpIbLdjXAqqF9Z539+U5JStanG/YdPsoQVAbqPbb4n2VCyU/Sjy8YqJF/FoiVZVQwqEKhNos9X2L871HSZMDEx+YuGKihf4W80se3Gf5vueWQNi8oN9zSpD02Dk096HnlJTp+4dM3Gvi4ETJgto39dzOueOuQqKER9+XoMnphyZKdJRkKJlQwqLz7Lg7zxIjzZgoIVLSouO9ZqKES4mg3qMER+2cLp6o9VbP6ZxLWvS89rHOpjg0wFxFxSjYCBAgQIAAAQIECJyggKHbJwjo5QQIECBAgAABAgROpcDSVmltcbTOpWjBvIRDQ55bYG9xv1hnULRQ/9SJFvBbUK/6oGRECYcW9ksMlGxoob+ERkmKKi56Xgv96+J9szRKHrx6OccSHy3kV6XQ60qSlBypMqEF/cdMlGAokVDipIRDx9Vzel2Ply77aqZE79PzShCUFCjh0fM6zhIgHXP7bh/9vucXtWfqdSUa2p48UZKk2RG9tsRD51JlxjqTIpOOMa8SKdl0HiVwavtUIuTgxCuX9+38+r6ZFL13z883+67DobZUe2EoecdpI0CAAAECBAgQILAXBCQs9sJVcowECBAgQIAAAQIE/kqghfIW7VvkL9HQ1mL65RMt+Pd1i/lVSZRQaLZFlQRVGVRt0OtbxO95BydKWpQQqbVTr6vy4EMTVSk8YXlNCYOSEA+aKDHQgn+JjZIZJRj6fQmIkh4HJlr8LxnQYOvea+O2DgcvubFxKwnQPttHSZaqR9pHr++5HdvDJjrnvu69SySUoHjsRBUir5noXDrfkiM9r3107iUr1qHaVZ6UwOg1/U1UxUVJi6opapHVOa0zOUpQrO2o1p/Nj2wECBAgQIAAAQIECJxsAS2hTrao/REgQIAAAQIECBDYQYFpIdVCfNs6B6L2T1U6VJVQMqJF937WQnztnkpK1G6phf9+VmVDVQf3nKhaoue/a6J5EC3uf3CihEQVGiUTqjooEVKciq2kQlFLp5IaVUiU0DhnokREczdKpPS3TcdesqXz7NirQinRUtuq102ULOlnJSh6fufZ0PISPf1snb9R5cTGwd6n4rzskwABAgQIECBAgACBTQISFm4JAgQIECBAgAABAvtYYElglFhowb+kQlUJLfZXpdGi/DMmav1UC6USGCUtSkZUnVFFQgOq+3mVGmvlRM+piqFkRgv9tWBqa8G/ZMHJ2Dbuq4qIkiz9/dIcjpIOayVGlRElImod1TlVJVFSo+f089pC1SrqdydK5nROJV2qCikRUsLlixIUJ+OS2QcBAgQIECBAgACBExOQsDgxP68mQIAAAQIECBAgsCcENgzvbsG+Qdct6B+YuO9EyYEqKB4wUfuj2i1VcbHOfegcS3j0fYmBXttW4qJF//bXVnKj35+MbeO+GthdsmXj+/b7Ei4lHNpqbdX3VVTUtqoWV++eqAKjJEqzKA4ux9z+Sm4Yln0yrpR9ECBAgAABAgQIEDhJAhIWJwnSbggQIECAAAECBAjsFYGl6qL2TiUBmlVRkqIF/mZF9PWjJh48UeKimRFFlQvrcO+SHM2nePNElQ8lO3pdf1+sraUuma8fv5jUuulI8/M2/u7353mPmFhbOa2zNUo6VMnRcV02sQ7CrlqkSpBmXxQlKt65HFfn8z+X4+rrZnqUXPmSaorlqnggQIAAAQIECBAgsMsEJCx22QVxOAQIECBAgAABAgS2S2CpumjWRa2eaglVdUQVCj3WAqrB17WDaqG/ORhVWTQjouRBA7BfO1HyouRG1Qw9p3kSL5t478QTJ6qA6PUHJqps6PVtzcioMuPgRImT9n3xRAO9nzXR3IxmS1T1URKiJMVFE5dOlCTp9e275/T62j99ZKIWUVVflDjpsZZQzby4cRIVJUBsBAgQIECAAAECBAjsUgEJi116YRwWAQIECBAgQIAAge0SmMRFb9XfBlVBFM28qHVUP2vQ9Y0TJQjuPlFbqM9NlCT4k4mqGkpslPAo6VACpKRBiY6qHvq+6ov229fNoGireqN9V2FRBUTv0YGUeChZ0vclJEo4lIjo+edPlPxofkXtn66ZKAHSfjvmEhK1elr3WzWFJMUC7oEAAQIECBAgQIDAbheQsNjtV8jxESBAgAABAgQIENhBgaV9VEewJjFKBvR17ZhKJjT/or8rSnAUJQiqaOh3JRVKcPR9P+/rfta2ft1rq/BYn1vio+/7ecmHQ7MmJppD0e9qS7Uew5qcaH/rfpfdf+1hEhZf971vCBAgQIAAAQIECBDYvQISFrv32jgyAgQIECBAgAABArtCYEMFxlqt0N8RxaHvq2KovdRazbDx662cwLL/9ak37XfDe6x/t6y/u+k4VFBsRdhzCBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgiH63eAAAA4NJREFUQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBAgQIAAAQIECBDYksD/B640zyYHlIM3AAAAAElFTkSuQmCC"}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO3deXhV1b3/8ffe+8xz5jkkJCQhgTDJPCjiBKLWi9o61qpXr6W11tk6Dx1oa9tbvT715231arXOdaooOKEogoCiAgKBQOZ5Tk5ypvX7I3ggEvVQgWD4vp5nPXL2dNY+x/PJHtZeSzOZTBuUUqMQQoivoGlamWYYRk84HLYPdWWEEIcvwzD8+lBXQgjx3SBhIYSIiYSFECImEhZCiJhIWAghYiJhIYSIiYSFECImEhZCiJhIWAghYiJhIYSIiYSFECImEhZCiJhIWAghYiJhIYSIiYSFECImEhZCiJhIWAghYiJhIYSIiYSFECImEhZCiJhIWAghYiJh8R1x5d33c9S4oqGuxn5JyS7gxl/+gdKxxUNdFXEASFh8B2QUTOCUk+eycdPWoa7Kfll84x188PZyrrnzt/I/2jAg3+FhT+fq235DoL0RfzAy1JWJmW71kuxSvLV8KfVdkBzvHOoqiW9JwuIwN++Mi+mu3U5La9M+8/JLp/PwC29y7NzZQ1Czr5eWU0B9RRkA3V19uOyOIa6R+LYkLA5jroR0fnTh2Tz4vw/S29GNLy5+r5LA4htu5cmHHuDMCy760rz+YrPZhqzuKWnpNNXVAWCzm/AHAkNWF3FgmIa6AuKrLf7Fr3jsz3cSCCt8Gbnc+Ks/RueZbS5K8jIILjiNwtJJA+Z94aN3lvLEP544lFWO8sTH097eAkCCz01rW8eQ1EMcOBIWh8BF1/6Sho1v8/Iry2NeZ+Ixp5Fi6eTVZW+TVTyVsg0ruf7qG6Lzc8fN5kdnncBdv/4z/++vD3D95T88GFX/t7kcbvxdjZidCZgDbfQE1VBXSXxLchpykBUcdSwTRiXxytLYg8LuTuCKq67gt3feigIM3UwoEBqwTEpqGg111fiS0mhvqj7Atf72LDYHgb4gJUfNYPP6VUNdHXEASFgcZBOmzmL5808T2Y8/rItvXsKzDyyhrrE1Ok2pgRtwuL10t3eSX1hM2ecbD1R1DxiTzUwwFGTuiQtZsXzpoMskZxdx/c03k5pbzHU33XSIayj2l4TFQVa2+VOOPeV0zKbYPuqZC84m0dTGy/9aFp0WUWEsNjtZuaOYPGsuC/7jLDweB4FwiNKjpvLxhx8crOoDkJiRx/yTF+wzfdKck8hITRx0HZNhoNs8TCjO5sP1nw26TFtjNa+/tozW+ireWLZnf802F1fe8ku8LvuB2QFxQBi6rt+klDIPdUWGq9ryLSTlTeTn19+I3WYlHA4TDAYIhUJEInvaTZjMFvLGTuGu3y5h2UsvMPWYEznlzPM455LFnHbGmYwsKCY3bxSJSUmEg330hjSceogpR8/j4f/5E8Hwnm1NPvokvHadpqbmf6vONruDUCgYfT1u5ol8/4wFvPziSwOWO3fxL+iu/pyK6jp88Qn0+f171plxLDPmHMOaZc+w/qNPBn2fcChAXV0dXo+bHdu3RaefesEVzJt3LG01ZZTt2DXImhojC0sIBXoIBIKDzBcHmq7rIbnAedApHv3zXSx9OptjTljAWT9aTGp6Oi63B5PJ6F8iorA53TitOm8uexWb08Wusk2semspNZUVaJ4M7r7pCq6+7LLoVqccfwbH/mARTTs+oqdvz/WMkqnHc8U119NZX8aPL/lPRpYcxbW33sF7Lz/G3x99nKxRpVx3+93Ubl3Lr+64M7qeyerkv665mZaGWhadcz5vPfcQ9917PwC6YZCWNRKTrhHa63yqqGQsHzyjccWd9zGptJD68k+57udXAaBpGqVjCrntJ+dzwpmXcOnll/LoH2/jhZf2nJKMn3kCV15/A10d7bjsZn563vfo9Icwm3SS0jJYfNufuOT6Xm74zzPZVl4VXe+ym35PcW4S8UlJXHrmQvyB8AH+zsSgDMPoAZSUoSujxk1Xj73yjiouzB90vtmZoh5+8skB01LzJ6oPttWqCWMK9kzXdHXv06+rSZNnqAf//oiyOLzq4ZfeVgVFxeqRf76iLE6fevSVd9WY4kL1l2dXKJ/DiK573e8eUueec5a64Mq71MIF89VjL7+pDA0Fmlry0EvqL/94SZ2y4Pjo8onZo9V72xrVjXfeo26/6w4FqN8/ulSNSI1TgLr4hiXq0ssuUiPHTlN/feIZlTNmmvrDn/60p/65xeqR519VCXEeBaiU9Eyl7bV/dz7wnCrJz1QXXvMbdcLcmdHpFneSeuLl15QO6g//WKYyEtwKUGOnzFEJce4h/y6HazEMo0euWQwlTWfB2Zdyyx23cfPl57BpS9mgiwX9rZgcCQOm1Zd/Rnn5DrZs3RGdNmnu9+ir2sCOmjZCfj9nX34dyx6/j+3lVYRVkO9fejVvPf0An23agmFW9PX1/0UeWTqDWROyeezxp3j/7dc4/fyL0HQdi9nEwvN/gt6+jRuv+hmLLvwvtN3v9b2zL6SuchfzTpzHf/9uCQBtre04HQ4sDi/zTzmV8vJyrr71Ln5701WYzBY6u9ujdb3s2tt57an/pbm1g5HjZnPV1Vegds/LGDWeEYmweXsVaZkZ1NbsOapY9MPLaWuoYczME3EG6qlp7sSwOLjmtrtRYTnCOJgkLA6CgnFTSE9N/tplRpVO4Q8PP8fkMbksPvd0yndVffXCkQCdAQ2Pfc+lJRUOsPz1d1l01iIAnL5krrzmKu79/RKsTjuGM5G5M8by9FPPYlicuNw+Tpo3jccf+wcAZkMRioDF4eHaW+4gGIygAWUfr+SpF94gM2sEDz63nLEjE7nzpptorS1HcyRhNevkFE9mYlEa765ay9JnHqWrpw+TzcXoURnsqqnnP6+7G4cpzOyTz6F+4zts2V6BAgy9/7Rr9inncdzcmXS09t/tWbDo++QV9D+ZarI6uP7OX/Hnu24hosDhdOL39wKQWzKZ+fOmk1I4lUsvPo+br/opCrjgZ7ew8p9/o6Wj59/4tkSsNMMwesLhsFx2PoCKJs3mpjvv4oPX/8XKFW9SU10Nmk5SagZjJkzmmBMXEupq4qH77uGjjzfEtM0r7rqfdS89wHtr9ixvc8Xxp4eeZOem9RRNnM5T99/NK0uXM2LsdJ785/PcetkZLHvjXRyJeby15gOWXPVDnnv+FQBuuOdh9O4acoon8cLf7mHE5JOJNzr4cN0nLDzrfB7/8+2sWr0eiyeZvz3+JJs2biYtzsyTz77CBRf9iF9efyX3PrWMdSteIyHOhe5MZsf6N4m4s0hzh/h0ZxuXXnw+Zx83heqGViyOOP727It8sm4tJaPzuf/e+7ni6qvYvGUHHpOflpAXe7iF5JxiVvzzrzzxxDMAzD9nMSfMHseH6zdy8ve+x+0//SGjpp/CycdNZ9nSpZRMPhqvuYebrvr5gOsp4sAyDMMvYXGQWOxO5hy/kMnTZ5CSmgpK0dxQw+effsz7b79OdXXNfm0vr3Q6hVleXvnXqwOmmyx2JkyZRn3FNioq+o9OdJOF0vHj+HjthwBoupmTTj2NZS8+S3j3D8psc3DU1BlUbNtIdU0tmmYw47gFZKansOad5ZSX77kLUXzUbM485zx8Hjeff7KGJx76X6YvvIBbbr+Fn/3gODxZpZwwfz4GYd5d9iIvP/88dk88GakJbN2y57H6pPQR5Oflsn71SvoCITJyCkhNjuOjD9eAYWbStFk0VJaxa1fFXnuoMeO4k0lLjuetpS/Q0tp/KlM0fhrjJ4ynavsm3n/3XSJKguJgkrAQ/yaNB/75Jh0tDTz2x5v4+LPBr7WI4cMwDL9csxD7Lbd0Jj3Vn9LS0Uco2DvU1RGHiISF2G8nnPIfvPbCM1gtDgL+vqGujjhEJCzEftKZMXMqK999H7vbRnePhMWRQsJC7JeknBL8tZ/T1RvC47DRvVcTbzG8SViI/TJ20hQ2rP0A0HE4zHT75dmMI4WEhdgv+YXFbN30KYbVhRHo5DvUh7D4liQsxH5JSEmhtqaa9LxianZ8PtTVEYeQhIXYL6FgCF3XmT3vRFateGOoqyMOIXlEXeyXla8v5Ybf/42+nnYWn//Loa6OOISkBafYbwkpaXQ0NxAMyVOeRwpp7i2EiIk09xZCxEzCQggREwkLIURMJCyEEDGRsBBCxETCQggREwkLIURMdKWUBIYQ4msppQxdKaV986JCiCOZUkqTowohREwkLIQQMZGwEELERMJCCBETCYsjmSbXtkXsJCwOYzl5BYydOBm31/ettpNXMBqr1caoohIMo39w4oysEYybOIWScRP3Wd7ucDJp2ixGjBw16PYKi8d+7fvpus6oohLMZgsFo8d8q7qLw4eExWHM7fGy8eN1dLa3xbyOrg/8SvMKi2lpbmRk4WjqaqoIh/d0WBNRETZuWI/VaiM1Iys63TAM2lqb2bVjW//2NA2X27NnvmlgB2val26qjR47npqqXYwuHU/Fzu0x110c3iQsDmM7yj5n5KgiAJJT07Ha7NgdDqw2GyazmezcfDxeH9k5eaRmZJGcls68+adhdzjJHJFLQlIKBaNLcDpdZOfkEQqFottOTEll+5ZNJCanMmn6LJob6qLzujo7cLrc2OwO5i04Dbfbg2EykZGdg9PlJj1rBBarlezcPBKTU5h74slYrFZy8gtISEohK2ck3rgEMrJyCEtvWsOGoWnaLYAx1BURe9PIzS+goa6WrNyRhIJBxkyYRFx8AlarjfGTp2OzO7DbHRSNHceu8jLSM7PZtaMMs8WCUgrdMEhOSaW1pYWK8jIsNhs1lf0jo1ttdhxOF031dWSOyCUSCVNbVQlATt4oOtrbSE5Np7mxHk0Dq82GUgqH00U4HCY9K5vGulrSMrOp2Lkdq82G3elERSL44hNoaWqkuamBrq4OWpoah/KDFAeIpmkRObI4DNnsNkwmM9B/WpE7qgi73UFbSzMeXxyd7W0kJCbz+Wcb+n+YjQ00N9STmJRCMBgkISkZXddpbKint7cHp8tDU/2eI4dAXy8ut4dIJEJDXQ2h4J6BghKSkolEIiilSE7LoK6mGpPJTGpGJju3byUtM4uWpkZaW5rp6uwgKTmVlqZGXG4PVpsdf083zY31eH1xNNbVHvLPThw8cmRxGAqFQsQnJpOcmkF1xU5cLjebPvmIYKAP3TCor6mmt7eXSCRMe2srPd1d5BUWU7lrB2npWTTU1WB3OAmFgnS1t5GQlExdTRWRva5X9Pp7GDmqCKfTydbNn6GUAiAcCpOVk0tPdxdtLc0kJKcQCgZpa20hc0QOTQ31dHd2kJSahscbR211JYkpqXS2txGJRLDZ7VRX7CQjO4fa6sqh+gjFAaZpWgRN0/oAJWX4lUnTZipd19WkabMO2XtOnDpTAWryjDlDvv9SDlzRNC0g44YMQ7mjCnF7vMQlJFE6cQrNjfUD5jucLnq6uw7oexaNKcXucOKLi2fi1BlU7tpxQLcvhp6maVqfUsoy1BURh4bH68PmcNBQWzPUVRHfIZqmBeUC5xFm5KiiARc7hYiVhMURJn733Q4h9peExRHG6XQNdRXEd5SExRHGGxc/1FUQ31ESFkcgu8M51FUQ30FyN+QIk5NXwJgJk3j5mX/sNVXDFx9PXsFoXG43Lren/zkSBYbZRE9XF73+HrZv+5ymhnqUXPM44miaFpR2FkeYndu3cvzC72E2W/DFxzN2wmSmzZ5LXmExtdWVhEMhEpNTcLrdBPr66Oxop6e7GxWJkDkil107ylj3wUo+/nAVtdVVhMOhb35TMSzIkcURxmKxcuGPr2Ti1JnEJyRSU1XByjeXs+a9t6mpqiASiWAymVGRCKFQEE3T0HZ3kpOUksakaTOZOmsuhSVj2bWjjPfeXs7r/3qB7q7OId4zcTBpmhaUsDiCFI0Zx8U/uZrE5FRCoSBP/t+DbNv8GTVVFQQDgZi3YzKbyc0vZM68Ezlqxmx03eBv993Dh++/I7dlhylN04LybMgRUExmszr3ksXq6eWr1BnnXaQyR+Qql9ujbrj7HnX08QuUruvKMEwKULquq+S09Oi6bq9P6boefe31xSmL1RZdNiUtQ5102pnq8VfeUT+94XblcLqGfH+lHPiiaVpAjiyGOYvVyrV3/Jb8gtHccd1PqKncxcJFZxOfkERXVwe6bvD8E48wcepMpsw6mleff4aK8jK6OjuA/qOIcCgUfSpV13WUUtHXX0hOTefqW3+Fw+Xm5isuob2t9ZDvqzh45MhimBfDZFI/vf42teT+h5UvLmHvvxLKbneojOwcNXrseHXiKYuU1xen3F6fuv2e+9W4SVOVpmkxvYfFYo3+2+5wqCtvukv95n8eUja7Y8j3X8qBK5qmBSQshmnRNE394MLL1G/uf3jQU4PMEblK13V16pnnKofTpUaMzFeapimX26N+9os7ldvjVSaTafe2dGV3OGN6X7PZoq644XZ17e1LoutL+e4XTdMC0ihrmMoaMZIzL7iE+5bcMejj6HXVVf13Psxm4hOTcHu8eH1xeHxx9PX2Eg6Ho312KhXB39MdXTcxOQWT2Rx9bbZY8PjiAAgGA/z1vnsYd9RUJk6deZD3UhxKEhbDkKZpXPSTq3nn9aVU7SoHwBefMKAX7lCovyu9V194hjPPu5hgMEhfXy+JySm4vd4B4fBlLc1NhIJ72lcEA4EBy3d3dfLUIw/y42tujnYPKIYBOQ0ZfiUlLUM9v2K9SsvIik4zmcwDlklMTlWJyakKUFabTZ146iJ12c9vUGecd5FyuvY9bdENY9DrEPGJSUrTNKXtdccEUA6nUz352vtq7MTJQ/55SPn2RXrKGqYWnH4WWzZ+Qm1NFVk5I6mu2NXfwErXo021O9pbo3c0+np7ee3FZwGwWG0Eg/u2uVCRyKDTu7s6UUrh9nhRkQhdnR1omkZPTw9vvvoiZ11wCZ+u//Ag7q04VOQ0ZJgxmc3MOX4+Lz79GChFdcVOIpH+jnqTU9OjI5IF+voGPUXwxcfjcnswTBYsVid2RxyabqCUIhzat2l3X28vAJ3tbdHbrQApqem89uJzlE6cgtvjPRi7Kg4xObIYZlLTM4mLT2T96vcBBrSorK+pGrDswOsSGi5vAjZ3JvFpyXgSMrC744iEgnQ219DasJOmujK6O/cdB8QwjOjwAQBKKTy+OBrqaqirqaJ00hTee2v5gd9ZcUhJWAwz8+afyifr1kSDwDCZBj0i2JvTnURO8QSmnxFHKGCmblsBkYgFwzCh6QY2Txw2lwNfQha1FZ/QUPM5JrMZh8NJR3sbmqah63p0aESb3U5eQRFx8QmsWvEGxy88fb/DQtN1EhKTaWrYvy4ANU3D64unrbV5v9YT30xOQ4YR3TCYccxxvLXsX8C+QWGx2r60hkZi6ijGzfoBI8YcjcWlsCdUYHE1oOsG4VAQND+6dQfZk1rImQQ5oyfjjc8gFAzSsXsM1lAoFA2K3PwCTjnjHKoqduJwuVi3+j1KJ07BsZ89dBWMHoPL7d7vz8Dri8P5b6wnvpkcWQwjiUnJ5OYXsGHtaoABQWG2WJgweRqrV74dnZaUXkDJtNMxO+z09YT4dPkIND0TlzcTpfpvrZptrSQk22hrdFEyr5awCtLTfhR9/k56/XuuUVgsVuadfBqB3l6efewhNE3HMPqvdUTCYQpLxvLRmlUx70vWiFxWv7eCuIQkOjvaBoya9nWS0zIo37alfxs5I4mEw1TvHrZRfDsyItkwMuvYE0lNy+SZv/8VTdNITc+MXnSMhMPRsU4BzBY74+acTGqRjfzpmzCsVYT7RkLEvvsHHuq/q9HZQDhcizOxAsMUJiXfoLujE1O4CIslREZWNlarjTnHz6ezvY3KXTsoGjOe9MxsfAmJ9PX1kp6ZRUJyCmtXvRvTfuTmF9LX20tTQz2Tps6ku7OT/KISps48msSUVJRS5BUW4/Z4KSoppaW5kYWLzsYwDFxuD3kFo6mtqiA9M5v4xGR88QlkZI3A5fGSnZtH3Zeu3YhvJmOdDjPZOXm0NDdGH/Rq2j24kMnUfwCpaRrW3acivoQsRs1oJmPMOoKBTly+LLLH1WO2OTBMZiw2B874MJg/JEI7XS1B6rdlsultLyZbGLsvhL9XUVhSitPl5tUXnuad15cyefocdF3DarOx8eN1NDfW09hQz4jc/EHrrGkavvgEfPEJAIwsKCKvoAhvXBxZObnU11bTUFdDwegx1NVW097ait3hZOf2rdjsdrq7u7BYLOzY9jmhUIiUtAyaGupIzcjCZrPjdLlIz8xmw7rVjBxVSE1VxSH4JoYnOQ0ZRqw2G7q+VyvN3YfuvvhEmhrqMJktJKakUl25i8TUPOy+LqxOneaKNFp25qGbVH9HN5pOJBKmqbIexSj8gXx6/RVkj4ngS7FgtiUQ7GnDV5fNlo2f0NXVSaCvD4CqinJ2bt9GXEIi516ymPraKlLS0rHbHdFOdMxmC26vr38E93CYivIy2ttaSUhKwW538vorL2C12cgcMZLk1GQ8Xh87t2+NNk/v6mynoHgs27dsonTiFJSKYLPZqauuorxsCyazmfTMLLq6Ogm3thAMBlFK4e/pwd/Tc+i/mGFCHlEfRn58zc344hP41S9+jm33j3OwZts2h48xU+eSP9uPNymB6s9KiYTMaFoApaygFOGIH4ujntTCXfR122mvTcXfXU3m2FrKPuyhobwHc2g0FWXvEA4Fo6c7SSmpzD3pFJ76vwcBSEhK4fJrbiK/sJgH/vhrDN2gr6+X2qpKGuproiGzvzRNi96qHT12PFs2fTpg4OdvWkfsH+mDc5gxTCZcbg/Qf1dA1/VBw8JidWCxhzGb0wkH/UA3zoQO/B1WVDAJNAPNqCFr/Ga8KTqRcBcWVwXrX0zGnWjCbp1OSqaP1sqtdLS1otSethxNDfXs2LoZ0ABFc2M9ddWVJCalsGrFGwdsX7/8o/+moBhsHbF/JCyGkV5/T7QRVn1t9YB5VquNUDhEJBymr7cLf4cNtD66mzMwO3poqbZhdyahIgo0ha5lUb9jM5oWxJNkJqPATfD4DnasKUDXvFjtrkF7+VZKsXbVyoHTIgq//6sfTPu2vrj7IQ4uucA5jLQ0NWF3OAadpxs6Ho+XojHj0Ajj7+yk/vMSulp0CmdvwJf1Bt0dDaBpKBVBKQsd1fOo+mQcjbsChEMRUvM1wqFOnN5EAv4uenvao0cVhtH/d0fX9ei/v2B3OGhp2rfl54HS2+s/aNsWe0hYDCMb1q2moHjsPoMI2ex2Ro8Zz8mLziYnv4BjTpiPCrfjb2+ivakNf1eQ5FwLhXM+I6w2ousGmqZhGBaC/kQCPRba6v1Ub+nB7hxFJBKhp62BtuY9dxZ88f0jnem6Hr37Av3XCcZPnsb6D947NB+COGjkNGQYqdq5g77eXorGjOOjNe8zdsJkTvv+eQQDAdatfo/lL/+TluZGTjnjXFqbq3AnNBPvK6RqYxXTFpkwzDpNuzroqg8RDPix2JxomhlXvA/d1IDVbga9GX97Hz1tjbQ07mm30dzYAPS35gzt1RgsNT2TjOwcPvt43SH/PMSBJWExjPT2+vngnTc49qSFzJp7PPW11fzlj7+m1+8n0NdLoK+PeQtOIyklBRUJUlfxKRanl7isPPp6tlO2po/26pmYrSZMZiu93e1omkblx6PJHNdMb2cKDk81VeV2KnesJRz65jsZpZOmsn3LZhrqag7BJyAOJgmLYWbr5o387Bd3cN7Jx1BbXYnd4aTX34PN7gD62PTJelateAN/Tze60YzHl47VE2bnhk62rizCm9j/OLlhsmB3mlEqQm+nn84GFxVrzbTV9VD++Zt0ddTjdLn3GVzIarWh6Rq9/v7rCPPmn8LS55+WOxHDgITFMHLCwtNJSkmlq6Mdp6v/Yaovbp1+8d/aqsro8uFQgLJNbxEMTqNlZwruJA+9HS1EIiEC/m7s7nhQivaGCmq3GLQ1baS2ciPhUB+6rjN9zrG8vfyVAc9t6LqOtrthmDcunpJxE/nvX992qD4CcRBJWByGDMNg2pxjaWqoo76mZsDj1rn5BZSXbd1nnWmz59Lb6+ev9/6epORUTj/7h/zu9uu/8b00LUxjzQZ6e0O43InYHF4Mk6V/fJCIoq+vi+7OJro6GomE+0NhwpQZbFj7AW8sfXGfIwa/f08LyXnzT6VyVzk1ldLEeliQPjgPv5KQlKySUlIHnTdmwlGDLl8ybmL09eix49XTr6/+itHBBo4HYjKbldvjjb622mxK142vrd8XwwjsPc3pcqvE5JToa8Mw1P88+pw66bQzhvzzlPLtiwwFcJhK2/20ZHxiEiaTCW9cPGaLhcTkFHRdx+P1YbXZgf7DfrvDycYN66Prb938GU31tSw4/ax9tj1p2kwys3Ojr0PBIJ0d7dHXwUBgn/4gdN2gsKQUAKfLRVXFzn3GNO3199DVuef6xYQpM8gckcuK5Uu/xSchDicSFoehcCjE9i2baWtpZtToMRQWj6WwpJT8wmK6OjsoGTeJzOwcACK7+9n88vqPPHAvi879UbT5t6bp5BcV88m61dTVfvUj2pFIhM72NgzDwGrrf0JVoUhOTUc3DPKLSvB8qU9N3TAIh8P07j4FMUwmzr1kMf946C9fO6SA+G6RsDgMBfr6CIWCRCIRvL441q5aufvHaycUCOL397B96+b+hQcZdxTgw/dXsPGTj/jBjy5DNwyUilC5s5xgMDjggmRicgrTZs/dZ32PL47c/ML+t4hEePeNV4mEw2xYuzraQxb0H9nE7X68HABNY95Jp2KxWHjp6ccP0CciDgcSFocZwzBITEmlsKSUnPwCKneVE4n0jw6mULS2NoNS6MbX91cUCoW4b8kdjB47njPPuxhd1+kbpFl0R1sbtdV77pDYHQ7MFgvBQGDQJtq6rqPre947EolEG2QBHHP8Av7jnAtZcuu1+9xWFd9xcoFzeJeM7Bz195ffUlfceIcymy3fuLzb61NWq22f6RaLVVltthik/k0AAAIWSURBVP4BhQYZNFnXdXXm+RerZ95Yo8ZNmjrk+y3lwBZN0wLSn8URICUtg+vv+h26rnPvkjuoraocdPzTr2Mym9F1fZ/+J6w2G8mpGVy0+CrSs7K5585fsHXTpwey+uIwoGlaUMLiCOFwulh07oWceOoZfLz2A9asXMGGdatpb235t7bndLkpLp3A5JlzmHH0cax9/10e/sufaGuRLviHIwmLI1DWiFx+ePmVFBSPpaerk7eW/YvV775FdeUugoF9hyfcm2EYpKZnMn7ydOYtOJWk5P4u+h554M9s/mzDoP1biOFBwuIIpWkaCUnJTJo2iymzjiG/sJimhjpWvrmM7q5OHA4nbq+XSETR3dlBX18fuq4x45jjyMjOpaZyFx++/w6rV75NXU1VTL1Uie82CQsBgNvjZcyEozhq2ix88Yl44+KiAaAbBh3tbXR3dvLx2g/4aPX7tLY0yYNhRxgJCyFETDRNC0o7CyFETCQshBAxkbAQQsREwkIIERMJCyFETCQshBAxkbAQQsREwkIIERMJCyFETCQshBAxkbAQQsREwkIIERN9dxdpQgjxlTRNi+iapkmPJUKIr6VpWkROQ4QQMZGwEELERMJCCBETCQshREwkLIQQMZGwEELERMJCCBETCQshREwkLIQQMZGwEELERMJCCBETCQshREwkLIQQMTFpmlZmGEb+UFdECHH40jRt+/8HK8lWxAMyFzUAAAAASUVORK5CYII="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydCaBN1ffHzaR5+DULmcfMZKikQaGBNFEaJBlKlIgQoiIhGTOEkFKSRmWIUuZ5TpLmNGow/9fnutv/us65w/Om+973ZPfuvWefffb+nHP22XutvdbKkkWbCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACKQxgaxpfH6dXgREQAREQAREQAREQAREQAREQAREQAQyDYGstp140smnkI4/8aST8h5//Am58xx3XM6cOXPlyJEzZzbbyLN37549O3/+6cf1a1YuO7B///5MA0gNFQEREAERyNQEpLDI1JdfjRcBERCB9Ecg/4WFi557/gUFsufIkePH77/b8eWm9Ws1QUt/10k1EgERSD0CbR/r3mfXrr/+HPvigKdT76w6U3ITOD9/wUI/fvftNwggk7tslScCIpD+CFSsVvPSx3o+O/i9t16fvPu/f/8tUqJ02QsKFipy7nkX5D/jrLPOQTERa62HPden+8iBT/eMNX9K5EOJMuClydP5++BdjeunxDlUpgiIgAiIgAhAQAoL3QciIAIiIALpgkD1S+tc3aF73wEXFileMrRCv/+685cp40YOQVC3Z8/u3emisqqECIiACKQSgSo1Lr18xJS3P6b/q1Uy3yl7dv/3XyqdWqdJRgLlK19cc8wbH8xftuiz+fc2qntJMhatokRABNIhgVy58+QZNPbVGdVq1b4yUvVMj/HPP3/v2mVd+7/08/v27d17wLaDltxx7OvduV3LTetWr0zLppYoU67ipHc/WfLnH7//dmnpC05Ly7ro3CIgAiIgAhmbQI6M3Ty1TgREQAREIBEI1Gt4S9Peg0ZNoK4/fLfjm7Urli5isla4WMnSBYsUK9GyfecetepcXa9VkxuuZpKUCG1SHUVABEQgOQjUtL6PcrZsWLdayorkIJo2ZVSvfUVdznzm2eeelzY10FlFQARSk8AzQ8dOccqKX3764fslCxfM3bBm5fKvt27ZZGPd7T//+MP3f/z2604UFKlZr2M5V4Wq1Wtx/Pc7tn99LOXoWBEQAREQARGIRkAKi2iEtF8EREAERCBFCZx93vkXdHv2hVGc5PneXR+dOGrIAJQV7qSY0/ceOHJ8qYsqVH5q8EsT2za7KSC80yYCIiACmYEA1me0c8nC+XMzQ3szahuLFC9VhrZtNIFlRm2j2iUCIvD/BIhHwbeDtt1Up2ppW2/za6LzKVO+UlXasGXj+jWJ3hbVXwREQAREIH0TyJa+q6faiYAIiIAIZHQC9z3YsStm869NeGnY+BGD+4cqK2j70s8XzLu70VW1dv7y0481L7/q2svrNrgxozNR+0RABEQAAsT0KVS0RCk+r16+5AtRSVwC+K6n9mtXLlucuK1QzUVABGIlMG3imBHk3bh21YqMoKygLaUuqliZv2ntmirWa6B8IiACIiACiUtACovEvXaquQiIgAgkPIFcuXLnvqpBw5tZfTZmyIC+fg364dsd2597snN79jdr+dCjCd9wNUAEREAEYiBQr9Gtd7hsuBGJ4RBlSYcETjjxpJPPPf+CAlRNCot0eIFUJRFIAQJlKlSuRrHLvvjskxQoPtWLPPmUU087P3/BQpx4/eoVS1O9AjqhCIiACIhApiIghUWmutxqrAiIgAikLwLFSpUphyAn6M/3m0i1+3Dmm1MJwF22YpWLz8uXv2D6aolqIwIiIALJSyCrbfUa3trUlfrt9q+2Ju8ZVFpqEShWqmw5zoVy3hQWS1LrvDqPCIhA2hFgvMrZly36bH7a1SL5zly8TLkKrh8zhcWy5CtZJYmACIiACIjA0QSksNBdIQIiIAIikGYELixSvCQn32mRB6NVYv++ffsWfjL7wwP79+8/8eRTTomWX/tFQAREIJEJVL/sirpuVf7fu/7685+//96VyO3JzHUvXrpsedq//asvN3MtMzMLtV0EMgOB7Dly5ChZplxF2rpi8eefZoQ2u/bQj1k39kdGaJPaIAIiIAIikH4JSGGRfq+NaiYCIiACGZ7ASWZfTiNdYMJoDX66a4c2jepUKbVBQUujodJ+ERCBBCfQpHnrdq4JP3y3I6IFWoI3NcNXv0TpQyuT161aLuuKDH+11UARyJKlaInSFzG2/W7H9m2xLMpJBGbFS18U6MfWrFi6KBHqqzqKgAiIgAgkNoEciV191V4EREAERCCRCewzswnqb16hYrKY+NOiFpISuc2quwiIgAhEI4D12cWXXH6Vy/f9jm++jnaM9qdfAsXLHBL0rV+1XH7f0+9lUs18CCz/5rBRUE7Lst/SAbKWz3eSmPkQKFuhSiB+xepliz7PKJBKli0fsBhZs3zxFxmlTWqHCIiACIhA+iUghUX6vTaqmQiIgAhkeALffbN9G408N98FBXLkyJlz3769ezN8o9XANCFgApfz7MQIW34yIcs/aVIJnVQEYiTQ7IGHHiXr7v/+/ZdVut9/u10KixjZpbdsdvnyFixUtDj1WqdAtent8qg+sRPg/VnU0nGWlltCcaHNh4ALuJ1RrBGwiHYBt1cvXyKFhe58ERABERCBFCcgl1ApjlgnEAERyIwEWI1mKY+lXJmx/bG22YL2BVab5syZK1fBIsVKxHqc8olArASCz2J2y1/GUllLJe033/FPMD/Pb7aQz7GeTvlE4JgJ5CtwYeH6DW+9g1gHn8+fM4sCnXL3mAtXAalOwNyolM+WPXt2Am5vWKNAtal+AXTC5CKQ1QoilbZ0enIVmlHLKVuhcsDCIqMoLMy6ohLt2bNn9+5N69aszKjXTe0SAREQARFIPwSksEg/10I1EQERyCAEgqbz9K9nWypv30/MIE1L9mb89MN33xK8j4IrVqtxabKfQAWKwCECKA55DhGysEo02naCZSC+Su5oGbVfBJKbwH0PduyKgHvy2OEv2OL84ykfP+jJfR6VlzoESgQD727bsmnD37t2/ZVcZz351NNO/99Z55wbrbystkXLo/2Zi4CNS3MnYUENin/uJca3eTMXsfhay7OJ4tm8nu5bv3rlsviOTp+5ywRdXKGs2Lt3z570WcuUqVVw8UrW0EUsIW7SUuakKlUEREAERCAw4NAmAiIgAiKQ/ASY1J1mqZClgMBJmzeBBbM/fJc9NS67sq4YiUAKESho5aKs+MnSWnMJFfC/Hb6FTEARzJDnYArVR8WKgCeBCwoWKlKv4S1Nsa6YOHLIgLPOPT8fGb/75uttQpaYBEqVrRBYmbx6RfK5Ubn0ymuvm7V003czP1u1tVqt2ld6kTnjzLPPGfnqzNmLtv6yu1GTu1skJj3VOrkJBC0MT7Zy4x2bMq7FDdR6S7uSu14ZqTxnXfHlpvVrceuXEdpWvsrFNWlHRrEYifOacO+fY8m5Fo3zcGUXAREQARFICgEpLJJCTceIgAiIQHQCeSwLgiZWdseyojt6iRk0x8fvzXiDplWpeWmdEyz6dgZtppqVBgRCrJ2IDPqrpXWWosWvcG4vsK7QOCkNrltmPmXrR5/o7awr/vj9t18ROsPj+293bM/MXBK57aUuqlCZ+ien3/d2j/d8BleKuXLlzv2QffbiM2DUK29Urn5JbeJDVa5eq3YiM1Tdk5UA7zWUFSdEco/ocUbeo8QZ+58lWe1EuCQZLX5FNtucEmbtyqWLk/VuTIzCiPta0tJFlrCe1yYCIiACIpAKBDQRTwXIOoUIiECmJMAK7S2W8POaqUyn473aKxYvXIBrKAQvV1x7faN4j1d+EYhCAMUDQt/zLRWxxLMZacPVBYIZnls9u7q9Uo0AroOurH9jY9wGYV1BsO3jTzjhRHyG//rLTz8mpSIogc865zzufW1pQIDrd8GFhQlUnGVNMgaqPTffBQVcc378/ttvwpvGveOEpuxbsnDB3DRovk6ZPgkgfGVxCG4S41E88G7EVSJBt+M5Ln1SSMFalSlfuSrFr125LEMI9wsXL1XmeHuZ0KZ1K5cvSUF06bVoLG6d1a1chabXq6R6iYAIZDgCUlhkuEuqBomACKQTApiAs6KbzdP9TDqpZ5pX44Bt77459RUq0uDmJneleYVUgYxGgEk2igpWxbEyFJcWkTYXu4J8gWfXXEhlNCZqTzokwKp54g288tKQ57GuOO2MM86kmqar+J6AzfFWmRX4r7wzb/Goqe/MifdY5U8eAsVLl6vA6mTzCvPP5g1rVydPqab8CApCt2xct6ZXxwePcve0Z/d//21ev2YV5/ti/pyP3pwyfnRynVvlJDwBlPa831A6xNOv/GH5f7D0u3s3JjyJFGgAfbizqsoo7pMuqli1Oqj+/eefv7d9uWlDCmBL70XyrGA5j0soKSzS+9VS/URABDIMASksMsylVENEQATSGQFWotWxdLklAvhqi0BgxtRXxrG7QpXqtQoXK1lasEQgmQgwyeT5w9JpjaVvLXkqLILuo1x+3GUwOdUmAqlCoPplV9StUvOyOjtNO/Hy8EH9OOkpp55+Bn93/pw064rLrq53PTExfvn5R4SM2tKAgBNcrlu9fCkBeJOrCj0fbdP8mW6PPtjs+joXc8+El4uC647r6lS7/dpLKrW6o2Hd5Dx3crVB5aQZASwHcY2Iy9JYLSVQcpSyVM9Sfku4htLmQSB/oSLFzLDtFIT7KBQzAqRylavVoB0b165awSKjjNCmJLThLzuGRQRnJeFYHSICIiACIpAEAlJYJAGaDhEBERCBGAigsGAVDpYWf8eQP1Nn+WrLxvXLzTUUEG5pdl/rTA1DjU8WAiEKiGJW4CWWUFRsNGuJSCtKEcrgPopjNClNliuhQqIRYAU+1hXkG/5cn+7//P13IKDtiSefcgp/f/3lZ4LFx70RmJmDVi1dtDDug3VAshA4vNI6Gd1BUbGvt27ZNGXsiBfcveJVWYL9rl+9YumB/fujWZUlS1tVSMIQOM1qekGctUVmUM0S7uW4nyRD8AFYtnxlOGVZt2rZkozy7F1U6ZCFxcZ1q1bEed9klOwo9lA4M0bEpZo2ERABERCBVCCgwUYqQNYpREAEMiUBFBasQGMFm/raGG6B1yeMHk62axve2hS/3zEcoiwiEI0Azx/KhwKWWFX6S5QD8OudzxJKi2jBuaOdW/tFICYCDW66vVmREqXLfrV54/o3Jr/8kjvoRFumy+ddf/6BC5a4NydkksIibnTJdkCpchUDAbdXLVv8ebIVqoJE4NgIML5iQc0OU+DHo8xi8c1cS2stJZu10LE1Jf0dXaZ8pUD8ipVLvvgs/dUu/hqdcebZ55yXL39BjtyyYV2yubWLvyZpegQWt1jorrOksWGaXgqdXAREIDMRkIY4M11ttVUERCA1CRCUEHceDHIROsklRxT6s2ZOf61Dt74DTjvjf2fWb3T7na++PPLF1LxgOleGJMBzuMnSuZZwDRXNXzfxK760hOk/SZsIpCgBi42ct9WjXXtxkkF9uz0WuiL3uOOPD7gT3LXrzz/jrUReO9YJmdatypRBUuNFluz5Tznt9DPcNVi7YumiZD+BChSBOAmY5aFzAYUVVy6+R7E6dGfg3fmfJVx2breUGeMYxES7VLlKVcjoXPKZZ6hde3bv3m0e4fYeNHdKofGIiHeR1SzssmfPlj1Hjpw5F3/2yZz3pr82KaYTWaYKVWtcUrx02fKTRg8bFH4Mbqns36nff7djezyWHryTstv2965dgTGQU3zzeVMwLk4s9Tv9f2edXbFajUuoA+3CKiyW49JpHsaSuET7xpKUden0IqlaIiACGY+AFBYZ75qqRSIgAumDAJM7VrExQE+SO4/00YzUq8XevXv2vGmri+9t+8jjNzdr3io5FBY2A8zBpO1PC2CbUf3uXlikeMmSF5WvxLz3k4/en/nHb7/uTL2rlu7PdLrVsLAl3F/8aimSwgJBDv6JmZgSXHR3um+dKpjwBO68/6FHzjz73POWLJw/d96s994ObRBBs/m+Z8+euO/FAoWKFqdPwJ3UD9/tQMgS85avwIWFb2p6z/1jhjzXl+Df4QdSbuHipcqYPOrcrZs3rPvh2x0IMI/ayFe2YpWLTz/jzLMWfTpv9q6//uS5invLbRK03Llz5zFDk99iPbhG7SuvqX11/RtOOfW003/47ttvZk6bPH7DmpXLox1/30OPPXH1dQ1v6dz6ntvCg2Sffd75F9CWH00C+MtPP3wfrazS5SoGBJfkjfcaRCvbb/9xefMev3//gf0E3Y61jHPOz5f/+pub3j1h5JABf9tFCj0uV+48eVhgbWFQvsPFVLQyuVZValxy+VnnnHf+VrMYWvbFp59EO0b7U5UA7zksgHF5iED6uzjOzvuURTgcg8WitjAC3P9FS5Qqy8+MzUjxQDrN+pdYFRaMbwePm/r28SeceNLs995+w/UxPM+P9ew3uFaduvVxN2iP7T9D+/fuNmHkC8/51SX/hYWLNr2vTfvL6za4kUVD5Fttbuy6PNi8ablKh+JXMIbesmFtVAsLlOUPd+nd78bbmjWnjhxrupq9He5r0pAxajw80lFeXEEVscRYUi4W09GFUVVEQAQyNgEpLDL29VXrREAE0oYAE0JMhp1VRcyCg7Spbvo56+uvjBlxd6uHH2OSV7n6JbVZlRVv7RCS1b/ptjsbN723pbnjqMKEDUHX5DHDBo8c+EzPSIoLVoSNmDLjo99/3flLmzsbXctEz52f1W8t23fuccOtd9xjK+X2jRv6/DNTxo0cEql+1OX50ZOnIzxksvblpvW4Uji8XXvjzU1atOvUjQniBzOmvfpst44PoriJpc2s3O327AujCNTr8u80qVLTBrWr+gkQYyk3g+VhgonPbVxBESgyWoBRJqNFLSHgDayIttWnGQyJmpNeCPzvrHPOveuBdh3pk57r+Xj78HrR5/BbLAGTmzRv1a71o916Ixj61wIb0PdwLAL7uau2HXaFZuEM9qPUHNS3e6d5s96d4cXiiWcGj6T/NXflSz+Y8fqU0Dx1rr2+UbsuvZ49/4ICF/I7K3f79XisXXhfeM0NjW+nbytgAWjJR5/U7IYrqpv2BLcaUTcE73e0eLBDA+vLz89fsBAH7Ni+bevAp57o+PG7b03zK4B2d+//4mgE8KF5br/3gYfoswc/3aNzpJO3fLhTd1vunL1ardpXOoUFfezDXXr1K176ovLu2DkfzJyOMI/Aun7lOYXFGg/rCuKL3Hr3/W0KFi5aAjYmUHwCpU5UMD4ZWGnduuMTvZ1w8bUJLw17uusjbWIpr0ufgcNQ8Hzz9VdfvjNtygSOQfDa9rHufRo1ubsFK65ZFf7uG69O7PnYgy28lCFwv+WuFm1aP/pEL5OfBlyZsaH0euGZJx+PpR7KkyoEcFF6niVcH0ZVuoXUCGU/ygqOZYwSCLpNrCi9I/+fUokyF1VASE8/N2rQs73sY06+05fbv5z8zZ6DXw595388W2aEsYv+Lby/jXRH4KgJZQV56PP5W7RkmYtGTJ7xEdZd7lie35btH+/hp7Cwfqjtw11798uVK3duFJabzYoCBQaurV54+fV3XNnbvty0IVLMHM5nxhSnDbfz01fy3lptrvDOs3cFY9yHuz7Vf/7HH7wTamGSKnd88pyEeRzPC/FfMmvQ8eQhqVJEQAREQAREQAREQATSjgAm9pZqWnrE0q2WDk/e065WiXPmweNem2nMDvYfOdFXKOXXGiZLo6a+M4fjXVq2/Y8D7jMKh0gkEGq5vKFm8AiwBo6Z8lZouXwOVRZ4lcvk0R2D5UhonmYtH3o0vDznGiba1WJSPG/N9l85fsH6b/8Y+8aHCz7f/OM/fEfYGO34jL4fIYqlbJYqW3rOUh9LN4W4wzgKge3Lbqm+pQ6WKlnKGQzcndFxqX1pRKDngOHjIj2ztzRr0Zr97Z94qn+0Ko6Y8vbH5F3y1a976RO+2PLTv+H9i/u++Kude66+7qZb/crkePJWv7TO1aF5Huz85NNeZVIeVhnkxf2H68Ppe9/7fN3Xrg9+vM+AodHawf5ipcqWe3fh2m1effjSr3/fX6XGpZf7lYOiwh034e05X/QeOHL8B4s37HC/oXDxOxYhvctX/bIr6pLvjhZtO7j6c+5ZSzd95/KguInUHoR95A3t+xFUUqdwjlyvCwoWQsEa14aioNUjXXqGvudc2YWLlcR9T9SNa8Qxda65riGZsUqcOHPuIq9rXaJMuYrhBbIo4MkBw8a6/FNnLVw1fd6yje5+ZMV31EooQ6oQsGvCPd7I0p2WDivgop2cd6elxpboAzpbOoP3o96RR5Jrel/rh7nvWUwSjemx7q/X6NY7OBfPGmUVLFysBMppfpv52eqtWEugdLi7dftOfmNV3LCSf9HWX3ajuHBKcpTpM+av2BzaB/CMR6ozx457c9anHEP/XcSs8MiPssKNT53y+VjbntrHW5uOt8R48mJLBXTvp/YV0PlEQAQyKwFZWGTWK692i4AIpDSB/9kJWFnKijT8kCfJFUZKVzI9lo9bqFp1rq5X+6p61+NW4sfvv90RSz1RVoye9v4nhcweH8uIkQOf7vnGpHGj8MPLJPKhx3s+06xlu0dZZeZ884aXi/sSfsPKgVVmbv8DHR5/khWxrF7GTJ5VrAiKrmvc5K5FC+Z+7Fc/Vx77161ctsTlu/iSy6+iPnxn9S0TTQKNU97Qfr2fiNRe3JIMe+WtDxEMfj5/zqxOre++jRXTl155TYOBY16dwUrZWHhlgjysTseVAXEpWBG6IoqvbtxksCqRIKS44GEVXQ6bmDJWwh0AQUr5zO+4RsGPMd/5y6pVVrRzTlaisvqUctjP786lD9/J6/K4lXrk4TfflXtaxZqx7lhW32MJhpukIc/27OLVOmcN5lxDRSLQ9s6brkUwxMpejkOBgWC/k7k2wi0PFgsIlPbbsldcFPn1gfS5btXub+ZPyp0TBSvWb3x/feKYEVgElLqoQmWE8pR7VYOGN8+Y+sq4YZOmf0gf/OmcWe9heYHfcgRd9G24kYp2FeFiK3RnUUKTsHkAACAASURBVAdzvb4NiwrciLAk+cnnho5B4dDS+mM/awSUzpzj3TenvoIFBJ/pK4e+Mv0D6lvQrN386lC0ZOmL2Ef/v/jTT2ZjXeCURQs/mf1hn87tHmAVNEoMfseKhPp5lcf7oUyFytXY5ywsUHz3Hznhdd4lnIP30/avvtzM6meUBHeYS5anHn/4gWiM3H7Ke7L/0DHcR/zGu3LG1Ilja15etx5K7XJVLq7Jb3aL+QZtP/vc8/PxTuF4AoOzGhv+JcuWr4T1yND+vczy45PZF1WsWv2AmdOsX71iaXj9UGRxfbG86PbwA3d98Pa0V1FijJ8x+3OYV61Z+4rpU8aPjqVdQQE44yb6w8Ou0NT/xUIvpjxwZXzKu4Y4Fp5bmCKCdxbvP1bxo1Tj/YbVE+/MPy0vrut43zHWxRUqZWOd6hL73fuSdyx1YB/Xl++4euNYymPjPco7d5sljuV+oK78zjuUz9zTnNPlpU6c171fOYdzAXkwte4fZ1V1LNZSQQZR/1xc6/IryfTZ3I/exw3TgFGvvHGyWdRhmfxIi6aNnAs9xqxehWGVx9gYK7l299x6PeW4fD+b3zus8PqPmPC6+y1aEPE2j3V7ioU+v+385efmja+5jP6bY3FL+N0327cVLFKsxJmmCNlhllxRG5f+MvDMXGsJl6vvpL/qqUYiIAIikDEJSGGRMa+rWiUCIpD2BJiAMbkrYCng1kNbbAQwGUcAz8Tr6usa3Tp+xOCoq4sxsMciA0EZE60Hbr/hqlD3Sy8PH9SPiRkun6rUuKwO7jy8alOqbIVK/I6wypm+o3S4p3WHzgiY2jZrXO+L+XM+6vr0oBEIs4qVKlMuUqtKmdCH/QgllyxcMJfPCKZ6Pj98HAKtYc/16Y5ipe71N93Wd8iYSQgLabdfHAqEQM8OfflV8qxY/PmnDzZrXN+5kHKT0v+Zw/HYSGf4XMdbC1nZ+5UlfOx7+tkPoYDfZvx64yoDtzX4965vCZ4IVRDU4OaNfLjYYQJbwdLnlvD7jkCG7+stca23WbrOUmVLuAJbaYlxF+6mOA/Cmh8tbbGEFRb5cDlAzBv2UQcUGShHdptQCIEMv+OawCk2DsfkSC2BjJ1b2zES4NnvaD7GD/UBT3VHwONVJAJifnfBtyOd1sJc7HY+zCnXBMWBvmfl0s8/o0+MtcomzyewaGD7befOQL3oAx/s1KMvn0cNeqbX0P5PdeMz7j5cXvPiV+bFiW+8Tx+MAgZXQM71h3NpFc21Ff0flmwoK5Z+vmBe++a33+iEbnbj//uiKXNRWCA8R0EdHl8DoV2REqUD/uPfeWPKRFc3ynj43ttuwPrijcnjfFc+Fy91yOXTlxvXr72waPGSj/Xq9wLfZ74+eXz3Dg/c7RRIVvYEFBbEHkHR7KX8wVqCOsLAAm4vphwsMlBWUJ+2zW6qt2rpooAvdOcarIIFqI31OnGNsdCp1/CWgFIGv/dPdX6oJXXBtRP7uvR5fhhKkOsvKY+bO88N11fsQEHPfdJ70KgJKCtwU/XgXY3rO7dYm9atpv86aqt5+VXXosyCTccHmt3s4rDwfd2qZUtQWNC+WNtl+egjea/SdyPUZsHCVuv/6I9DhdBHFKn+L2bC8KU/4F3Fu26zz5G8e3iHFrDEu4/jUPZhtXOKJVxD1bTE+wnlgRt3cM2IA+XeXSiqGAPzDg23bhphv3H/oqjwctfIGBqFBe++Ny2h1ChoCaEx70fuDZRtvItxH4obx1rBen5mf3m3slgBay3eq06pwbsaJUayu/YpXb5yVSs7y9LPP53H35TcKlusGMpfMPuDd9s/0ee5AoWLFl+26LP5jFOjxZvBIs716SPNdVWossLVeb4pinmOGXfyG2NOv/ZgTUxfw34UxU5Z4fK7dxgByFOSSQqWzf3PvcY9qDldCoJW0SIgAiIQSkAKC90PIiACIpD8BJh4IVRkgsbAFtc0rE4jMVFCCMXEm79MmJzQ0U3YPAMDJ+KEHJcmBYsULfHME4+2jdVvLVYMs96Z/jpBX1m1G4vC4p5W7TtVurjWZSgZwpUVXF7ObTKczSgsEKh5KSxQJDhzdbcfn749+r04mgnbgF7dHkNZQXlrVy5bjMIC//CRbh/nPuPTOR++5xQLHbr3HXCGKRXmfvjOWygrXHmuHMr0U1jcfGfzVqzaRVD3yP133BQa78IWUDORymLGJb4+1ZP/Vk/XJSJIIeg9PPwEIqENINYFyginnODZRFCDlQYrr/3GTAHXMSEbQp0bw35DiHpb8Lf59hehSui2zb4U8KCJYgThEArQMZbWWCJwML8jJMJ6hDr/ZX0Mygz8WdP3oAgJCGUsudgdAeFMFCsTjyokz08+rkPo81xyfKkzq2uddQrfETqxypbfEDqF9qNcWwRrLvYLzwFCM/pbykHQyb0Q3q+SH0GM64OdMDTF+18E57jqQKn66sujXvQjbDrSQJtMJh5XIBVi5iD03/nLTz/GG8+G/pFzIvD6yQTYWE/gZo7V/B+/N+MNp6wgz0nWWbm6X9Wg0S0I0bE4QEEc2ibnLsoMOyLGrzALirH00QjJH7r75gbhioCvv9qyib6c/pjVuuECNBS5LnbHf2GxJRDGv/RCv6ci3c0lyx5yd7Rp/ZqV1AXLFqzYuj/S6p7Q2EcomFiVDJPj8p5wgpfCwllXfP3l5o0orLF8Q6CHFQLxkUKVPaw+5rzxCPaJL+GUFbwjn+/d9VHXtlPN1MZ99rOkcfsrB91rLZj94bsozimT+6bFrfXrfLNtKwJf3w1rDOJfkGHsiwOeDg8an9fYsO/ff3bFI6TkeUS4zEp9rgcJRTECafo9lLv85Zkmb+gYKlJ1j2lflP7Lle36Dmdxh7CdPoj+in6L/gthPmM/9pGPfSRnPcBn2uaEohxHPhL9AeXR37l8rr+Eg8vrmByO2xQinOedgXKB8iKNX9hPn4uyifxcQ44lcX8FAjMH20Ob3OasJNy+SHFU7g85zusj7WSDRZMoeVG8zbLEMdUt3WKJRQqMAd6whHIV5lh58X7AVehc+8u9RFthd1TfH8+4m7gRxBbDCiseJXGUdnnupk9FYYo1MX1iw9vvug/rOiwroikrKBBXULly58nD+2GsxfbxOglKcGJaMDZmTPrVlo0sxvDc2nft3Z/+8O3XJr2MNVpoJvplLLnoM7/eupnrcdQWfL4YC3Avcd9xPfjOPewsXn3f0fFcpwjnZ5ezdg3PxhgMBRmW0hpjJ+Wm1TEiIAIikAQCUlgkAZoOEQEREIEYCDAxwg0UE3YEZwy6MaFH+MmAl30MyFlpzV8m6CWD+VitzQCd31lJFnA1YwN6BJHsY7LLBItzMIFlEO9c07h9bvIVWBkVzOOq7SbTfGfyy+bM9amrc1fDJNGZ+jPBo2wnBI0aaBGXRwSURbjzbPfHHjpokxVXgWh/P3r3rYDCwq3OjDT5YyXrfe06Btwo4YIkPLC1O5fJTBBcZmHy5HX+0ICqCG/Ic+f9Dz6CYGz54oULJo0eNsgdd9CkV3wmgK1fWxB2FSp2SPg3P1heucrVaiCsZIVtLwteGl5epDJZyduyQ5cnyTOg5+MdCLAdem78vvN966YN66LxzST7uc6sxuR+Z6W4exaOar49W+xDEMNElGvr3Exstc8Ia5zQJjnQFfAoxE8g7QJnIiDCHQ/9BnnDV6Nyb0+2hAsalCOTLKHY4Ll1yg3aUsHaiiCQewThMX0KfYVzecWknOffle+Uq+FCfadkCO1fQhUjlOH6D8qmzgi8OA5BF6zZcA1Bn4L7PNwtsI8+D+UR3LnH6fMQcqAIoq64raCe9KUIx7hmWKdQDkIpgkFzbo5x1/JX+8zqUPpLVsByb9B+BCOc7+tgOex3K3qdyxL7Kfk23BPhQocSUeRGsjrYvXs318e3z/KrFcoQ9q3xcQUSqTWFih+Ke2C6lFUImG5rfn9bYiHgRqrno22ahx5rsrlAMGw2FAUzXntlXLiygn1OEbx1s3/fhFujqrVqX4GQrLO5sfIStFMfk/f/i6D8ZJMOhrcjVNH7PxPmxXvVnIK5uJnGsWL4WzNV6Njyzps5b3hZWYOrjr0CUJO3bIg7KIJQ97BA4Pzet0uH1qHKCn7LYZF3+WvCwcA7KtqGUgG/9OQj2HmosoLf6l7f2ClHzV3MrMNuXrzKrVitxqX8joUefvdpa8eWzW6OpqzgmKbN2zyMOyncfo14/unAuyl0Kxq0QIzzneQElPQtCO7pE+g/YEQ/XsASfQmLB7gHGDudGhR40l/AkDLc2Ig+x41zuI58dsJ9pxR1K+9dXsZB9C3kpX/g3PRJ7Mc6wQlV2U9fh+IO6xj6Diz6nBtAFN4I0qkTK/7rWCphiT6YvodxHn0g/RPKIVxScr7XLBEThr4cxTR9lYtHQl3pK7HO4Z7iGeQ94ZQh9Ie4qaTvoJ9EgI///WX2l42+9ipLtOk3+53nxClIKJvj9pgAeJ/to168K9z4FasM13cHizv852371CD8R/vumHvsyrLCfoxopep1kP1GG50yIzQLrJ1yjDbBHOtG3gm8L5wLKq4b70NY8xv7V1uivdx3XGOOj2tz7qBWRrBEiKvACJkZS7J77cqlix/p8fTz9L9PPtL6Xj9rvdCiGFfjQpTfXjSXb359GAt2nHtAxsB+i45437i+G1eB4dWub7E2+A3rD9zMxcCA54P7k2cEBSXPD88k15zPPF+MC3jeeD64V91chfK5j+kz3H7KCSwes+QWr9BX8I5nbOeeY87BuTmectxndyz3MotXuHe+S6vFHzHwUxYREAERyDAEpLDIMJdSDREBEUhnBJhEs5K6iiU3kWQChEkxAgLcK+CygwksSg0Gz2d7tAEBJZNFJrMIIN2qYX5n0M5gnUF1AUtzLTGgphwm9p9YQpDHZIzBN78xyGfAzwCeQH0M1HEXwXFuRRMTcOcfmEk/k2WOd+8M8kXcEKagrPj9152/PNDkhqu8BD6RCliycP5cVqUi6KlcvVZt/JH75X/AhPgoB/AT/tarE1iF7rk55YJ5j/J89zn3TghqcK3Cue9s+eAjCBSf6tSuZehk7dTTD61gjeQbHGWFC2CIiynyt3qkay/+vvB0j8749XUVdeVFKvPmO+9rhYuRLRvXrZk5bfL48EY6P+afhvgh9gJhEzsnlDlCCJdRJl8hK/VYSVnAEsJ7hEKR7lvuee5xBBabLc2wxGo6JrgfWGLyyz4mwAhsEPrwbPFsMuFFOE5ehFYczzONsmqcpbmWWPHJfgRbWD/wHPNMo7C8yRLPIv0C5UbamLx7bfQBocffbt9JkTYENTz/9AsI/mjbq5aoOwKbAsF9CPNpH6tVEWZxLo6lb0M4hNAH9y30aQif4IYLHAL44u6D/oiyUZzQ9wRc9gQ35/IFoSSWJNyTlIPbLMpyK8Vfss/0l/RbCOdgifCMZxk3IFw/2kAZ1BdBIfWgfQganYKX+nINyMfzR70497ZgXtpGmfSvHOMUwfYxeTaUFTzvuPDB13ikUv/79++AcIeVu/GcHT/i5I/mc9yrTGdhsXHNyuW4WLq3zSOPk++Zbh0fdO6Z3HHESHCfUUb0ebx9q/AysZhgdS2/+7kUof9u1aFrT/JMHjN8sJ/Smf2R+nEs7LZt2bQB1yjljMEHM16fEis36oAbKPKjrKC/797+gbu9+njigRy25LAVzl7nKF3ukGsYFAHEqMCqbtbMN1+b7vGOOue8fIwLsvz43bfc9xE32tal76DhZJo3690Z/bp3DMTscBsunohf4b5/sWBuwCrQayMYNm64WKVd++r6N3Cf4cqLmCfR6gED3CyS78V+vbqGWvvxGwp0gu5yTVYs8Xcl43Mexhy4x0PgTD9KYixCn8lYCcVsPUs8HzzjV1iin2GcgOKS/fStrl+nj+ZZp1z6N/oxjmVMRp9EH3aZJfoNxj4I+tmHkgD3kfR3cKZOzvUReXgXhP5mX323Gzz2oPhwQcwRtruNcWG0DeUG5/eKyXKvx8H0fQGLF9t4F9ImxoOMB7Dc471E/0oiLsUmGxPAiID1MEdBAiv6SPpMXHViuUA/yRhzmyUsJngHko/rwTm4l+DLu4189L1cM5QVKEPoj+nf4E1fzX7OyzmddR3Xi+9cU9415KVP4dyhgmnqRv9P+dwrPFdw4hzkox6UST4UR5RF29lQ3LCPvp+YD8Rq8bS2C+Y/6o9TWCThfvcr0vd3lA7sxAUeSvAP335j6mfzPmasEnXDhRuZ6GfffePVw67zwg8sUqJUWecOatnn/n3CrXe3bMuxjNOdW0JXFpYgLdp16sZ34sdFqRy8udaMSbgPuV9RUnCf837neaGPZJzAs0l/zXiBdzlWqyjvuI+5/ixWYfyAcoH7kH6BMSH3GPePG+dxT3LPMrbifuRcPIsc4ywIeU64rxjDcK/SB4y252K9PSNxK7bsWG0iIAIiIAIxEpDCIkZQyiYCIiACcRJgssZEkgEvE2UG4QzGWcXlzP+vDykTASaTqfBVowyimRgzOSExiCav2xgsM0DnPAzSmZBzPnxxMxFlYM1EjEE/x1EWglcmBAzUEeox6Ccvk0Qm3y4AIoN0JrnUnTq7lYkhpz/6IwGlcVeBoKJV0xuu3rh2FRPTuDaUBAjzEKJUrFbzUj+FBeb35jYK0/8s+E2P5HYK4Rv5/vrzd88ApM5/Ob7Tydekeet2mMK/+vLIF8MFaAh6yBPJxQmrdMlDgEFM9WlH5eqX1MZXOMFWQ4Gcc/4FgfIw5f/LrC/CYTFpRGHB7+OGDXw21D0Jv9W55rqGl1mQcphPe2XsSD/YQWUFwgYmdqwEZeUYk7qTbB/3DtcZARxCA+4jJoLufkXI4YRzCI+YNB5e6X+s/qCDigYEEAHrlWDZbiW/M9PnGSKPswLgs6sDn52bH+eigueHex+muIDgHg6UZfUNVdjAgecLLnMt8RwE/PdbPp6vLCEuQTgPK/mZ6PPZPRfOqgBenIN9zhUI+d1qXtdGp0AZa/uc9RKTZZ5XJsZw4L6gH+EacS2utoQAhs+0CRcNCKe4t2kzzzMTchQOCOkiba4fcQI48gaeJZ+NNnBfeAnIopwqsBshUfjGakcUpihsnCALdrSB+xEuMEHYhGAJgQOCKphzXeizsIZiFS2suAYcw33KPoQW9F9u5SzHIUALrC62BDOuEQI2fkNY5WKEUJa7F+3jsW8oEnDdgTL2ObOSilaiLbinD85y+hlnIqiLeStf+ZAiIZLPca/CEMJfaMEo2GdekZbdfk+rh1CuEED2I3PTF35MleqXXu5+Q1nh5YqkStDPOpYTfsFf695w0230qay+RWDu11Dqh6Cc/X7K4nkfvfc2Qv3Lr2nQEIu78L7Sr+zCFoMjNLg5ym/3Lgg/5iyrrKsD7Qrfn9tMQMyzVkAxx/vm1rtatMH6o2/XDq29zu/ibmzbupnnwHcjVtPTQ8ZMhgE+4rs8eN8d4e1r8fAh4SAb71ECafsVWOqiigGhJ24YUXh/v+Obr/FnH8uNhhUH1ooo+MPvDdrfpe/AgFJl2itjRrh4ULGUG5KHZ4/nkvpjlcqzSx/C2MpZfNEX0WfzG30kSlqefxQ2zjWRE7JTNEpQ3v/sC3VdFFo112/SP9MntLS0LZghtK90lgb8FsmKIM5mx5U9nr7YKSs4Ae0iYanB84QQFuUewmDGBwFL25B3Hn0kbWSMSh8JUwT69NH0kyiz6be5LliHuI19TujPghuEy6Eb+Rljcl6O3xB27OHxRbAcxiwkNpQK4fvdOMHVBaE04znayvuXtjqlN/cL33lncq15t/AsO2VWWFWjfy0TjF+RFEVx9NKPzFHM/NfxC8oKnnPGv7GUgUUU40XyvjVlwphI/WOo1fFSHyUmC3uuuPa6RpQ39eVRQ0PrQJ8+csrMj6njO9OmTPjEYmLEUEfuCd7fJJ5V3t28/xmPMZ5zn5krMd67zBL3Ju9ztyChgH12CxUoj7ED41l+owwUoTy3vIO5Pxg/cJ9iPYFlkxsXuOeac3J/MN5iXMF+xvf7g0oL6qFNBERABEQgBQhIYZECUFWkCIiACBgBBrhMfJn8nWhCzz2sWLPPTPBmWWJixAQOAQaTwbcsIZzCVJ+BMINnBt8Ij3D1wqQZQedcSygnEPKxn2OYLCLQYvLK+fAf+6klViVyPvaz0oxJPRNOVpsz6eMY9rECicE8G5MCt7oQZQj1DAh2wwS8wexH/mHy8uSAYWMRLPV6rG2L9atXOjcEnvkj/bh80cIFKCxwR+KXjzgSCPOxOnDxJfzyulWs4YFaXX7nvgKhGgKh2+994CHckni5ushXoBCTmiz4J/c7n3PR5IR097Y9tFIZH+/hk0Tn4327xdnwmkBWrXnZFUw0EXrNevvNqaHnrH5pnav7DBmNFUEWVtviuiUKbCZXXFvGAAh9EUCwWp57CiEM954zm8dKiPsN9wEIixAAcM8x4UNQhJAYYRICfcpD8MDkn0khEzvuN6ckQAhC+dxr3PPs4xlBmOBcUrDCFWG9c92AUo1y+J0VbhyDwAGBIccimKc86lLAEvc135lQIlRBoMpEEz/aCCZY9cz9/YvVl7ZTX87NMawApa2s5DxKCBniI9kJsY+wULFj2AIufHw2r/xkDayiDwqHeP4CipLgRvsQ2DnFDH0BHOFHnWE+0BLPN3yoG8zoG2oHE4oVBNjkRdHRNVj2guDvfOWczpoB6wgm807Zw7nZWLV8LBv1QzAAdwRK3FMwoV9EuEnf5YQO7to6ns59B23mfuU47gPKQbBBHSnHKRnYz2fuXzZ4OcEZ1/eILTmti6698eYmhW1l+W9mQYVFAoJ1FBQWa3RX92eHvBRwnTT1lXFYS+HmDWGTbXtNZrz377//+ovV7q5yWKjxmZXvWGshWA6ve/h38iKwR5BOrJ1o+UP308c4xe761cuXDhn/xnsogU25EgimGrpZmIQzXZwGLAf8hPtVal4WWC2OGyQ/1yONm97L+y3LjNcmjgu34gg9Jz7b3Ypfv358+pTxo1lBTN5LrrimAbGCYmEQKpzjGoTG6gg//vz8BXjGTGH9He/Xo7aSZcpVRLmAAocg4Xwe2KfbY37uWoqWKI2gLMsWi90Rqa5YLfJewWLx8bb3NsG/fGh+rCucsipQnr0XI/mzd1aFvLfJP3xAnx6x+L8n7w233HEPf1+bMHp46EIB/OIPeGnSm7iJ+WrzxvWUGQt/l8fHFz0uX3iG6Zd5B/Cs058xzmLcQ99N/0E76McQcvI7/QVjEN4XvN9wj8V7gfddqKWXVxV5L7kNQSXvOvon3oG8R3jXzLFUwBKWBliAsVKb/pj3Jy57ENDS33A+LF3ou6kL/TX9EUpaFAks6qBdfOY961zQULYTqiPsp1/mfeaULjCgb6S/Q/lE++kz4eFWg/NuZIMZfTDWV86dklPUUh59KbyoO2MILyEsbacetIF7L6CQCF4z179GUvL67QtVbASrG/jjynS/xfrd5YMLyb3P3WIVxsC8c92CCN4fqyzBkz6WtoefK7Renp9LlatYhTFjJAuxqIXEkIF3iFNykh1rvVhcuJGXMTWxJuhDIlkuk7dk2fLc0+aqbtdfG9auYr5y1Fbz8quu5ZnHLdz61StQYgU24uF0fmrAiygrCOjdw9xVRWqaz3PvFFq77FoxFnL3KGNKxm08/4wpeS65t+mXee54DlwcL8ZCH1vimeLZ4DjmPXzGksItlHDzKZ7rCZacEpT5B88tYySOoY2MK6gP7+q475NIHLRPBERABETgSAJSWOiOEAEREIGUIcDgmcknE6WfghMjp4RwPnZxNfCOJQRvbmLFBJfvTM6dSTSTLEypGZgzkXJCYAbzHMekE+UDk1n2M1lnMjnXEquQqAMDejdxYx+TMt4B+CpmJZ1bqXZMg+/GdzZ/gMCh+Kp9/63XEa4meXOTH4RvfoVcY8JB9k0ZO+KFSCdixee5519QgDxMrMLzsrK2YPA8KBiIM8FEa9hzfbp7CZkspi3KoCxbIwQhLFrykBBq9fLFX6B0wfIEqxEvs33nhsWvPIRelGWxPaa5Fb3U+f6HO3W/u9XDjzEBHdqv9xNe7kZC2xq81txP3J8I9RGOcK8xWWeyx73BvcLkDqHMZZaYpHEvIlhHmIFAiPuEiRxuFfiNe/B6SwjwtlnCzQX3I/c3k0qOQeDjrH0QGASEsbYhPEEBxOQPQUuooIgVlygREEYhRGGlHPVjoulWuFIGdePex/qADQETdWOjHlwL7n8EE0w++c0JbRAocW5cSFAuv7tnNFhEyv+JEDQS1k7Z4YR2VMgJtuG4LWQ1LIoZNgRLgy3RTyC0hSvP+RhLbgUhwiz6KZQACPDgwspVOHF9ETZz7REQuNWplIuVAtYL9C+cHyUr9wHKFc7BPUYZsEUggLADJSr3EvXgnnjaEvcN14381NOtkLWPR1jaOKEYv7stoOiJskUV8EcrIJ79CJOfGvySr4sNVxbKUJJX2SgwzFDqL5Qce/77L6CwQUDVqXf/IQQ9RQkcyWVPuUrVapB/3crlS7xW/0dqj1MO0+fh0gilxAdvT3t107rV4Sujs1xuq3Sd8mDMiwM8rSLoly678trrOOe8D9+d4XVu4ls4xQfuoCLVz/rowDONUvebbV/yvB61bTMlMn0silxc+sWusDhkEcf25uSXX4oUNwmFFPkQyHvVwbWHGCSX121wYyR3hVjPwJlyIin47fV1YYuHDsVqGjHwmZ7hq7i55q07dusdWh8/IaPLU9R8R7nPxOuY+cYUBHVRN97xtBFFxQczprEyP7DhiqrXwJHjeZ9hrYE7yCRaV0SqA/0hfQaJPpA+hv7IWbsxruHdQHLvEvbxHqG/QZg5zRLPFkoM+j+U7gUs0YfRf1I24wTy0v8xpmJz4yP6T5S/9EG8Tyjr5eBn6kR/yWpz+msSi1T4y+Ys7FxZfHfuOF3/nMS0DwAAIABJREFUx/FOiO/m6k7Y7xTIfHeWJpRLWzmGMqizWxhAXV35tId37H2WuHdxIUSfHRhLBuNWfB0cJwSre8QfzkF7qR/cjmm86HWC1PwtqKh2Sm53fZJUBWKpoYRm4UysVl1JOpEdZItv8qPsdsdPfOnF52Mtq1adurhSy0Jg7J2//BSwHvXbKlSpXot9Nob93M+tqytv9nszUNoFXME92KlH3+qXXVGX7yhTenZsc18syvYY2sC1csqn0L7XPTe0h/EL9zzPDfm5rjyf/MY+Zy1EOSgyGNcwvnJjK8qin+Aepz/gOCyQGA+jkGQ8Qx/Bc8O4JKGfgRiYK4sIiIAIpCkBKSzSFL9OLgIikIEJMOBlIOxWAGX1GdgykQwVqjGIPmLVZJDR4XgHPsy2msCSlXahGyuCnFDHS+B3eMV3cgy6EZjg+oIKTHppKKsMj2nDlRIFoDhghWp4cFqEI/hG53cvdyWhJ2e1J8IzfvMSCuG7nBXMCPjwgf7cyInTsGZ45aUhR00EcROFwIaycO/k10i3Am7jmlXLm4T4+vbK7xQgmy3Qrdd+VrHxu5sUIgRr07HbUwQEZyI4+Kkenb2C3XqVFbzWTgATyBJUWCE0RtDh3CpxL6Jg4C8CSwQxCAwRhLAilPsWRQOr91ltRj6E3pTBRA8FBQoErFAQyDFp5Bg+kxdhD4Jy53/YWUU4ZQpCFBQWKIeYJKKoQ8DEfhQjoQoLBFbUGyE7QnjqGupiDcE752R1HfVAIUE5PB9OIcPqZiycEMQ7qyL7mBhbiMLDTaBDBTChnw+7RLPrTvtdflYAB56R4IZCtY8lJvBcC8aM7IczfBBe8deNJZ0gwFk3uN/5HipYo7yjBCVRFDYJcRG+sr4D1xwIl08y4RUr1y1o6YkoS3GtRP+Cy7fs1qHRp/GXT/RNLt4NP9HnkUIbjTWZ+96k3qWV161aHrBsCt9cMNblpjSOF1qoD/Y7WrRpj5BquCltvcpp0Oi2O/kdd1EbLN6FV56KVWtc4uJvzH7/7Te98tQ2V3b8ThleyuTQY1zbsESLJAgf8XzfJ1FYYG2AG75osUI4h3MJiBB+8tjhERXgTrFjYTs8LSJc0HN3DXFN5eeuED/xnB8h54Y1K3wtEol9wkpmlCQvvdDvqXCWWPZw/TgPK7ypY6T3E8cTY8KVM3nMsMGxxprifcT7HqsZrEyIU9KiXccnGt1+dwvuX96xHVve0fjH7791ytN4b8Wj8kfoHwL4rC+jj3FCR94t7twBYaY7PmRVPf0e7w02PmNxFijLklMqHK5HhPOHKrf9FN2xKE5DBZ+hlgh+lnnhjEKtAkM/o+APbNZ2xoS8I91Kder1X+j4z30Ob68dS/143yPE5p2Mv3+n7AivS6b77p75VcsWLUzpxpv7usNWxyywidXtKu+YitVqXEr95nwwk/e774a1nVssFMm1oOuTUXI/O+zlqVfUu+Em+gYs5ej3Zr5+dLy1pPCJ8vy7Z8ct7vB6Dvkt/PdIFrFU8+/gQhDGqCzCQUnCexkLjUiWRElpoo4RAREQARHwICCFhW4LERABEUgZAqzIYcKMwDdVNp8Bfaqt/mFVJW44cCkxf/aH+JU/ps0WGaP0CWy2mOykcBcgVWoccjWCb10/9yDu+Kq1LruCzwQE3Pnzj0e5hHFCoy83blhbo/aV1+CiabAFxsYUPrwRTliFgMlPIMRkD8UGwqNf7HwIk1j16+XbGGGlmxh6TTxdYFTOd5wtq5s4c+4iF3AR5UrXdi3ujNf1S3ibgisqEXKECjpw34NQgg0BDgmlmLPGQRCCYAi/wBz3qiVcCCDQRnDExJ0JHgIXykIhgSUQyhcE5bgu4zvWF6x0Q9GBYoSJNMo+FB4krCpY1clkk/t5tiUUHZyXFf4IYTgfn1lF69xRMaln1TTHjrO0yBKKDpQZe1lNan8Dm01KmYRixcKqRep0lMDK5c1If41B6KTbrTR1TYwmZDvKbVYYGz+/zqnWJ6X2tcLl0egX+qPkObwhtJ46a2FAEdnz0TbN3/EJcoqQB4G0bfaYn3gSCg5SxyefHUR/hEDf9B3//Wwu3whw7de2shWrBKyMli9e6ASwMWMoW7Fq4NhTbck/58RlCBYL4QXQX7nz4Jvc7wRX1r+hMfuw0GAFv1c+5zJq9vszPRUaocdUrVk70I+vXbGUZ9l3W7V00UJnZXF36/adoikssBQh0DYF4toqmnsVXD6Rd82KJZ71cBYW5MFdFvXxq6xTbG83yz+v9w3HIQy9sv6NAZaD+nbvFK5YMAPCvG1tVTP7sWx0iqetm/zvE1Zou1hM3Le4KYv1RnFCShQj7br0evaWZi1aUwcWD4wfMbj/kGd6dgkPwh1r2UnNF6vCM2RVPacK7Yv8FAZJrVJ6PQ5lMc8aY9Tf4lyswvuR9yp9P+8OFNgS3BoE1x+ujPCsJ9cN4Sy8KG/Ga7E/t/TpuXLlDsSu+mLBXMZcvttV9Rve7HauWvqFZ/9FDBtnudy+Wx+swLMQh2jS6KGDWEDjF2couTikYjmMYRmzMkZ1llWpeHqdSgREQAQyLwEpLDLvtVfLRUAEUo4AEzjc1yDwQ4iK//0UX3WVcs2JrWQ3Ydu0bs1KP1/lsZV0KNfxJ56IdUpg83Jt4la0Lf70EwTYEbdLzZc5GT6xgKxeGZ2wauPalcubNG/VDgXIq+NGDPHKWyi4ug2hlt8q32JB4de327dtveaGm29nkjhy4NM9vcrDlYCbRG4wa4zwPCXLlA8IxxCq9R8xIRD49odvd2wfYeUxWY11VWw0RlEUXgQXDF/pyeo0t0oPAT/7cfvDhJjV985lEdYW7ON3EquXURY4Fx4IP3hW3Op+5+oHxYiL1+DOzTHOvzSKDOceI7x519gPD1vCyuI9S+M5RwThDBYzJCwwcAUS66rWaFi1PxMTQAnR8/nh484657zzPzZ3bn7KChCh3ETZS6L/Iagyvze46fZmCJoQ6I8a9EyvSDhxE1fK/I5TVryBX6mrE3SXKlehMgpSv/MROJx60C/7WU6giMVtFPlmzZweGoj3iCa4cy7+bF7EfhxLDfeOIbB2tNuK/hYrC1zx0b97ubVyZeS/sEgxBO58x4VJpLK5lihs6HdXLvmc/u6IDes78vBjLMFwLX5FwMLCXMR7Wsyw776HHgu4gkIJNW/W0a61cAvIOREWojCY/N78gKWGxfD2VWwVCokNNcfifMQjXCwRVNjccOudAb/03G8oSob2790tmrIn2nXT/hQnwOIBYjdhseUXeNyvEs76d5tlOMq1ZorXPB2foGyFKhfzHGB1lNLVtLVBgT6D/gWFaKznw5KYvL9afCVnwex3bL2GtzR1+/wWxOS/sDAWr4ENS6up418a+vrEMSOwTo61TgmSz7law7qIfhrFhTYREAEREIFUICCFRSpA1ilEQAQyJQFc2OBaBlc5rAbPsKuK3dXFLQSfWQGcHFf8f2eejT/9LCg/EMSEl+kELusjuNHgGCw/3CrWOe97m8FbSIpDAThNaFfp4lqXEbvCTxnh4k1EMsMvUvyQEAoXMTff2bwVK3z9BIiuPCaRXgGz8xcqgs/pwIarjUljhg764K1pU9LJCla3utL9DXdxRrWjrcSPdLtEW+V/1OrOoMsP4nHgGgoBC1YeB6KsJOU5xa85z+xRFjjJcT+rjMxHoHnbR7tcajEcsOzq1emh+5NCwNyMB/pT8zCF8jviVqJsuYpYaWAVESl4tVchFxYpXtIFX0bxQewKL+sK3IrUb3jrHZSxZOGCucTa8CqvUrWalxKfgX0fB/2bh+fjnYEiAuVINLcmVzdodAtKW5Qkn875ECVkxI3+FndVVWpcenmjJne16NulQ2u/A6y7DsSvQOA4b1ZkZQiBrcmLKxYviwinSCfP29Mmj8d9VaSKOus+gpx75cOiz7kEHGzWFeF58Bl/T5sOnfkdBZPdJlisZSFwuF9QcPY7RQmf358ee7wpFFtOUMl7eea0SeMnjR42yOteiXaNtD/VCTDvx0qJ9xz3fLxu43CjyLuygKUKllhAEe0dneqNTO0T5j3++BN4nrB4jbffTUpd3Xg2YF0ch3Ign8UL4nwb163GpafvhtWbW8SD4tyvTeecdwEWsFm2bFy35ra6tSokU5yKpCBJ6WN4bojZghUei3GIA6ZNBERABEQgFQj4rUxMhVPrFCIgAiKQoQmwChxf/wx0cUOT4TcXBNA8muD655g351bD4syykv6IDaGJha8ITJZwSxHpZA0a396M/SgDELB55XUTQIRRKCqmRPBhXrhYiYD/4EiTPhdwG2EUAVVHD3nuCDcxoXVwLqb8yiPAIvlZuXb7tbUq4hM4tZUVx3wxU6mAoL9h57KKsyKUwfVFtI3n9HJL9S3h1z20jGjHar8IHEWAODMPPNKlJ6tgO7e557Z4BEuhheEbnO95Q4Ks+uF2cRiiuUzyOt5ZL7h9Y4Z4B9K+5Iq69XFVRb75H703068uda69DhdrWYhLQbBwr3wm70JwmuV78xflpZQOPcb14/M/en9mrIGcp7486kXKqHt949uIreBXV4T+7EPw5uUyMPS4qxoccpWCxYxXeaXNfRO/o/wYN/T5ZyI9GtSJOETk8bKu4/fGd977QCCIullghPuSR7HUa+CI8SiRWAU9fuQLz7m27Nj+1Va/uBmU6xQlcMd9VqR6hu47zZRQziKwQc2LCvd5vH0rKStipZfm+Zj3o3AjbgwuHeONMULsK6yFsXw8HEchzVuVxhW4qGLV6liUJcUNX7xVRyGdv+Ahy4Y5PnGB/Mp0CukdX28NxIfz25q1fOhRt88vPhH7Tz3ttMDYateff/6RgZUVNJF3B65Gue9xO4rSQpsIiIAIiEAqEJDCIhUg6xQiIAKZjgB9K+5w8IvParbrLGV4Aejvv+78hStti2YDAamPdXNunLwC/uHjnYkb54gkCDwub97jb7ytWXPyTXtl7EivSRWrgFEqkIcg3tMmjR0ZaZVcbBYWh4KZUh5WEV/Mn0NAY8/tsAJk7SrPVW+2YjYwKfzdJJfHyjSTHI81E4Glv7DEalBWqIcGnT4Cgyk5eF5RVqAYcsHAMwkqNTMlCLA6tfegURMQNPd/stPDkYKWRjv/b2Z6RR7i+ETLWyBojbXBXNtFyxu+v2yFytXcb4vMv7mfC6X6Nx0Kto0w3C/uBO3GsoR8Xi6M3HnMGCDQ70ZT5lxUqWp1F7dnyriRnq76vNo719wnofAhjog73iufGdgFLCz8Apm7Y4hNVM1cTKGE+nDmm1O9ynIurpbZ6udoQcQLmCsqJ/z34o1CAssSzsP7K/x8bTt170PgbNyIEcuIejnl+4/ffYvbH9+taIlDMTs+mzvr/XhcOLr3EcfqnRTvU5bm+XG7iOCVBTXElMEffzwbglpn8ck71S9OUTxlJnzeimZNRiNSQ2FRyMyBnfKV/i0eeDZuJgZJwCWU33FVa9W+Ald6bv+aCPGC8tgAm3xeLlvjqVcC5IUbimXivzCmZHypTQREQAREIBUISGGRCpB1ChEQgUxHAIEp/SsTQoSl7nuGBmGW4wRkDrhgOiPozimpDaYMF4z1velTj/IpfpzZ4FM2fsQjrcxtfEfzBxBWoah4feLYEV71cStNXXmTxwwb7FdvlBtudfHm9WsDgXTDNxQpxKVwv08c9cKASBychYVfAO/Dk8Lde47FtVJSL0UiHueUg9ut8ijPcFUWSWHI84m5PwK+WZa4rhnehVsiXthEqDPKiuGT3pqFshSrqHgE7F7tM5dQARdl5+bLXyBa+52rni0b1h1llRbt2FALi9cmjhnulT+3Wc85YRbCOT+XQ8VLX1TBxXH4xCwi/M4NI/bt+vMPT7dS7rh72zzyOJ+xgFiycP7caG1x+xHgr1p2KOB1sZKHrCi8Nuf+5KvN3pYg7phb77q/DW6p5nwwc/qP33971Op0FDUlyx6KOeQX2yP0/O7dQ0wirxgSBLcmsC3vOc4Zeuy1N97c5I4WbTvwG+6ucEfDZ3cPeNXPHU89nWIjXqGni/WBGy/4xnotlC/dEOBdiPD1Kkvx+uJnEY6zrOCdKdfSBgG3c1zdpZ8vmJfSV9m5cqOvot+I53zu2d2//4BnjC4stTr17EeMscNbpJgc1i0FyjlofUE89UjAvLhjRHGMwg7rlEB7feK+JWDzVGUREAERSL8EpLBIv9dGNRMBEUhcAgg7iWGBgHm1pUyxMp6VmvjNxjT+lrvu8/UXHu2yIkx5vM+AoeRbv3rF0kgrvDgXq1C9ykRR4Xx7T588frRXfAiOY4WqOx7hzfc7vsFPs+dWqFiJUuz42xy3+wnrChUtVpJ6kW+nSRs/fNt7JS77qTsBdfnsFyA1E00Ko90ase5HCFPFEqb7BAbH2imahROm/pdYamwJP8/R8sdaF+XLRARYXT9q6jtzUGoisO7b1T9uQqxYXD9DjAnXr/gd6/qSaAFVw48/0TrLgmbqxe8ogOd//ME7XueoWvPSOigt2Bcp2GudYLBtXDfFEvzbKWW9zsnq5Vp1rq7HvpcG9esdKzeXz60mPvHkk3knH7Wdefa55zkldCRLD6wrbrv7/rZYloz1cfUEQ6z/OMmnc2ZFjbPhhI8oYrzqVqFqDfqkLJs3rF3tXIPxHXeJ3fu/OJrP06eMH/3W1Ilj3fHnB/3UO4tHr3LPPf+CAs6F48K5sbuDoiy9j+K9A9NVfsamxANDiYcVFu/HeDYUFLiSYkNZleld4zjrLWI9RBo7xgM5Ul5TBgeswVYs+fzTeMt0MXfOOufc872OveuBdh0LFC5aPFTZ6beQhuN//vF7rA2yoFSNty4Jlv8vqy/9ubNc9JxzJFibVF0REAERSAgCUlgkxGVSJUVABBKQAMqKmpYqWUJgmtFXIGVBODX91QmBYHT3tGrfyVlIxHvtHujw+JNOUPNcz8cDK0jDN4Q3zr1TqDVDaL4O3fsOMJ3FaSgXhg3o092vHoWKlzzsi3marYiOVF9TWATymnvwLb7lWZBUt2/GqxPHRvLty+TQmfd/s+1LzzIz0aQw3lvFLz/KBlY/4+IG5QUKqEjPH/mZgCLQxF2GNhGIm0DD2++6b9TUd+cgwELg37n1PbexMj7ugsIOMOFRwLUPq2NDAyV7less26wrRsByeKtc/ZLaTe9r/bBfXehvURSzn4DWuBjyylvr8kOKA4T2H787wzOGA/tdkOgVZoURqf+zsEKB+E4I2d35Q8+Lu6SufQcGrD1Y6UsgcK964TLq3raPPO4VpyJ/0E3WLz/+EAheHr65eEP87pQxXvke6f7081jPfTBj2hQ/11GlylWozLEomaK5gyKfs3L46stD1hHhm3mMKslvm9atWen2YQ0yaMyrM2CDMogYEm4f7eedx/dIbg2d0PObbVu3oFT3Orffbz//+ENASMm5nHImnuOVN00J8D5ESYFFE9c9XktC3qsvWSJAPOOVTK/Yr2UxfVAkR3L7mZxXvGipMgFLsa2bN6yLt1znKrBG7SuvCV/og2K4ZfvOPShzwewP3+UvFlR//P4bcUs8N6cYz1egUGGvvhNrtHoNb2n6wsuvv4PCPd76pqP8PCcooulbsWqRZVk6ujiqigiIQMYmIIVFxr6+ap0IiEDaEWBCiPATv/i4BwqsuM/o2+C+3TohBGEC98K4qTNxWxFPm+9u3b7TfQ899gTHsGrUz8QeIdi6lcuXkK/OtdcHgruGbnWvv+m26xo3uYvfnun26IORfPY6CwvM6z+fPweXQL6bc9/0oy2l88vkykOo96atfo1c3iEFiOlU/nCr38Lzu0mhzfcOW4KE5jHvWCfc92DHrs+Pnjwdk/54eGfQvLiqwN1FwN2MbZtiaOfHlocVdHODKcMrGGNgoiwxEEBJ0H/EhNefeGbwSJQK701/bVL75rffmFx+vem7ULpSlUhxGNifO3fugIsXF1yVz9Vq1b5y6CtvfvBwl979/ATMlS6udZlr6qx3pr/m12xW9rOPAM9OkRqel3M7QfwqUzJEQrhhzYple/fu2UMMofJVqtcKz9ux57ODUeqiQOneodU9fmV1fXrQiDYduz3VtPmRSplLr7ymQQUrF8XRos/mzfY63gUqZ5+LARKej5XHWI1gtdD/yc7t/erhrs/yRZ/Nj+HWORz4ese2rzyD4J4SjF/k4piYu6lKzoKHFd0d7mvSEH7uXHny5AlYv7D5KZ3YV+wYhJ6/moLDuWE0l1ae7yRcWfUfOXHalfVvxGJNW/ohwDsR90VYIDJWiFehinUG9xhKD1zVZXo5QqMmd7fg8tLXMRZDEeClfE2OW4Byi5nCkrIiWR77nQtFOvFqiK3WqXf/IW68yBh68LjXZqKERAnq4g5xvkht4T2AVQnWWrc0+3+rahQVxDCa8v6C5cRyQkFywkknJfJiEOZxWEKzsIV5h9yzJscNrTJEQAREIAYC8j0ZAyRlEQEREIEkEDjLjsHfLyvQCmSWiR2CjPturld7sCkrWAn61OCXJl5/yx33TBw1ZMBn8z7+wM/ndbFSZcu179q7v7PKIEjt0107tInEndgW+F1v1vKhRxd9OvdjF9j28roNbnxywLCAiwzcZbz92qSX/cphMlbAohiy/41J40bhlzvSOV3A7UjuNtxKssWfzpuN8uZYy/vonemvP/R4z2cqm5/kMuUrVV29fAnBpLPg/x22KCsQ+OHOJGeunLkirWhOwn2ciIewEi7gU9o2VoTuitIIVs8xAWUVM5NS3BtssxTv6tNEZKU6J4EAgnBbfLqvxmVX1m3U5K4WrLznuRvar/cTfu6CknCaw4ewWh9hNckr+LLL+OvOn39CgUIfOH7E4P4IjfoOGTMJwRT1coqP8LqUr3Ix1oABxem8We+97VVXyriw6KFVspHiUpxzXr4LEFiR76stkWNCoKT9xM6HwKxL3+eHtbzt+itRhHA8CgiEgSh+e3du1zJSWYsWzPsYZXKrR7r0xGKA/hmrkib3tmpHPWa8PullP3/vxUsfCrjNVq/RrXeMHzn4Oefahet6f7vHuuFakHdDj0da3bPTTAz8rmXJshWwqMyydsWyxdGuN5Y4Ls7HP//s8uyjXFwLlE5Nmrdq17L94z1QCNG+1nc0vCbcOgKe1O/0/511dq0rrqk/c9qUCVzT8LoUK3XIrcya5UsXRatn+H44zH5vxhuwQpHTfuntN7r3psXxrtCiXadul11V7/pDHOIvP976KH9cBPZabix+UWyifCDFs6GoYGX/z5ZwKxWvwiOec6X7vFh2la98qO/s3m/ISyRXaca6e02beOj/ew79tU+HP9tvR+xnn23Yr9HXolwmTtDgvt07uTLPu6DAhfzOc56UZ5cx4msTxgynL8Ei8Ip6N9y0d8/u3fQXnAPL5a7tWtzpzsfCI1zm+cXDoW9+beLo4Q926tG3XZdez/JexLKLGEYoRSiHcz71+MMPrFp6KJZQgm4o91ygbbmDStCLqGqLgAgkJgEpLBLzuqnWIiAC6Z8AQgIEoBdYYmVnphF+Mrm5u+FVNRFc3H7vAw8RkJCE4GTDmpXLEb45Qcz/zJluKRPCsYrWXVLcfvR8tE1z4mFEusy4n2raom378/LlL/jS1HfnLvxk9od5baUXK2o5jpXOvTo9dH+kMhDusSqOc73+SmR3UJTjYlhYfHFfRYRzUTXBlDTRbtPCQXdUkcojmDnKHoLdjnz1ndmLP/tkjs1nc6K8cCupv9y0fm3nNvfeHikAebS6ZJD9KAjzBtvCM4jlRDShilMqYpnBpJTjMs3zmkGue6o1A3c6A80lT+gJEcYQr4L+LSUqgjIWZUVoP+l1ni/mz/0IQTLCI4RILubFh2+/MXXIM08GAleHb6wIdsGfp0+ZMMZvZT7KCudGZMHsDwIuQ7w2k/EfXuX//Y7tvvGA3LEjBj7T8xITdKHonTZ70Vpcq6B8oK1YRjzb/bGHZr4+eXwkri8PH9QPaz4sEno9P+IIBTXs+vd4LKC48NqKBX3Cr1+9chkC98nvLVj22dyP3idvlRqXXI4wD4F8r8cebOGnzCEvrIuWKFWWz1g/RLsPQl0ZmmGMZ/BjAoxj2YHyH5dUlIlQsVXTG692QbbDz/PK6GGDuPa8L54b9cob99/aoE54Hmdh8YUp+qPV02s/QsprzdULCrHXPvp89dZNG9bhestZFyKcHTds4LNcl6SUr2OSn8Dyb/5EiVjAEkoKXLFhURivaxvyE1gai2FiWaAAybQbygMUEzz7uERlAUyOnPafDdCwVjjkou5wdxg3p3/CXPs564q3TQGb1IUpQ559skv+CwsXxW0fSlNXqWVmFfbkI63vdRa9KG3POT9fftzS+SksOBbFeMky5Sqi/HCuXPkdy8BpNqaeOOrF5yO5p4sbStodsNZOjdtQLNo0Pky766Azi4AIZDICUlhksguu5oqACKQKAQSgDGoRfG60hM/TTLUxeRv41BMdp748aigrueo1vLUpQUtxPRLqfsRBQSC0xATxCDlQPMQCCyVDu7tvuQ6hDMIf5zed1acjBj7dc8rYES9EK4cVYqxWe65n5/ahQU29jmPVb3abgbJvpQnB/MpG4Ic7K+cHOFIdnEm+sw7xy9vD3KEMn/zWLIR6LgAtefFjPGHkkAFMYP2sV6IxyID7cT3A88dfFBARrWbK5zvpgAlzcLmzwhK++wM+2rWJgBcB86jxH30PfRaWXfRxsfZZSSX6usXWuanp3fevCVpX+ZUzpF/PrqUs8DeujRCi4f5jsvWDg5/uEbAQ8DqufNXqtYiHgBJ5nE8waY6z0AiBwKoItNavXoEPe8/tG9tPX/S7dagEi47WZoK6dnnwvqasTib4N4Ivjvlq88b1T3d7tO2iBdGF6sSMMCF+XcrAWs8dP23S2JGvjhv1op9wj/NZ/OkLyd+9fcu7+plrL4R519zQ+HZXb9r7pClGTR63AAAgAElEQVTQUR5EassZpthwftwjuSB0ZWAdASeEmhamxHOM8MYr40aiBMACZZ8tzcaly/ABfXv4CRB7T1ycdXiPu55DiX/jrXfe6xYGhNabALlYdhDom7gg0a6P137cxjzfq8sj7br27sc7yVkVcr+9bzE+xgx5rm8sMTyScm4dc0wEWCmOkopFNDstMVaNV/i61Y7BtRTvysPuyI6pVgl6MIrNi4ueffyBgwcOhI+/UO6ivM1jprC4CrR/eflOX2v/8tjnPDntgz3+puLImRPtRpZgHCHGkMSK4TkLRbP9qy83Y2E35JkensrnWDDy7mrb7KZ6KN7NuLiUGXrs3rRu9crw53X4gD49Lr60zlVLFi6I2O/R7kdb3tkYd3j0vbSbBTRYh2SgMSkKOmK+4Ar2qyQ8M7FcGuURAREQARHwIJDpg2XprhABERCB5CZgwk/6Vnye9g1OCCfb33dMMBrvarbkrlqalsdqrZJlylc0uc65J550yilZTQHw15+//47bJAQnkYL7Rao4grlylarVMBnMBT//9OP3q5Z+sTCadUZSQaB0wdQdf8XJEVAXCwkC6W4yoZ2X647QeiLYqlrzsivOv6DghfgYwIcxwr6ktiUjHmfPHs0qZOlRS5dYesTSB5b22/Pn22Q7Dlc3rDYkWDEr6QJWGZGOyYj81KbYCKBo3G/SGBSesR1x7LnwE+4X5ya0dBSrZ517Xj4EYybH/yZSLAOOI+D1nfe37fDem69NQsjkV1NWD9e+uv4NCKOiCaNZafuLRdRGwBZry7F04zhW/fJOoH9LCl+ORzkTrT+lXriNGvnqzNm4UbqiQpFz6I/r3tD4NtNhFOZ9ZC6NFi/6dN7H0VwFujbiissO27nsi08/iaXdxPrIZRcKX/DR8psy4ogsXZsG4nsHNhQV9ofkYgoceHvcM3ka3PWYWw3MvgN2zAGUKl36PD8M6weuZbTzRtp/rml7KlSrcQmKn+++2b4NpY6f27FjOY+OPXYC9o5jsQXui5zV73/2fvsl1pKD71aXHQEuCtBA/6f3ZKwUlS/RCATve8aH1S3hDhCFH8o63feJdjFVXxEQgYQkIIVFQl42VVoERCA9EwgOcE+zOhI8+lxLKC5WsZI7PddbdROBRCcQfPbwwYBQhoCwuL0I+OmOorDAHRQWGfjoZuWpJqOJfjOo/qlCICgsP+JcJhhPNUXOsTTyjhZtO7R/4qn+uHpqd88t1x1LWSl9rJ/CIkRZgRAZoTTKVhLXAAUGq+rZx2/0b1kS5fqkNNPMVL69G7kHiNGE2zIsejbZOxG3TtpEQAR8CATHlFjh8dzg4hBXv4G5nBR1um1EQAREIOUJyCVUyjPWGURABDInAQa0Ljjn31JWZM6bQK1OEwL41UYgg3AuIKCLttnzucsmpuSNFu8iWlHaLwKZgkBQgO4WPh12LZNIwvASZcpV4GIlQnDoUIsKd4MFlRUEgSVhwUn/xV+3OAKlRcC6wpJTaOzjuES6TpnigUr5RqK4Khq8P86yv7hA1CYCIhCdAO59sRbc4fpWKSuiQ1MOERABEUgOAlJYJAdFlSECIiACRxNAgPC9pQ2WfhYgERCBVCPglA74HI55pXdmd9mWaldHJ0p4AiHKiiOer0QTghcvVbY8F2PtyqVRXTKl04uGBQVjDf6iqA13O8n14XeUFsz5nMXFfruGuIiKuX9Mp+1XtWInwPXfZgnF1V/2vtsd+6HKKQKZmgAKCxa06JnJ1LeBGi8CIpAWBKSwSAvqOqcIiEBmIIBbGvycsiIHv/jaREAEUoeAE8Kxqlhu2FKH+TGfJcS1kKcQ1WuF+TGfVAUkiUDwWoRep4QTfBMIN78FJwdALDEkkgQqBQ+y58UpH3Lbaf62axIpRtZBy48iF2F13mC/+J/9ts+Ok1VZCl6ndFQ0iqttlvibqYNlp6NroqqkcwJBS4p9ZoGrsWQ6v1aqngiIQMYk4IKzZczWqVUiIAIikHYEdtmp8Xf6pQ14JRBIu+ugM2dOAjxzh4UyMt9PmJsg4QTfCUNWFT2CQNGSZS4iQPmOr7/6kgDbiYQnqKxgDne8JawnogqgCbht+VBqILBGcYGiI5tXDJJEYqG6xkyA6/6PvQsJti3ha8zYlFEEAvEqDgSTYlfohhABERCBVCQgC4tUhK1TiYAIZCoCKCy2WJJ1Raa67GpsWhIIUUxI8J2WF8Ln3OGBg0Oyyad+OrxeGblKJUoH41ckpjsolBTOwgJBdKyLIsiHWxMXz4IyDscfycjXO7O3TUqKzH4HqP0iIAIiIAIikHgEZGGReNdMNRYBEUgMAggR8HsaqyAhMVqlWoqACIiACIhAghMoXjoYv2LFsoSKXxG0iEDJgIVEHkuMNWLagjEr3JiERWscnzNosRFTGcokAiIgAiIgAiIgAiIgAqlBQBYWqUFZ5xABEchUBIKrvGVyn6muuhorAiKQRAJa4Z1EcDos6QRKli1fiaPXrFi6KOmlpMmRPC85LRGLglhZcS0+wzWUKShwIUWwbhQWuImKFP8iTRqpk4qACIiACIiACIiACGRuAlJYZO7rr9aLgAiIgAiIgAiIQKoQ8AmcLfddqUJfJ3EEcuXOk6dQ0RKl9u/bt2/d6hVLE4yMe15QMjjXUPEq/f6zYymH41hcwV9tIiACIiACIiACIiACIpBuCMS1Kifd1FoVEQEREAEREAEREAEREAEREIE4CZQoc1GF7Dly5Ni8Ye3q3f/9+2+ch6eH7C6A9j/BysSl9Au6hsLKAndSJFmEpoerqjqIgAiIgAiIgAiIgAgcJiCFhW4GERABERABERABERABERCBTEGgTPlKVWnomuVLvkjQBqOgIBYFCguCaMe94RrKDiIxF8wRjI1xuBz7noWkTQREQAREQAREQAREQATSgoAUFmlBXecUAREQAREQAREQAREQARFIdQJlyleuxkkTMH6FY4WyApdQWEkkOf5EUGkRl3VGql8snVAEREAEREAEREAERCBTEpDCIlNedjVaBERABERABERABNKeACu7tZI77a9DZqpBucrVatDeVcsWf55o7Q66c0LJQEoOd1ZYWaAA0SYCIiACIiACIiACIiAC6YaAFBbp5lKoIiIgAiIgAiIgAiKQeQiEu6HJPC1XS9OKwDnn58t/5tnnnvfrLz//9NWWjevTqh7HeF7nEsopLpJcXIgCJMll6EAREAEREAEREAEREAERSG4COZK7QJUnAiIgAiIgAiIgAiIgAtEIBIWl0bJpvwgkG4HylS+uSWHLvvj0k2QrNJUL4rkxZV9yWkXILVQqX0OdTgREQAREQAREQAREIDIBKSx0h4iACIiACIiACIiACIiACGR4AhWq1riERi79fMG8DNBYlBbHbC3vpTi03zIAHjVBBERABERABERABEQgUQkc8yA3URuueouACIiACIiACIiACIiACGQeAhWqVK9Fa5csXDA3kVsdomQgBoU2ERABERABERABERABERABERABERABERABERABERABERCBRCLQ8clnB7Vs37lHItVZdRUBERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABEUhlAllT+Xw6nQiIgAiIgAiIgAiIgAgcRaD3xMXut2z2IZelfcEfDtrfA5b467l1bVpZREVABERABERABERABERABERABDIAgRwZoA1qggiIgAiIgAiIgAiIQIITQOlgSguUFSyoYYya2xKKC77vtbQn+He//SVpEwEREAH6DUchdDHeYQWnFJq6SURABERABERABEQgsQhIYZFY10u1FQEREAEREAEREIEMS8AEiwdM+IjQcbelPJYQOvI9r6WcllBaYHmBwoLPES0vMiwoNUwEMhGBEIWEV6udkoK/pOzBfoM+gu/qIzLRvaKmioAIiIAIiIAIZAwCrGLTJgIiIAIiIAIiIAIiIALpgoApLVBSoJT429KvlnZa+sXSP5b+tYSigjzOGkMuTtPFlVMlRCDVCYQqKZyy4jirBclZaGVDCRpUhKZ6BXVCERABERABERABERCB+AnIwiJ+ZjpCBERABERABERABEQgGQl4rKAOj1fBKmlWTLN62llYaOV0Ml4DFSUCCUbAKStQXLqECzkss0Jdxh3+bP3MgaBCNMGaquqKgAiIgAiIgAiIQOYiIIVF5rreaq0IiIAIiIAIiIAIpDsCPj7mndLioAka+ewEj6HKDN9A3OmukaqQCIhAchFAWeEsrOgDUF6izERhwYYlFr85RYbLj3WW4t8k11VQOSIgAiIgAiIgAiKQQgRkQp9CYFWsCIiACIiACIiACIiACIiACIjAsRHwsMBy7p9YfBdqYXGSfccCy8XBwY0c7qGIf0NcHL7vk5XFsV0PHS0CIiACIiACIiACKU1AMSxSmrDKFwEREAEREAEREAEREAEREAERSE4CzGOxqsiWI0e2XDmyZ8O64vhs2bKebOlE+3yapVODCcUGSgvcRWVXPIvkvAwqSwREQAREQAREQASSn4BcQiU/U5UoAiIgAiIgAiIgAiIgAiIgAiKQDATCXcY5i4tcObNnOy5Pzv0HDmY57sC+g7mzZd+fPWvWrCdmPXgwy559B/7JcvAgSowDBw4e3Gt/mfdieYEFhuLfJMN1UREiIAIiIAIiIAIikFIEZGGRUmRVrgiIgAiIgAiIgAiIgAiIgAiIQLITMEVFtrzH5cp1Qp6cpx2XM9v/jj8+5zkn5s15Vq7sWfNlz5GtZI7sWQqapUWxrNmyVrK/ZawCZ1rCIgNLC1lZJPsVUYEiIAIiIAIiIAIikHwEZGGRfCxVkgiIgAiIgAiIgAiIgAiIgAiIQAoSKFrgjKx//b07a47s2U/JljXLSdmyZTt134GDBQ8eyJI3R44sp5vJxUlZc+b4et/+A79mzZrlxOzZsv20Z++B/fv2789t5hbEssDSgkTAbm0iIAIiIAIiIAIiIALpjICCbqezC6LqiIAIiIAIiIAIiIAIiIAIiIAIHE1g+Td/Zv3jr/9y/PTr37nN/VPRA/v3n7Z3f5bTs+fIUvC/f/advnvf3rwHDmbNa/v+3L9//7a9e/fnzZI167cHDxz83dxE7Tt44MBPptD42kr+zdJeBeDWXSYCIiACIiACIiAC6Y+ALCzS3zVRjURABERABERABERABERABERABEIIoKzY+fs/uXf/H3tvHqxZkpb35Vm//a51a6+u6qV67+nZeuhmNmDGDAwgVgtJSEEIB0TINoEjrH9kKUJ2hI35wwrJIcIOY8uCsC0MDiNLNgIsQNIwiPEwg2aGmZ7eu5au/d6qusu3ndXP76sve25XV01vtdzlPVFZ59zznSXPczLzZL5PPu87LlKpJmbjODiUu/q+IHKLcvt0XxFXc1UQSUtRl1XlFqIkTsd5Wbuy6iishQ5xJxXAgvHvqlJfiXgWprKwUmYIGAKGgCFgCBgChsAWQ8BiWGyxF2LZMQQMAUPAEDAEDAFDwBAwBAwBQ8AQeCMC5y6th3lZJWVdd2tXH9Wvh/Kiev84Kz8wHmWHh1mxZzgqZ0fjcq6oqo5cCRxvpcnxZhofiuOwF0dhHLgAwuKgUk8pUABv8zhgBc0QMAQMAUPAEDAEDIEthoApLLbYC7HsGAKGgCFgCBgChoAhYAgYAoaAIWAIfAsBEQvhxZWNpNtptKSJ6NV1fU+W1x3FqWiKoGgHoRu4OlB8ironyUQauiiVyqKZJsG4KkPkFedHRdWMoiorq4myIlVqKw117VLrGyot5DLKXoMhYAgYAoaAIWAIGAKGwB1GwAiLOwy43c4QMAQMAUPAEDAEDAFDwBAwBAwBQ+DtITBVQQT9YdYK43Ch20jmKueSUZYtjEbFbFVXnSiImmVVLkkuMRMGwdC5slQg7qQogzyMgrAOgp7kFfeVYfhqFFYSatQd3T1XGlkci7f3HuwoQ8AQMAQMAUPAEDAE7hQCRljcKaTtPoaAIWAIGAKGgCFgCBgChsAuRECxBzY/9cQFzweOzFjsgF1YFt7lI1NmwtG4aAZuvJSPy0WREIpTUe/J62omrOsM0iIryrQoKpdEUa6YFQMF3u4Egf4Mw4YUGaM6DLpaPxJqR1WXp3UMcSxiESI3jWVhCot3+cbsNEPAEDAEDAFDwBAwBN4DAkZYvAfw7FRDwBAwBAwBQ8AQMAQMAUPAEHhHCEBUWNyAdwTZrj+Y8tJR/OzZICv2RXE434yjjlw8NYqsSIlrcc1NVNAWi8F2JwiDUmRFKfIizfJyRoEbAykuSpW8A3EQXNKPl0VeNHXdRClTkmjDAnDv+pJmABgChoAhYAgYAobAlkDACIst8RosE4aAIWAIGAKGgCFgCBgChsCuQaCW6gIjtFdbYCy2xRC4KQIKmh1EoUviOIpEQsyUtdtTV/X+2gW9WrEq5OIpjuOgTOOoEDkR6veG9g3rqgzC0LUS6SykuFiXd6iwqqq9Qe1e08106GQJzC2UFT5DwBAwBAwBQ8AQMAS2DgJGWGydd2E5MQQMAUPAEDAEDAFDwBAwBLY1AlMi4u26fIKwSHQOQY8LcxO1rV/9e868XDPd6BoTUktsQyHCoairajDOi7Ao6wVREFmaRGtSSgwCkRadRhzpwErBK9K6KFFOxGkSDgIXQohdEeFxwsXu7Dhz64ppseLqWkG6J6SZuSd7z2/PLmAIGAKGgCFgCBgChsCtQ8AIi1uHpV3JEDAEDAFDwBAwBAwBQ8AQeBMCNzHEctzNXCO9wYC6zfzov10DMM/o3UOlgCHiwkgLqz83QqAOw6AoymqAZycVliSJg4FCUVyQymJWRMaeSFRFVpZ1Piprgm0HLkhFUJSoLIoyh/Doyk1UjxgXin0x0k28CyhzUWZlzhAwBAwBQ8AQMAQMgS2GgBEWW+yFWHYMAUPAEDAEDAFDwBAwBHYFArij8W6R/LY3oqI48Mu2mf3t3TxJKfF2XTxxXK7EmIQZ8biKKk1psSvK/5se8ibEXC3CT4qKSmErQikqwpFYiJHiWPQVu2JGKomRVBbDvCwDuYYK5fEpiII6TMJgwGZVuZ4qlwJwO3EX9ZLIiheVMlU86hUKCx+/YneCbk9tCBgChoAhYAgYAobAFkTACIst+FIsS4aAIWAIGAKGgCFgCBgCOweBzYZYGV8hKSAoIqXG1FDP38z6Zk3STHIHacGxGPXfLgGwFUALRTrUm0kLbX+7fBVTl1CbCZxtQ9JsBcB3Qx6kjCikknDDURGHURCndXS1oYDaZV0vKuWqKIpuEcptVN1UjIraaVuuoYb6LdZvmdQYp8OgXgld+NKoLl/VIdQxIyt2Q+GxZzQEDAFDwBAwBAyBbYeAERbb7pVZhg0BQ8AQMAQMAUPAEDAEtiMCzBSfEhKoCSAs5pS6ShhP+Q0Cg/45BAX7Jts6DxXCTY34W8hllCdi3inBwrNxzsRFFkoNU1lsxxJ+2/JM2RhmeSkeIrgQhtFJ/X2orEo5gApyxbDIg9CNakksRGzUKkyhU7ALMRWrCsLdyIsykhLD6Zc1eY2CzxgqXdU1IAlZUHG8KfNbqF7dNmDtwoaAIWAIGAKGgCFgCGxFBIyw2IpvxfJkCBgChoAhYAgYAoaAIbBjEJiqKngeDPrEa5hVarGW//2mJo5DTvSYCS5jK8b7RRlU+d3PAMeQz/ZWVx5gWPbKkHf6/jbHtHin59rxOxgBEQcQCpQruXVymerLJRETx4pJhQouB5FrKISF3D4pckVYH0qiQIG2g7J2dZHE7He5jt/Qyefzos5Ut3x9wiVUzfV3MHz2aIaAIWAIGAKGgCFgCGw7BIyw2HavzDJsCBgChoAhYAgYAoaAIbBdEJiSFRhIISraSi25tllSAOB52Upnw8D1ZFg9JANrImvrOfncH2lfGrjqhAys2GQ5tzOxzV7zuf9O1Qt3EiryinKEhby/m2USBNlUFu8Gup1/DrEocgXOVkG7KtdQK0EUrVZFXUSpa6iCdLU/yPNK3IWOVIDusixPxzH1SuqKonq5qqtTQumCEgQgy+Z4MTsfQHtCQ8AQMAQMAUPAEDAEtgECRlhsg5dkWTQEDAFDwBAwBAwBQ8AQ2H4IbCIrcAE1ryDAPfnZFxkhV1CBW5I//YeD2jXqMLgUR8GCiIuj8lxzXscOqiocK2LwabmxGWl2OMZVCI9cs8G3OmHhY3S87Rd2gxgXNuP9baO3qw5EHXFe9QhXTiPpjXoi9y5WoUvk56kn91Crcht1WYVnJAJwSa6i5kUOigis11WvzunvFUXlPl+58orOn5B/pq7YVeXHHtYQMAQMAUPAEDAEtgkCEz+xthgChoAhYAgYAoaAIWAIGAKGwK1FYBqzArKCdFjG03aSRLPqgO+T65rDgQufTJMwaTTiZRlUFzUdXAqM6ETg6ovafknuay5kWTEoyuoFnQ9hgeuowVYlLVBFKH9MiEJlMbY4FLe2PO32q00JQMpWKtJiSQqKuTQO5frJzadx3I3jYC4ryrZIjW5d1kty/LRXdW5V5OCLUjN9RQqLc0EYroyzwsiK3V6Y7PkNAUPAEDAEDAFDYEsjgLTcFkPAEDAEDAFDwBAwBAwBQ8AQuPUIYMD3AbabMpwe0YzwQ0kS3N9tN/crLTQbcVtBhA+3G42Hu63G4U4zfrjdSB5XsOB7kyD4iJQXD8ZReHBKAhCUO50SIbc+t7fmij4Wxa25ml3FEJgiMFVD4MIJpYVUSFVfbtOusj3O84GCa6OcOKMA21dEVpzV9pfLqvpyWVZ/JuXFaRcEV0RWfNsA9ga2IWAIGAKGgCFgCBgChsDdR8AUFnf/HVgODAFDwBAwBAwBQ8AQMAR2GALT2eBMDiJuRVcu9R+II7e33Ur3p0n8xFyvVY5G2b2jrKiTNF7tNNPHms24kpubK5oJPnNlY/jcaFRcCmoFCq7Kk8NReVpKi5O61roSSotiK7qzkcqCGfCk3BQWO6xQb5HHmdYtiEBUR4nUFnu0no/CYBJEW8QEyoqhBrprRVUNoiBcH+fFmn4rVWcgLGwxBAwBQ8AQMAQMAUPAENjCCJjCYgu/HMuaIWAIGAKGgCFgCBgChsD2RGBKJni1geynQUd+9SMZU5tBUO8virzRaMZBs5F0e+20kqKi30qjWC6iDsdJeKjdiB/utNLOnoVua6bTWpzptTIpLV4Pur0VyQrelEgKZsAXRlZsz3K7HXI9LfsQD8SykNKiXlY6K7XFQGlViooXFPflVZEVr6niXRBZsUGZnKbt8IiWR0PAEDAEDAFDwBAwBHY1Aqaw2NWv3x7eEDAEDAFDwBAwBAwBQ+B2ILBJYdHV9RcUbPvhNIkacgG1T8TDj8x0GnGnnTY0HzzMyypvJvHRKA4iBd4eyuDaGA3Ls3VQP99Io/PDUXFKhtivnr+0MRxn+Yq2VzDWbtVYFrcDz9txzek78peGXNo8Nno98Ldwvh23t2veAgSm7tG8qoc1hNn1bslQVrDfFkPAEDAEDAFDwBAwBAyBbYAAQfFsMQQMAUPAEDAEdgUC9e9P3JQcDz7tnuOB9fc+rVb190jbLE2lWaULU0Ae1vpF/W6Gjl1RQuwhDYFbjgAGcMX5lbYicFkjiZoz7caGtsNOO1lMkrgZujpMXVRFYZgURRmmaRQVaqqGrpit6+rh9X5Za2loxvjeRiP88yBM1vqDrLrlOd3BF7yOmOBJPTGB2pzxEHjSzk/e1/Rv9r1OWuxgeLb1o01Ju0rvGAWFf7e8w9dJi62qRtrWwFvmDQFDwBAwBAwBQ8AQuI0IGGFxG8G1SxsChoAhYAjcHQREPuDbGuPFvBKkxONK9ypdUir1OwFsv0fpgNKc/iaQLQvuVq4qnVP6Q6XDSs/o9yWtX1X6uhJkBoE9YxEZ5gv77rxiu6shsOURwEgqIypG00yExVUREplYi2EziXJZwq+Ixph1VdULwiBtpPEFKSvqyoVzURTNiKAokzQs8iJoxXF1tK7drFQZF8IwfEl++ofLQVCt92mubAEB4XwzIG6kJmcf5DXvhnVPiX0A6g3duBqifYfQ4DgjiLZ4UdtEShjJtMXflWXPEDAEDAFDwBAwBAyBt0LACIu3Qsh+NwQMAUPAENjyCIhQwMh0RGlOCbJiM0lxWn+jlIC8uKgEWfFn032HpgYpb+36kP5mH9fhmh9UOqu0VwnS4/j0PhPyQveFvMCoBclxWgSGGUq2fGnZnRlUIOSJ4dbiCtzx9+9neQdRFIwUdLvXaMSNqq5XRFwcSqIwlZ/9tCrrZqU3lIahYlzQ+tQjgl604qgXRIHc89enw9BdyvM6zotiZq7XvGKExbfe5fUumzYpKjaTE4x7PIFBIHTIChbad4iJU9N9qOwuKxHQmfeX63q08zclLcxl1B2vV3ZDQ8AQMAQMAUPAEDAEDIEdjIARFjv45dqjGQKGgCGwixBo6VlRS/yHShikMEYRZBMXT5AVrCEsjrkoHboyQ10BsZEpoZZ4/xQrtjFWHVWC2MCghcqCY/kNUgSSgvt9RGmghEHrv1Nanv69i2C3R90qCIiQuFlWvIF2suY4Iy3u6FubGLzlzimUQmJVEopFxaA40GqlcTNNc5ERYTXOJbko5+M4HNUuGFdlpUPDdquRykJelbE8RJVFNS8Fxrqam3F/WMxJgfHaHX2K7XczyjskBG033wP+hoCg7WYhrgjjIL4BENR8I/gNgprfOA8XUavT47xbwC2ptJjW/8Dq9vYrqJZjQ8AQMAQMAUPAEDAEDAlOZYsAACAASURBVIE3I2BBt61UGAKGgCFgCGxbBKRwwJXHp5W+T+keJRQUGJowPj0wNT7hCmrddR7Z48J27OY/3nJRJ3PpfpmqruYu6bXd1T+66Fa/NHDjkx0di1oCwxaJ63vf5hiu+Bt1BWTGS0rebQgzdJmd+7tKvy+lhQyLthgCdweBzf76P/joQYy27sBSD8M5BlrW3vham4Hz9r8jvQ+Iz0arEc93Oq2D+xfbh7qt5IONNPlYGAWPZHnZqKs6jCI3UPztoeJbBLGUFVVRl6OsyKKwvjzKy2WxGKclunh+fWP8u0kcPfdDTx2m/bHlOgQ2BWHG1R+Jdh2FBN+FPdPtOQQsIn58W00bDrFxUol2HmyfV8JNFNcgyDluBn1A5zfc9W4rLDxhQaasTluVMAQMAUPAEDAEDAFDwBDY7giYwmK7v0HLvyFgCBgCuwgBERQYnFA/kB5TelQJgyykwteUcOHEt40YFFdc5+GDbv57apfsPeDSPbELZXcavjR2reNtF7YKkRhNl1+qXPuBwHUe7bq1LyVu5XciF8u+VfQhLJi2joH32kzdeGHFVaMlVw1QW2DQQtWBEQsXUwtKP6j0WeXzWa2/oYTx6yRBvXfRa7JHvUsIQFSImAh7nUZwdW0UNRtxNBwXwXicVzJwh/MzTWaQyzAeYoTFgDuWobMyA+dtf2G0T+M0ja90G1HDhcEBxaSI9F76SSPuS02h0BV1opZGREXYlCuoUIb0rKqrPIp0YBj2GrVb03srtH88021KdRGGeneh3t2WnPF/2xG9yQ2mZB0EkVdWzGgbIgI1HPuEXNAVKbSkd0B9EPkcjIWr+ItAbXgtjCfHUz9QsUBUD6ftvB833ZC0uFvPzH1VDliZS8K7+RLs3oaAIWAIGAKGgCFgCBgCtwwBIyxuGZR2IUPAEDAEDIHbhYAIAAgDyImnlXDxdL8SM2OJVbGo9IoS5AAzYQeued9ht/iphus8IfJhflZkReUGz4cumInd7EdLl+wLXbGcKcZt5rpPLbrm/ftERFRu30+l7r7/ouVGLxbuyp8ULkhl4CraLmhVrnnPuitWei67sOza9+3Rb0dcOcjc1X89clXddGtfWHTFVVQezMQlH59QelnpOeX/C1o/K+LCjIu3q5Ds8utiqJ3tNeOxZutHo6yVJpE8CkXFcJznvXaD+AndjUFWySCeySAbQmbI6E0/sJDhe2ikxe0rQNPg29Vst5nPzLRyxa0ogjjM4yhYC+rgguiJbhiETYXcbsriHCqJpqjFW7hEAbiLMHAbUlxcUSCLdb27V5MYR1LBRDljy7cQmJIVlGnaXwhntlFX4OJprLKv0CBBqf86wnhJuCqFErc4BQmpFA89yLVfm3VLpn+2n6L9ViIOEgsEB2Qf7gZtMQQMAUPAEDAEDAFDwBAwBAyB24SAuYS6TcDaZQ0BQ8AQMATePQIy8KNWOKaEsYnYE0wf/ZQShidUFny/ICk+oMTsVwxKEBiPuMUfmnWN+YbrfaTl0sU5VwxecN2H92nibNs1DssdVFt2qFhGq1kZs+rS1ZmsWA1dt9SMWpmwXLns6v4Zl68uyF18w619ed01Dsy5Klt1dS6SozgyIUCK9cCVV6SckOEwXz3h8pXArf4Jx+u3lS+5usIVFTNeUVdg4PoDJRQbqDP6SidEYBDY1RZD4C0RkDH22x0zUVb0R3lDoRF63XaaKEjzHqkq5FKoHGOM7bZkv601i1+ltdNKg1YzCfX7umabD5tpzCzy191E3ehG0xncb5lPO+DGCPzm518NG2kcdTvJohqce9XQPJqmyUdFTIgsrY7VQdjW+ymLuirERrREVrgwDGPFs7ii1u55VwenZFtfFWHxhbKqXi1Ld1aKmb4pLK7hPSUr+C5AVviYFazvU1qYkD9BOB8lgdryoF25+qgYIdF2QVPVQ6k+I0XLa2qx50sIC7XTejevCW/aaFR055Ugo4lxcUUk1Dsmn79dnBkjDK3lMAQMAUPAEDAEDAFDwBAwBL6FgBEWVhoMAUPAEDAEtgwCIiqYEUtA7MeViBMBOYEhFQKDGBGQAPgXZx8GIwz/uIdqurj3ojv4cw9KCdGRi6fYjc+ed53HDruoN1TMitrFe2SxTSKXNCE3jikxQ5lrMRP3BSXuTcBt7gWpgIupl93w5Rm5jzrqRqdLF8aLioOxX6SFVBVZKoVF5KJmIMJiQ9szbvzchsv7592VP+67/ldGIjEgLCBSiHuB+gLjF+5KIDEwfH1d6Q9FXGAQs8UQeMcIYKh98NieKC+qZL0/TpuNaDFw4XynnczKCLtPaa9+0+9lniThRqORjGW5Vfl152SYfa3bSUMRHJdFYjBznHrliYs35MUIi3f8at50wr/4szPR3Eyjq8Db9xeVu0/06NNyRdQrK3dvFLhDZV2jvkjl+kkGc+ktapfpGBGpwYkwdH8uY3qmBuWLZV09L+P7OREgIyMsrsF8nboCYpuFtv0BkRWPiyR6QKqURNv3y/tTLYznpVRRsO060L/BKC8uiZzoS4nUFPBD4fyi6s5J7cNdFEQz35oz08T3oUA5895LhV3BEDAEDAFDwBAwBAwBQ8AQMASuR8BcQlmZMAQMAUPAENgSCIis+EllBB/jP6f0fytBWvA3RqIjSg8qYfxnpiukQjbN+EBkxUvuvl/8lNv46gkRFj0RFR0XNS671oNjF8284qLkO3Qs3zxmznJdDFoYoCAP8FV+XAmlBgYu7oebqSWle13rfgiO2jUO/pmryuOuvHzODU8kLr8yp2gAIjDmOi5YkapjYdUVS4HrPnPQdY5nbnCqcOd/7Vk3eIFgrriw4voYuA5N73lB67+jtFfPnou0+I3p89jKEHhbCEyNtCFkRa+TdqWk2CMD60NJHB6SexuRb/WDYeRaipAQ67f1olAchCBfzVy4Ns6LUK7M5PbMlWvr4/FIkZ8pn6fOrVZmiH1b8L/jg6aBzwd6X6sKWPFaWdbf1Cz+xaisB4qgUJZiMWRQn1UIC5GxdR66eigFjF6py4qipL1aiaNoHAfhQPEwMiMr3vAKmIRFoo2FfIOMhuCmvd0rQBfiMGiTpD7qSQGn+hK1iAsSRqFL6no/8UEIZCHZnYQuCisSBJmUGCu64iVdFBUSCgvqibnjesel304wBAwBQ8AQMAQMAUPAEDAE3j4CRli8fazsSEPAEDAEDIHbgICM9e/XZVFJPKGEwgGD0yeVDitBFmgW7MRAhC9xvlvEsCCoNq4/+m7xM203/31Pu5lnOq73wUOu+6SOj066mcNPiVDAuIQfcgxYJ5RwEYLhj/0QHhAYkBSoNzBscX1cUHE8Cg+OwfBFLAoFy41ec+HSWCTFgisufNGNL35kkp/GEREgyYKb3R+4uCWjWTVys9/VFtmxx61/+QV34X9/1Y1Pcz2ehWtCwPCMPCtkyqpwQHVBgO6vaG2LIfC2EFica2viuEtlZ51TXIqDmip+n3Yc1uzwg0HtFoMwHMgeG2uGfqwZ+Zrc71rDYTaT56Vs5W7h/Gj9vArhWCmY7TTGMqrjvsyTgW8rD3bQ20ZgMiNfhBJt0FwYlH2FEynyuhrrXSRxHMyInVBw6KovY/mqLOa8F8nC3KgOo0LCgPNR5JajKKZ9escuid52LrfngWDrlWoQ0pAVT4sAylQ3RPSE+6We2CvCJ1ED3SgK3KNRHVwoMq+hYzpgr4vkOmesD86sIoUc0pfiUCV3UiIz/pWO5VsBKcJ9+IbcMmWc3EV5suWG6JvCaXsWSsu1IWAIGAKGgCFgCBgChsC7Q8AIi3eHm51lCBgChoAh8B4QkHEesuHHlFAykPYovab0pJIMdhNjHAZ8DPwYhvZPbwexwExXXCv1XOveU+7Y33rGtY+3XNBMXdCbcXHCtw3FBOdDUGBkwsDHPVijqMA4hHqD6z2gdGB6fe4NYYELENxRLU/Ph5jgeO57RYqNposOzykmRunytROyW71P4TByNz4zdkE3ct3HegrUHbuyv+z2/+QxN/sd97mzv1a5K//ypLgM7k3eeEbud0zp80qf5n7C5mNaM5P3t0RekF9bDIGbItBpw1UEzf4wa4uk2COhxKNVWe9vNOKWjLSJVBRzYRSUSRRv9AfjhgqfvEPVySgr9ur4Nc32f0XGWQISF6NEc/3rOv4Hv/XVqwrQnZvS4rYUPOo9pFBfZNJJ6Sdm0yRsyj2XlGPRhlikWbkvUjsSoLIYyog+kuG8ioN6UFXBebkzok0amLripu8GgnnftP2mbiypbJ8QUXFKvp/ukaettoKDVJFa56Kqw6Ks5CYqqBQvpJQaqVD5z5M0KVWP8MnVVfjzy2VV9FRv7hWZARHCN4DvQ4jCyerIbakjdlFDwBAwBAwBQ8AQMAQMgV2OgBEWu7wA2OMbAoaAIXCnEZBBHhLiM0qfVcJNEgQCs2EJsE1wbRL7Mez5GazEmEANgbH/eaWu2/vjz7t7/+5nXfPonMiBF0UiQHxAKhCdGLUGs8QvKRE7AoIA4gOXUlwH5QZGw/dNn597s0BwMFMXoxdriAwIDE8u4IoKFQhkxkNKX3fJDO6e+q4qEhd0ui5/9ZSLDyifxYzb+6N7nOyMrnlvw7XvV3yLv/mQO/XfnHFX/jATmQGBQl4wfnEtSBmUJCg92F8Jq98TaXF1mjdbGQLXIxCOx0UzCoMZGV73N5L4vkYSHZCxuyW1xUgqil5VBw1ZXvNYFts6L1r45E/joFeW4ewor5Z1LmU7i+JIXnDqvtiMSgZcFACVDLKlGWRvXaGbBlYuNZseovKkVBSX9K6Oyki+SJBtvZsVvYxuUAezIi5o64YiLzCQV2EQXlLQ7YFcGNE23jDOyK3L6ba8kiehIcNpu4kzQfsvkiFIBW4oRHM53SoTxbJQfBBQHGvdVKOrsl8pfkWYC/dQkc/RXqje1J0gdKdVHwBEf9Zgz7eE79ItVbhY0O1tWeYs04aAIWAIGAKGgCFgCBgCtwkBIyxuE7B2WUPAEDAEDIE3IiDjO0QErpCIVQGJAHEBEfHdSigJIC0wBEE6KAZFZ9W1jnddY1/lZj+euuahsSvWUVX0XPuRnmvc85BICs7D4I+7JUgGDP6oIVhzP4iIE0oT458SMSv4DXdTbEMMsMZ85RN/+4V9GMDIF9tcE8UGx5BwN8W3dE0BuS8p7XfJY0uau9vU0YGrNoYumFeMCzntad7bdtXzI3fv3z7i5j/Rd6f/wciNznjjF8/O9iNKuB7hGb5f6THhRmyL0yIueE5bDIHXEcAdVBSHcssvOU+s6O/aSJJoWJZVrLSkWfsdWWIDGWJVHuWtzAWJnPNr1rj8Q0VRmSoySx0FSbORHNJs8myYFRdEcpQiLiD2MMheM+vacjsQAN+J2ksLqjGFsXBjkRVn5fpJM/rDvhQBalukrwhcX2TGRb3HizqOduyWuSK6HQ92F6/p1SuQzBC9L+IOSuTDYi0RhZrsfhjWubDsqXTjBipQVWiKowNj/l4XwScvXdW6C+QySm7WdNJh7b+kuBe8qEykBWQe781ivdzFF223NgQMAUPAEDAEDAFDwBDY2QgYYbGz3689nSFgCBgCWwIBGd1x0fFxJQzxKAk8EfDo1PjTd+nBQ66x94xb+tFlV6zucelS14VyN95+ZMGFCqBdJd90Cw/ud439zDjmehAGJ5Vw6YRaAiLBu5JCKUFQawgJHwOD33HpAbEBgcExkBcQJJ6s4PzrCQsMhBwDWcFxE/WDkidXwJhrcgzkRuJkRdb6Jd16n8tH65q/m7jiaiUCZlYuoQrX/cDI3f9LsYKEn3dn/7GUFysQOLiB4jww4Trk8ZjSTyt9URj+kUgLnskWQ2CCgAgLubKRg/0ojIbjYkaBmdkeaacUQIqpXZZrimkh4UXY08zxhbKuWiIx8mxYiByrJaoIU9ETipNQr2i/zq8gxeZkvN0nNzq5/i6ksjDD7K0vb5sJUgzrBHueuK8T9qr3GM5rVBW+HVjVftQCEEkE257EwrDlTQjQfoIN6/uE2WNabwRBvaAY2scVs2KhyuteEVRqrwONgRRcW2zyNFQ3UiNCnCuGBbjXV6Rxc4pfIY9q+OdSoO5r3wba/kmA+tuFvxQ4XHoi6/D3sRgWtwttu64hYAgYAoaAIWAIGAKGwFZEwAiLrfhWLE+GgCFgCOwgBGRoX9Lj/IISJAMLhh9mqeLC6bSL5x52i5+dc70nMze+cEx/i6zYtyIVgiiBlcglR8+7xkHc3Dwk2xLXwhjllRJcg28Zhj0MfxAS1xQP14gRDHyoLLgfKgbcRHEsBAcGJ/mNn+TPu5vi2n7xBiOuCZngSQk/89wTGygjvKHMz0z3Bq3KJc2hCAv5TT84lgFs7KJu0/WeUsyNaMF1pMZo3bfszvwPX3XrXyUPPA+xPB5UYjY1eWc2L2qLDwrLvy/SAsOlLYbABIEkjsZyZ7MyHOcXtK3A8EG3Lqr2aJwVURj2FGw7zauqGWnKOGqMsiqluHBiAiNt16mUFUezrByqsJ8V+bGm+Bevqa6NpLKA4Ju4vjHS4tYWNggHGaV94GbaINos6j+kBW1UKrEMRCt1n3aN9sTH37mlrohu7ZPd9av5tpk2Gbd9OHOSW756v1xBLdWliApJJMQ/5Crr4vEUtSKopEhSUAv59AvVUAdxWCs4t2K9RGkVVK+JBIxwE6XrLOiDsVfXhDCHnL5tKhfIiSlpwTfqDcTFXUfYMmAIGAJbHoEPfeyv0m7QR2VN8t8N38fdPEmn/vLn/9fbRsBuebAsg4aAIWAIGAJbFgEjLLbsq7GMGQKGgCGwvRGYBtb+Tj0FqgqMcCgVIAtIGH5G7sBfkyOOozMKXi0Vwih2s08vu/YDiQvbMtTFV9zMx3AZ9R1K55Rw+4ThjvMxRmEwwojHQAvjHgG0cQXiB2SQDAzUUEZ445J35+FVFsSo8LNmOc8bvDjPD+D89fkd3/Oe3PCGJIyMbJMvFgyM3I/EvraIFgXqDld0J+JTSEGi568HG3JzJVdR//6M3EU96U7+0tfclc8x8/2MjnlYCYIFVzHkiecEw58Rrl/U+t9aQO4p2rt8td4fla1GOhA5cULExZKEE+NGGhUbgxxyoinDdzYeZwPRFM2gDEpmi5d1IPdPeaxCK44Dv/3X6odsufs1s/+CiIwNERa+j0jZMyP5eyxnUwP05quAKe0G+HrygjaSBFnkCQofw4Zjc1NX3PRF0E575RtkL+36IZXnh/QDxO9KJMJbH5BxFLhVpUYlDk9niKOrCTYvPrlOA/mECqOwjGMn9VE4JKaL6sKymI8VHQJZTJt8y2O73KB8bP7++G/NeyyFNz9dpOTmH6+/X61YNrft3nZhQ8AQePcIiJygb8o3wxMTrJlow6QdyFvvwpS4PvS96cdChhOPDdXuuq5B/9K7Pn1TZkRovPsM2pmGgCFgCBgChsC7RMAIi3cJnJ1mCBgChoAhcHMEZFTHiP8ppe9VYhsjP4MllA1fVzruDvzMcTfzxAddcrDlGodCuUW66srLQxf1vu5SuYaKZ35Axz2u5A16zGrlu8XADGMO2wy4IDEYaHnXTxiUGKyhsoDYYHDGgA3SgwGcj0nhg7OiioDUwNjllRI83PUzW/ndu2jxv5MP7k1e/GxYr4pAKeF/J6g2AbuvKTziJHdlO3NVS880StzMU/PuoV/5iDv1Xy+7i//0EbnE4riJD3YlnptnRnWBMZP4G11h/AciLXg2W3YpAi+cWK6XFjquKOo4TaIkTSWnSJLDCqStieH1qcEgW1PoipEMsAuNOF4kkHNRlrHc26yXZS3vUYp/EYaDcV4OyrLMtG8gsiKRYdarmIyouL1ly8cI8YZ2P+uVNs2Tp96INGmPbmDYnuRwt7sMIji8jO7eHRTfhbbK8QkRDUeIVSFdRanyP5bPpzkJJqSoCEZRXTelnajC2um3sJT/p6FUFXU+rksxe4r/Ut8jl1EojgbaPj8lLWhzb7m64i3e352Y/ey/d9evKV4e28n2jaqEERq3t6Gwq+98BEQa0NcjVSIIIBpeX6aKCf729ZPjPBGxh/ZOie82RATfD4gJJuY8q0Q/mD4q3xT6yR9WekKJiTG/r/R5JfqcZ5X85BjuP/n+o77g/qbC2Pll0J7QEDAEDIGthsBtn7Gz1R7Y8mMIGAKGgCFwexGQIZ1B019QIoA0hnpcLqEaYCD0kEv373EzH0ld97HI7fuJlsuvKCBwrYDVzefc7HfOSo0AqYDywc8Yw3CPsZ/BGYQHgy8Sg6llJa+48OoH9jHYYn3f9DgfkJvZZOQHUoFjJoPDKSIM6K5XVng5PQNA/9vmtf+O+tgXnmhQ/IqJmoJrejUH25ApGNMweEGgtOWFZL8rRkO3/idn3MbXm2747HPuzK9qf8YAlGfm+Z+fPifXZJYvf39T6Z+LtDCj8vQF7sbVf///fCOe6Ta6ijlxpN1Il5I0/F6ZFBf7g/yl1Y3Rw61GdKio3B6FEk7HeT6bZSp6QXi5KqtCLvq7sj5uaHb5VxWv4lRWlGvapmw9q1nlwEl9g/jLMAhvZXyvM+S/aYb4VjfoK//XE6Te5dyEuNjq+d8KZUOEBRjSzkJAsxBI+1EFK/+EyAa+KXKMVt8vDUVHPp4aIjSW5P5JHtNcv6or2ni5SlOjK/mFiLxcRMXZIi9eFs/3bFFVKNvOKObLZdWFNxgTt8Kzv5c8THHb7ELG1/Ww2YDTDKokiiq1JxNXh1u9LXgvWNi5hsCdRmBKRqAO9mpf359kko/v39HPpR9MP5o2DsKBvizbR5ToU9JXpO7S/6QNZHIL6UfVlhWq4BKR1cf1N/1nv9Bn/S0l9v8vSs9Nr8N9mHSDKpmFfj3tHu0E7QDL630CU2BsQtQ2DQFDwBAwBG4ZAqawuGVQ2oUMAUPAEDAEpgj8Ja1RRjDDCyMRgyMGPU0XJG239ENDkRZ9N/vMUVeOz7v00D0KsH3ZJYsY8hkgMUOMWWAMjiAtcO0EscAsMgZt+BD3AzXuwfEMphigYVxlUIcSYeJ/f3oNXISQFwaFfPsYcHEeg69XlSA2vELielcc/A3R4IOuavMNSgyvzPBKD/LBzDWuS4JkIC8E1oZsII/HlFCBnJbxOHFJe8bNfvJe1zq46vJnDrqgXbvXfvnPFROWexL7gzyDoY/RwfX4DVLjn5AhW3YnAk8/eaR88cTKqNWMrzQasSJqF69JMTEny0QvTsK1LK8P5pJOlEUtOYUKrkIIa6Z5qlVW5FJUlHKMU9dyH1XFWoeaSa7fJ4QedYh6RdmbBN/W+g2kxRadVe1Jxs2kBTEjMPpvZdJlc968a4/dWajf5VNPVRa0jRBt3jXgmkrtNwgyr+Z+RQEsLkdhrTY2OKL9IoadCAv5hRJ7IWJjLHIiC+qw1MmnFI37lTqMXlP882/oS3JBdQU1Ht+NnbZQ3rySrxD52RBh2ZVSaz2Ookgu5hL9XXXbKW1CprYgN9JipxUBe567iAB9PO/Sju/t5hht1Dn+xiXqJ5W+poS7UPqskAz0lelj06+kf6lmK3hMRO33aP1EEOjUulTItERRqxJXZCPNkZl8yp/Tmn4qfWz67CyPKf2OEmQF9/yyEn1Y2jz+pk8OKXJCiQlBkB02YWYKnq0MAUPAEDAEbj0CRljcekztioaAIWAI7FoEpK74jB6emV+QDxjXvRHkg5PBT7p34Br797l4X9O17p9x2aWzrnX8qgsjjO8MnH50uvaDIa7DYI5g1AzoUFFgTGXxBIOflQZhgAHfG/cZXGHkZxAHWeBnq3nDK8chgec3rsH5GLrIC9uci4GKPHBfrsc2x/JcPg+sveqC+5MvnoXBH7PbmJkLieEVHQwwGYQywPSByOUKK+669HjlopVD7uDPNl26p+nWv7LqLv/BuiuucPyHptclb2DLYPEJMJfK4vem+bHVLkMAI/xvfv7VYjgsNhQ8O83L6qKMi8M8L7t5UQ1lbB1pvniQpjLDBuFQzm6act2/VpTFRReULcW50CFuoBnk+PHPVJLFZ0zKNwZfypgnALY6sj6f3tjj2wf/HLhTmtTTrUhcXKeg2MrEypYuB5tIi4l7FZXpRGQcBr11OYbKxUucUlTtURqHnVKMsHxBzUrhR3RueU6TpyjVAdF7ZVAFl4sgOCeSYk1V46o4P9rgHRXPZaqs8N+viRu4Rho3FLZjr1QVMzJ6ro6zois3cmmrkaxLhbWCe6y5meZI506MlUZcbOnqYJnb4ghIXcH3yrsGZE1fEcUEfUn6n/T16JM+qfRR1T/6j/fRYGmmwRM6Qc1WhLu7lvY8qQA894VIxPTZjtLUJQ11l3VslCQK1lO64dVlrSdzdcRg6MZVMSEw1ASSDdpJ+uB+eVobn1PyblhpU5lU9KvT/NGn9jHb7Ju1xcuaZc8QMAQMge2IgLmE2o5vzfJsCBgChsAWQ0BGc2JU/GdKDGiY9YUkHeMOQbdZGCGdck/8+jOu/XCkEdKGaz3QUpwKb3zne3R+OghiH0oIiAmUESgUuBZ/cxxunSAZ/MLx3p0T+7zPd4gJzodseGV6TdwwMTsN4xN55tpcl8RxXJ/BGddAyQHZwXE+QCH54rooLpjxxuINo2x74sLPOuMa7CMfmuU7uS8ur3CVdU1hcQ0vrs99/z+lJ1zRH7rs7MANX113w5cTd+GfvOyufp6BrCdK/q22UZs8oEScC87/RREXXN+WXYaACItQBEUiA+OsZkfPj8bFcRkav1NGx4OaOb5XltheGoVNWTYG/YFCp9T1hoy4pzcGGQaKXH+vyGbxioy7l5UwQlBeMZZQ7yDWRjJMejcQdw3dm8VvUIYwtvpZ4hh6qL/ePRAGIZ6DBSMrdcW7WTIjy117m7f3xjKo802g7cbYd0iF4UNBKOlaDXHhHlaw+Xu13VIdWdB6pDqgePROMS6CyzL+ZYp5cVZSoz+XsOC0/n5ZhAXfgrHqwY6ZUbzJXmUX1wAAIABJREFUFRQvoycsltrNNBSDmYjczITX/DjL56WymE/TKFebclrtQ5HG0eXhuFzO8oLvjZEWt7co29V3MAIiLOh70vdjMoy4hYB+4WelvD2g7T9RXXxKPUx+k1vV+seCKH4xTpsvaj0s8+z7VU/fHzeaUi/jxi5aD6OYNi8usrFLOz2XNK/N7xHp6sosc/loXSHUdHgUOZ2vNBaBUei30eRvjpuyFx51+rC4ifrXSke5ttIfKzG5h+8prklx+YoSeuIy7kavy1xG7eBCbI9mCBgChsBtRMAUFrcRXLu0IWAIGAK7AQGRFcz4+nklXC5h5GTAgssmBjQY9nHldNYd+9uHXb5BzIrAzXzsjzTlC4M7g6v3K2FwRJ7OdwklwpeUGGlh3GcGF0ZHBnUYSBi8oX7gfB94cPMscK7ljUqsITgwNmGcxZB5Qumk0qeVMMaSZ67jXS95wyx54978fkoJooNBGWQDxAXXxBiGAdSrPrwbEm9AxfiLAZVBKIEOmZ32BSWuzTUgTMijD55NYO3IxZ2BC+9LRVYsuCAO3NKPLrhibc1tfA0sUZ+AOdcEa3Bg/9/Uu/iHIi3Isy27CIG/+LF7q3/0e89NfFi3w5S68JqMHc9OJlaG4bJmRjerIJzXTEr5gSo0MVNlDJ/WoWaRF5Mg28SuWFHCsE+dpZ5RrimXNzVCbBGIN7uAYrulWfESmtRDBSLvSW0iL1d1qR8iVZYU9Qm7mmmciQApt6LaYovgut2z4dtVysQVvfvnZYi7R/ViLwQFSgvVga6M9GdFUrwmki8RMdHUfGXKvfym1CdFeb2gukM7T53ADdKOISs2vVy+IfKGFbQVrKILMTHf61Lv21fXBw+UZfhYEodjtQ09GUfvFyF6Tn+fE7ExkipL7rTqUsRHaUqL7V5dLP93EgERFfQR6Rsy+WastujBIHQKGBNpO/q+KE7vkVpij0iEz2jCQSuMkt8QmZCEcfJQ2uz2qyJ7Jmm0HtDf4h4SNVdqmoKgp7+lp4xco6tmL9RnXhcPwnBCRMRSXIThzOTvKG1p3pA0ZkoQFqP1Ky5McleMh/Ig5VUXNA01LlaZeETfl7zS5/2EEkQFfQ7axj9VQuXL5Bn67zYR4E4WJruXIWAIGAI7GAEjLHbwy7VHMwQMAUPgdiMwJSv+su7jB1/MuMKADsGArB0D/Ddc2L7HdR9vuc5jp133CYwhH1BiVhYkB4M2CAgGPqy9/1wf6Jo1Bn6Og7TgfO7nVQmbY06wPXFtMV1jYML4+htKj07zA4Hx3dP7QYhAZPA99IoMyACufUIJUsDHv4DcgFQhn/54xoMM4Bik8dwsXnHBmhgbHEu+yRODP8gNyBzyxbN4lwDci2uTn54Gmxfd4vdpStzKftf/5hG39qcjV41fc4PnyQPPSH64Jwls2PeX9U5+3UiL6ZvYRav/4DMPlyItXCOJRD7IOF8peHbgKlQXURzMyIC/NsryObmJKmUAGWka9ZqcQKn8VpTNZRkkKcOUR+owC3WAba9Y2spoemWUvF5Ulfz8dIejrKjrNMjyMhpqmninlcovv2vpOXMZXN16fzxxFSXSYvJ8Rlxs5df7zvMGuSBDOu+Y90s5vqh64eMXnSVmhZi7gwpIn4i4O4MfNBQXdVnNaXNFxsPXZAP0hDVtNYb5G2Zki8Zy+bagTdUV4OMJbwj0/VJgfUDE5pVmM9F3LbhHJMZD+pCN1Z7kcqm1R4SFvpM4xXdLUlqIAC37B5Z6fLfvugLrnZcSO8MQuHMITEkK6hx9PPqZD2lSwYNxI7iq9feq/XkqjOqZuJUccVUoMsHti5J2V2SFK4v8r+mbnYpcdSIrHpeSQrxGLBKiIaIhVXXEC5T+V8M16YJqe0JiqFkT8RGI3Lj2oH7NtlQWLJAWE2mwMsB2Ph67cf/KRHVBfJ+p4uIHdAj9Ux+z7YS26YPirpUJM/RraUtoa60tuHPFyu5kCBgChsCORsAIix39eu3hDAFDwBC47Qg8wzhH6WPTgQrGewZijI4YDZ0UWTF2+386c3Pfc9A19mL4QbHAMQxykJjzN7JzjsdlEwYmBjzM5uLaKCr4m+MY6JEw0LOw/9qo61uzutjnFQ7cg1lff12Jbx4KB0gEVBIYZCEJIDBYcx1/r69qm2d5frr/helv5A8DL/lmYIbaAZUEAzXGfH4GrncNhRsn7/t8Ml1NCVdSzFb7/PQ6H51emzyjyCB/XIdzP69g5AOXHui5I//xXnf+Nzuuzs+74SvgR/48ScK5vIP/U4l3QuBEW3YZApAWcg8l42K1ojDCG7I9XMLlzWCY71fB68puf0CubVwk46PcQ52XAXJietRvGGa9L2rWlG3v8mEru3x5PW6FiJg0ywrNUA3b8rm/T0TF3qwcpVVZReIuDuR5HSRxoEmmcaljB8wYF5mzvro+6s/2muU0vsVNZ9BfF2Nil5Wsbfu4tLe0817519N778iWJ+UNxHitsq5ZySIu1DJnKkx92ezOaP2q/j4j9QB1oS9CwpN42xaIm2TcE/sdGThn5fo+lkH0nqyoHqsGeSpib6gUiNyRi6igUvxtCPfHFLh8QUTFTF3Wf5Yk0em1jfFYBMhWbid22nuz59mCCIiQuFGuvPtt+o30M+nX0QdM1Q49ql7jD8Rp8ERrNjg4FB0QKPzE0lF9o9OqGFyN2uvLasKYgaAvV5A2NY/lmlfQuKUqqzUERRjStRUBK0UFi9o4VdEJebFZeXxTxDgvadM0atJCVSqKTTsSK+JKESHZsC9XUTShNcG8J/F+Jjdz7lNKryrRRtInpx9LBug70+elH2+LIWAIGAKGgCHwnhAwwuI9wWcnGwKGgCGwexHQTH5k4gTZJrg0oyjUEhjimWk179qPlG72mS+49n2PuYUfuODiBb45DGRQOrAwcIPYgASAZGBUhPEfcgAVATM+IRC8YgEDvVdQcD6DMQZIfkDoj/NumTgGtQaDQ/ZxfwaMLOSXvDCr3AfKxijFccwW5bq/qoTRFkIDd1EQAV5NQV5xFcKzcg/O45rs9ySCJzC8T31PpHAO14GkwfUVOPjnJSYFgz8MQ+TtfUpXXeOeSoPFV9zeHz/mkpkvuAu//rgbvMzzTAKfKjHLDfLkx5W+oXezKpUFcS5s2WUI4B5KxvfshRPL5dmL6/jExjC7pnVHRsdL8o2UitAI5QziEh6i5KOf8khZ80ZdSDOMDaTtYISk7qUypODeR259qo4IisbqxjhppjKnxm4hy6pZxR7V89X5OC/SbjNZ0cz6NC/Ki3INFev4gda+DdqJbn92fC24ifqBbwLlmLLt4/soEL07rLJAub8gu94rVT35drGoTa7P6+9z+tLQ9tOe7+TZwnyjQsXzUHzxQER50JOC4opIzf0yXqbYO8VWtPX/DEwgLub027rwq5IkyOSLZlb7+q1mMu4PM3AyI+WOr2n2gO8AAb5N9GHpE/r+rnd/ekz+Gv9Oe7528wdrxZuILskb1ELSqIaNbl2MB625YhxMXDTFiZQUClMRy40TLp8gDVijoJDyabIWOUHdm9h1pJJYl/qC+72TBZJDvqLiXBkMwkYjVN9gQpBI3XGt512LtPjWwqQd2k3i1ZFQYPyQ0j9T+hOlZ5XWFLvC3EO9k7dgxxoChoAhYAi8AQEjLKxAGAKGgCFgCLxjBGQQ/2GdhFslH9eBAQoxITIXzz3nWvcdd40DQzfz/lhuoM4o0PaCBkIYAonjgBGIWVkY+EkMrCAp+CYxAOIYFvYjQce4z2+QCFzDG+oZBGIkwRAFEeFVDQyQcG3jFQgMGFEt4IKK+x1TImgghIt3x0RQbogFjvFEw8e1jSLjaSXIBWbIoVx4Sgljlo8/wUDRD+TIG/f2brH8tbiPDw7uFSQ8348pEe/Du5jyyhAf+Jv1ZUUiOOSS/RddNTwt0uJ+19JY8dVfPKOg3AwUcWuFNP/3lSBVeCd/Ue9oSaQFg0dbdhkCuDfCr7zcIMk+X5YEE1ZBLHAHRVnVf1ktlYFmkIMMdcIb6SEuvAudLWdouF7lsCkIt4ypQUNBgWc2hrlUSG5mMMr3SmXRkNea5jgrm8Jgj1xFjaS46ATzbYJaDLNRsV8upIJmIxnqAoliXhDTwgiLnVVfKMe8U09csP26Co9pxfobQsO7i4Kwox5M3KFthWDzt/l1KNh4MCRFodvfSOJGGVV75EJuIc/RY01i3KTE+BB/UUt20VeTsjeO5SVf9lR5YPuagm8XimmBy6yNXYDXbX4ddvntigCBpaWy8KoG2hMm3aBEGKt+5Wpq6Kei9v20vDS5mf2p2/dA6Wb25bUEDfMiB6LO/LA7Hoxc2irksSmecAQD9ZbzUaE0cM3e3ERJId+HIhMUo8Lri6dkBdgpRgWTaN7p4t3DqYcg3iJM6irMgrTdnRAihdxDXReMG3kHEwVw+8qEGSYrMRmJ+BZ/qPQ/K9H/pK9siyFgCBgChoAh8K4QMMLiXcFmJxkChoAhsHsRkCH8+/X0kBVe2s6QCSN5z3XeN3KLn3rYdR8rXeOBddd7eF6TM1/T9DAIA4xAKCoYTB2frtnHTNfvUoK08C6WMNR7l02b3R55NQX7vCEKRQKLd7mEQYqBIUQGefRxLzjnmBL5hVwhNgXHsB/S4OXpmv3MDuM49p9QYiDGfTB0kX9v4OI7CjHCPbk/53jFBqQMZIlfyIcnVcABzDAWQ3BgTMPNE8+PKywf6JiBICTE8y5uH3bBA2tu9MoJFy/Ou8P/0YI78UuPuXyZPKDIAGOux7kMHr9b7yoTaWHuoTa9hN2ySRBcGRC9AofHRjlEOfOKHx8DhrLCfso1+3zMinqbBNKtNbu7FhnRGGXlweEon2kkoUvj8NhABEbLxbXsOo3xuIhUSQsZYfeu9UczcRyf13zSoaINK7RHuab54wXBuEWCTNoRIy62V015izgSxLPgvWI887FaaCtp02mzfd3gGL4JEz/su8D4Tl1XbApXi9hbjfWfotrs19+Lcg/VEGmRaXJ1W6RnLsdxmeyp8qzvmgoMfF9eFpmiWTRkiM3kXm5d4XohzfmW7WRFyvaqFJbbO4rAlKygXaE/Rr/ykIz6D0icdFAswoeCuvrwxAGjuotz+yu3dIxA2MSNqOSrsIqrMnLtOdxBuf7aBdcfD9zeZi9wSbrhVi9K1lRd88g0UT7JRZsutFnxcO1Z6/pr6okuvK47fhcIILRIO71ccTKCIh9HUmuEuVxD5UOaz2tCZgJ1qx1AzRGLiMH1Kn1Vv9DvRnHRFyb/L22qKS3exYuwUwwBQ8AQMATey+fM0DMEDAFDwBDYbQjIAP4RPfN/qoRxHOMELoyGrnnkObf3Rz7sln4ydcMXM9c6Hrp4/nOu+yiujnxgaUgKjKUYiXy8BgxF3iUNhncMpqeUUFpwDIMyfmdAhLEfgz6GfQxKPpA1rpkwOnEcBhg/58wTDFyHPGyOL8G5GK5OT6/FAItr4/6JUZmPd/HE9Dz+Zj/EBWQGqgsMvBAjDE69kWbzAJL8QmywMIglb9yXxOLdZ/nnZD/X4T4MdsGCPGFAkwsT9+Xp/qsuv7Doln+3587/2rq7/K9QgYDtN5WeVIIMQXkB1pAvf0+kxRen97TVLkNgU3Bdr2iiXFCeMTB6dQVljfLKOidg8XaBSQRDpDgU8zLiEDB4/+Wrgz3tdnJUE1gf6A+LvUVBvS/HMho5GV6XpCrJOu3GOI6DvuJa/Gm7lf47NQ2XNUN8tdWMITD6cg81MVhbIO7tUgreXj6ndYFyTvn3bgK9ym7iqJ33roQrtF1heBcmSRJHh1U9Dsu10wMC57NFVT1c1UFXttVQCopUBsmBDKRRQw7WcAslD/ml9g0l0NqIk/Arqmt/UBTVF6XgOinyMNsmROfbKzTv8qhpWdt89jQastsuRPC7fPLdedo0oDbtCn3V71JiAkwkNcRfSZrtj0dJ430iJvSV3TgZhuXR+58eu/nDtVw+iU3v1K6zgIohzlozuYiCen39UrT27B90k/b88MjMUh1vrHTdlXP7xEf0yjBM1WbVaq+CawEt6vrfiMFgoguTYPziXaS+2xdypSrzLxXj/kw5Ht9fleNWPh52ikwfVJEVlT6sKDyuuaWadBcURCPItcO7WQULlMw/oUQ/thJpsW36Fe8WNDvPEDAEDAFD4NYiYAqLW4unXc0QMAQMgR2LgMgKXA/9DSVk7j749Cuudf8xt/hDH3AzH8nd+FTPpQqs3X3kqmJWMHgifgSDFbYxxHvlAIMpDPQYTwnch/H/fiUM9RASDO498eDVC5zDvbkG53mDEoYmjP9cj2MZuEGEYLiHJNis0PDBwCEBOB9i5F8pHVFigAn5gCqC879LCcMlg0IGYfcpQQ4wIIUQODb9nbyTV+9SxCtJeAbySZ4wDnNviJNrg8xrz+JdRpEfH+ODNS6ouC6xM84qQYxAwDyudMIl+865pR/b72Y+fNC98J8susu//zXtB2PuiXsrroc7LfL6N/TuTom0OD+9r612IAI38eHPk3olEvWEsuhnZnqf85RB76ZsO8SseP3tTQNlRzKU1gPpJERGyPVTIJKifjiv6qPjomrLmCJXN9GGZo83ZVSd06EbQmQ8GhWzg3F+uKzKMzPtVlOGF80UdStSYKyKsDDDyg6sI1NDOsojT9DRvnvVHk88ee+7xeD+LTKzhpuI5QBKjvFdQ/VpTgTfSMjIc00g5zO1/slrTVU3JrEtnARNVSAPUjo6DhdEatxTVu4Fnce3yhM/O7AEvfUjbSLFODhqNxNcbtUz3XQymUHu59w/++KpQu766pWrdAdc9ZMfv8/am7eGdksccZPA2rxb+nP0tx5R+qze+delTPi41p8VYeHiRkvBq+XqqRkd3aOeWqMbydNnIddP1bgzXwW9pSKuq1xqhhpSsNmaKRbb88X6xiXXjxt13FkoiiipX11fTg/m42SPnDteVj28KJJA6g3FK0PlcE11AYFRSLeBmzf1JUmTQNwn9Td95GNvAaTvH5yO4ngtijvjaK6Sx8SoDuPBk6vn241inLjxxtqEqNB91DpMmgcJSKrNE3K4zZPK02cmhIqb9D/pG9tiCBgChoAhYAi8bQSMsHjbUNmBhoAhYAjsegS+TwhgsMfIg6F/j1v4VOi6jy+4+e9ZVRDohpv/7jUXNmXo6KAs8O6fMKRjFEIyvvm7gxEeBQAqDQgCjPsQD96QiuED5QMkgnelhCGe67KwD0UE5AGkB2oIjPycA4HAtr8fa2+4Jf+QGCTUGe9XYjAFUQFxgRsoCAZPqGD4h0CACIAMQcnB8Z4wwfUTxAL5hYwgf342pZ/N691WkTdvIGNgSD45lv08m1dbsCb/5Bl1BX8T24Prg9eyxqFfc9mlRXfkF7oKbP6ke+1XvjLNB8d6oghcwJh396tKtuxQBN7CJc5k5riMaZv992+OUcGs3205o1wuoEL50G+oUjVFSsymadVJolCWm2CUiMGIo3iIYUXunpqaFi6jbNnbkAspBTxtaWa53H0HseKKqj6Fp3XaF+Mooq76WB5bLo7HDi2+d/SxPHFxR2+6dW+mmdHhUCqJVF8m2SgD8Q7BQK5r9D2T7kIeaTSJWt/MulmpAqn+VFIzyQjvSlWePAy1L3cHZRA9onPoH4xxv7VbSJ/Nr3VKVvBNjxTrQ3HKXSqc2oqNEwrDWKROEjZdKRUK/Z1hmkZlllWVCIz8ngNz3hXfDUvK9fF7tm5x2rk5uwFZQV/Ox36gD/ghpSMiBn4qjFOXtDrXXCfpAxM32iIn2iIqYteaW3brlxbrKO73Z/cPVpu9cjYICXL/LewIf92aqfKk4V4WYVE0VwMR6mXZWbh6aeVkeLl/tUM/lP6yvlfBD6ueEkvi2hUgJqp6LBLhigJmP8/+KE5UpyPcNL3VouxzQvmIotksqU6f7y5WCvlUDprd/Pfas8knVk435qJ40Y3WVyexLThBqqsbXTfR3r+F8kLtw/8l/Hwcujd8V4n9YYshYAgYAoaAIXAjBIywsHJhCBgChoAh8JYIaIb+L+igTyoxiwzD/Lrb/5N9t++n5jSOSVzUzd3s03s1aPq8ax476KIG5IRcrThFh37d/QbnYUjHGAhZgUEeAzyDLMgCSA6vrOA+KDLY7wc5nI8x0RMRXiUBweBjYaCC4DzID4wCDIwgEDDGEmuCxbvBYYTFuf5e7Oc8Fh9zg/sxMOR83EfxN4YF8gXZwX5IDh9E3LsawTDsSRbWPAMEiR+Ski9PTnA/nsn/7l1SQQqBCWSGJ0M4luM+qeHsVTfz9EWXnb6id3DMDU9VbuV3OQ61BWoYngWyiIHsY3qHs1JZ/LdcwJbdicDUiOiJix0xk1zGkoDZynL31BxlRVPevRNN/2aWqojGYEaBuPdLNdHTFNFxnhfdMArTWBFFNZeeeMstWWe7Ij1eiFrBcn/kStkWi1lNip7WWZv5vDurym566kqEXl6H0Qi9hAzrkgIEfUkrxEUEikBfJ8zMVv1hLjWO67FPKmxFoBAXdZLn8r2vK0xcR1WTbw7fOr6Ru2rZRFaIBw3V56jTRpLsFY7Mui/lOmvo1NasD/KOGqCVoC76MkqP5YZuvdVI6MtsnLu0Xn72g4e2JXG8q172tYf1ZAX9RlTBn1D6y9r9iWsEhaInpQ2pEBSXehpeTU7VZLufc1k/WSuLdKU1lze7iwNiVhQ6ZKgr0i/0fdChKuCyys9vKFTEA63ZKmmtuouDq/GR1ux4eTxofEYupJjMskfEBHWX81U5Q/qrBN7ulHl2SUzFcblu0qSf4G0F4lbdlpiiGoVqCSQMGsZpGbdns1hRKy50FsN/J9okbXTWvuPK2Xh+5WRz4hLKiayos6ELEz0rkwNE0kwXFFkP6Yq/HMYJxMa/UJ7WLJ7FLqwt9siGgCFgCLxLBIyweJfA2WmGgCFgCOwWBGToJkA1gZ8xoGOYP+WWfvio2/dX7nFNCQ6KlcsuWpxxyVzuGofGmsWFkd3HkkCR4N0/bY5JAZnA4t0tMWBnoIaSAddMbPMbaggWPzjEGMK2Ty9qG/LAqyG4r3ezxLkoDPgNlQbX3Bxjws/yYk0+ITR8HrkOKgtPpJzRNnlEzUEeIDk4BjdWJ5WIIeFdUnG9zYoOT1ZMgvlOk8+//9vP6mYNweLjcXgliL+eP56/uy5qZq55f+XG56+4pb/4iBu+8nU3eMFjhr8JH8Sbd/eM3uU3RFr8vrZt2cUI7KDZz/JcE8Sa8d0cjspABlTZCoN0MC7mNRt8QS5u0qwsOrKhtDqdZE0++Jsy6YizCLONQTYQsbERywXOaFzMSYlxQZVvToTFusiPgayOmVxOEcfCSItdXFd28qPTDqCGkCExl3LialVV40Yar8pIOlMWZbvApczEDZTi/YZ8u3BupD/kP0rHKraFvNzkwUycBANtN+qq5nvJt9KT9TsOvpu43vP9E8m1wqYwXJDhd0HG2iXZcw+I2alEnA4UH2dfmVcHojQ+WSguyHiQD/rD/NTivLss0rSS+6jsN/7olezBY3ssfs7WLjm8b/qn9Bnps31WibhmH9fHRc7VVG0Urb4qU5EWrYnSIpIxX8RBXWRRkA2rbntuoPgV+jzlyUbgsjXJnPoy+6Oe9W4bW2Hs9qVx/Rfox0mBMZo72D/WX+3lV8/NHFWcC1xPTZdgXBXjNbmgSvR9G6mWTuK36c/DqrIcQ1+VfTeNazE5LKjXwkgyoEbxOdXgTpwWi4tHrozbc8Oof6XdFj95rw77dwv3jI7vfWC8cfJLyezyqWhmuCZBR0kDodB1jcZEdcHzv77U9bwozb8fREkpIuefar/vo27tt2y5MwQMAUPAELjrCBhhcddfgWXAEDAEDIGti4AM3I8pd7gi+roSJMOTrveBR9zcRzM3OotwPHUtiRrqYiTy4qv6HYn6iekToV6A4GBQhzHfu2Qi/gUGdP5mVOPJBk5DrcCMRPZ7109ePcHvXrnAfXDLxMAHIoG/cQnlA1WjUsDoj8Ef/7kfVYJcuN7Fix94MkOOvPqYE+znfFQUDPSOKUEAgAEDVe6NCoN785wcj6EGRYnXxvugrp6c2Jx/7yfYkyuTQK9KEDZse9dRPv4G5/rr+hgY7OtqKt2am/u4MNK7QPHy6t8lMLj3JQwRA4HEu4G8+bDe6TmRFt/gZFsMgW2OgGykdan/1htpmFV11CnkNUNailK1ZSD7Saba1I5Duegv65ZilWpCaK2wwGWuGeHqA9dLMs6KrBCFIVpRM547jTRq6C/UVLQpZljZ5gXEsv/tEcAVnIzwYxF9kNsnVXVekKe0nupVHtTB7JQhz1VvIC7kHqrSzOtAs79lJHXVSLPHk1re7eVTv6v61tNXjG/W25rNvcPeTSCXdO1EMT2UDgq/ByeKFakbNWl9LgriK8Kwo8ZqTi7sumKJFHOnPCEj72XF3IFsTZqNeHlxrr22uj4KjCzdeqUD10XT4Nr0CVEL0z/GLSn9y5+WusGlbc3dmbiC0idIPsEgL+K0WYhUV39QtIMKxOBqK5Q6QkS7uyIFQymSIE3b+XLazuhL0s/EjRP9Wfqx1KWL6vxxz4ca7fGB7mL/iFgOl49jKRqQRAQNBfVe1IaurxhNKKEIyC16cdr/+0Otb+gOSmeQq680OuNGo533db0LSSv7RqOTPSaXUL0kzZO4me+X2iNpzYxP7D++9rgcREn5UaaNbrBc/Mv0ybTVCRXbwo37Q1cW2bXZRHq4ifpiuqjd2Fu5/K8mSfuPP/r9P3/uj3/nH5qSaOsVccuRIWAIGAJbDgEjLLbcK7EMGQKGgCGwpRD4gHID4QB5cL+LZ9fd7HcuudaDCq69T96tF6R978kwOIthHwM9Rn6M+BAAJ6aDpU9pjaEf4x8DMgZ6fqYXhnUWH1jbz8zkOhAV/M692e/JDR+nAnUFCwO5jygxi4x4DdwfIz154hzvDsob/P09Nq+CUUjRAAAgAElEQVS5DioMT6JwLRJ5Jm+sca2E6gKigkGlV0VwfYgGH6fCx6bYrKjwz3v9zFP2o8Dwx3Itvs08I8/tCRq/Jp/+OTAMQV6g9ui7zlMN1zyiPGaX3Kv/FYQK7w0MIWIga4jFATa8UyMsQNKW7Y5APR4XuYysmaQWLfmt6BdlPR5lZSgDoCaDK1VM+5Q7jMCN5bcmlAuoXAG6uxP3NdpXF9XlzBV9GWx1YLKm2eMXdG5fbnF8YOY7gpEMlN/uPr7Oc8z1pOvkPPNxf0de0069icRG9YbqwEiV5qpcvFxSCAbcrGUysEYqcXJUH0q+JEuoBEqyRGYKZD/AHCrmL1Y07vmqDl7Vn3y3dqMiKZBrJ8iJtoicroiLGYX6ONZqpgMptpKNUTYnu3VTNGo7y6sl6VKaaSMG80JxLNYhUa9ujIKZduO1mU7jFbVnQ8W52FCbkKle37C+79SCuJWfa0pWMKmFvtVDSt+vdEjpB1Ey4PZI5IRLmlJUyB3UxGhfVWsiFFQnAtRHk4V4D9kgaV85M3e0GMevduYHF/SSZ6O0uBjFk8DVfHt8P1bfrXCtzKNo3E/PZYP0oLazupyQERP3UVIvbOg+me4vZU+Au1X/neAY+on0jzdPdJkILyZkRVBvaH1Cfw5EmDTm9q9dTVr5C8O1ZiilRVMERjzuN6ScyM+IZCEmy6G0VZzVt3O5u1jfd+9T2R+O++Wx019tP7B2Qb6titjlQzmQKiqRF1KZTJQmr7uI+qQw+XGd+4+EZd9cQ23l0m55MwQMAUNgayBghMXWeA+WC0PAEDAEthwCmomPxJ1ZXg8rMdu45eY+oRCSDys8576R3BHNuuz8OZcsXnVxGyMFgycM7sw4+5+UsMB9TOkzShAVGOb5fbM7JJ57swKBbT/g2uwGieO8yyXIDGaeYYSHOMCw/zklgmdDYtw7zQtqh2eVfmi672YDf08m+BlfDOzIOyQFv7GN8oP8ExuCPJI31vwNOcJxflS2OeC2d0Hl93niYfN+no2FASrPCH4QPhAuxOQgX1yfZ/ZxOHyevXuqrkvSNRcI5v0/c4+7+FuZ638TUoL35wkbrglmMe9WKosv+Bvb2hDYjghgzJNRr9KM5HSclXsVE/jwaFz2pKgQaVGoXQiG8sF/WU74E/mJj7O8VODSeqDaVCVJJK8sUmfI97eMrk6BL0RgEKZbc5/f3EbdLXg2ExW+ndxsEDZj5t16Mzvwvir7A1WFdX3ZXiqrsjkl7uokCUs5x+/L3QwMxaIM7bKWyiWU+gXa09dxmZQWV1WX+B5PvnHEdNhBrudef9t6pje9eZ51OCqChdmWmpVI3uWCbhagtpTxOQhnhdE+ERhMHFAk7iDVpPi2SIogieLHA808FzlxPk1C8JvRtsjV4IzcQ0H+FLRvRlrc/co2JSvoe9KHIkYbRMUHlVQgpHIQjxclCo1UFRNlBWSFln6Zj1+YOCGMQrl7ClDOThZIi3wUu6vnZrOLL+/5ldkDa39JREQi9UQhd0+5iISvi0iQKifIBquto6vne/s3lruFiI60f7ndGm0ofoQKEouu3+X+37o2Cgs3EHlB39j3PekHvn6QvDOJhCicyJIVqSvqZm98bgH3T7PDD+t+T51/YelS0izGnYXBsTgsN4YbzcWyjFrzB1YrnXtU+WuKn5nf+0A5FmFyeuGeYvnklxtPj/stt3E5dQoMLrJi0vd8/Z7KY0MxLB6rxuV3aD8x7pjoY4shYAgYAoaAIXBTBIywsMJhCBgChoAh8CYEZNBmoPMTSrhuYpB1LTD1wZ990DUPdF12Zd0lMo63Focumkwc8+6S/kzbyNmJ9cCsrv98er43rHmjmzfEecM7az+42ewuySsSvAJjc2wICBJ+5zyM/VyDIISeGIFw+PemefP+e/2zbjb0+Tx5EoHzuDb3IqG84B4QKSgWyAsP7dUYPtC2D5rt1RLcyz/L9c/PgJLz/HNxb54BFQTbXt0BecF1yT/398G3N1/Pu7+aUdTDDZce7rhHf+0B97UfWXfjs15hwjH4R+Y5wOgn9I6/KtKCe9piCGxnBGp5dBrXdbGC323NdA5l/Oskg+ihrCxjuVspZFCdVcyKrmaMVzpGsXCjAZZFGRFpQLI4DC/LGHtGhljVl5q6Tz30ROEdwea3/83zrxO3x48uOrmGmbiUk5uYWkHFN8fe8T7OOb6wGBt35PXs9JtMVIQi8M5LYdSsFfxFhastNzaqItViVAeFTLLdMi+aE0JDx0jJpH3uPMoM/X1WH6TTEzLwWwrAnY7Z688322uGAgq2Qi7l4jnFz9HM9CIYZvVR4YPrueY4r9WPqHIdwze3K8BnY81uH5eVzNaunyTxOdzRZXnQa8opHW5+NvUDjJi8Q6VJxMSN7kRby/uAqNAEmOD7xWo/I6ZAxMLEJZML4lSqipZcQvUm5IWWDZEWZ+Ueqqtf1f8KcDPoY6W9fg+5Vzp05tn9D62cnn81beVzhx479/Wkmb8qhcNSnJRfTjvZ8Nxz+/661BV7B1fbPcXAUNkSGVBu5rLfmGVlR9+xwE+AYQKOdznqyYNc96hETkTdPRsjkRZzC4ev7te+/cReoWe7cOTqE6P1xlG5r+rKHdTcaNCA3KA/elGKj24UlhOXqFHkGmXtpAypw96evDl3ML9/fqgy3E7ca19vRHLTqNAY+s5C4CgCuWLj/KzYGvqi/1hY/3NwktLC3EPdofJttzEEDAFDYLshYITFdntjll9DwBAwBO4MAj+m2xBIGsP8C0qH3YGfOyT3T5ox2Ahc99HS1WXukoOxIgn+a/3O6Ol9Sq9Ot39bax84e7PRfrOawpMVm1UH3p0ST7l5dpYPtu2fHkKFfQygiK/BvbwSgmvgvgmjv3cf5e/lCZDrR3veIIArJQZ6kBQY+SFrIClIfDO5p5fWX5niw70hBhjQbnbddLNn4RneIM+fPhT5RSmCcRJSAZIIlQXbzOxjNhqKjuufhbxey18Y632VA9c+3nGP/I+R+8oPcKx3OcXzvKYENpAfvOP/bXpvWxkCWxqBb+Myqe6209FwnF9SzWhEQdhWsNIvy9XKaLCeH5R7lX2qAAtyTCE7SR1pirOTYTDHVUtW4/apGruwll22Toaa3SwfLucU02JNJMgtJSxuEqwXzCdtkQiKSLOrEwUAxxQVrg8yeZTRfOygDBupAm5E8t9xrX0hX9R36vWEvBA2gc3C3tLFd6tnzpPvq6oHL8poOZDJfEMz/q9qbni3LOqDZVA+qoMUwaJeUz3St6/Wd7Je1jF8+1a0z8/k5jtW7UR1xc1e4t7FTjAYMinepUVRHiQkjurrBu7p5Iau0W2lkKbj4Vhz1EM3EikUCUcZgt1GndfrMgjPjMbZbFakihkywZEQBSeKomqrvaJ+51a/71oVon1G+co6l+UdXcMzuH+S66ckjBRgW/Eq+DVOGlJZNM6FUdISibEmpQXn0S8koTKeuHC6bumKAPhLw9XmS0r1+nKHYz4slcVDim3RDMLqtOpjlA2TVMctSFVxo2tMLzlRDyqIxITsos/o3ZRClLBM+rkqqIWiztCfPSFVx5nuwiDWdQ8O16RDbORy/FTe09uzMaPjussnF9bltkpuy8K18Ub6pwr4PZrZt/5oM6726Xf5vXJRlLj3t+fq/sFHy0zen06P+9IN5W5x7WJ44PKZVEMF4llM5/FopU3U2yeVvqh0buoeykiLu1bE7caGgCFgCGxdBIyw2LrvxnJmCBgChsBdQUAz7xlkEUQQl0LMhHqfax0L3N6/cFAjs8pFPUUS1Hgoml8TWfGcfscVEwTF7yh9VukHlZDLM8DbPDPYkwLXKygmYyglv5+BC+f5c/1vHOeN9fyG0Q5CgQGcD37Nfn8814OwYFac37c5T5vVHezHZQNGfWaJ4noJoz4DPsgFruHzAzHCPj8YZNsTA9c/y/UuoG70LJ5EATOw/LISbqZ4PvLPtxoiiNgTBCT3Po79N5x8kQeuk+mdyFdA57Trve+I2/MDy275t/kNgofzIJVOKaGA+aje9f8hlYUFFuat2bJdEZgY8mUULLOiXC+L6sK4rNNUjln0X0M1c6/8ysvVTRVhQEyTaE3xLkYiMjDGaupnuKYJoKM4CQeaHT0WkRGIKJi4XbqVRsKbuZKh3s52m9FglLeVt7Y8V4XKZ7OpTAauznO5sVrvj+skVmRWqUJkDB0pi5AVEwWGjJm0E44gveBws5doMS62a/G+/fmGXBCh5pWKCqJdX5FRvaPyN6940Hw3cJ2mGeP6xigYtyyefANxE3kOhZIqIGQ63yxiVe06w6PamgAHWRJwMbe+sTDTnl8fjPuKXVFKvTUMI83yqMOw2RD9WJbzZV71dEpT2OaC9EAuScbqRr7ebecXhS3kTy7Tsay+tQJ5b+5C3f6yYHd4EwL0s/Ypoab4sN7Pp4lR0ejOqquVKBzJeOIKCnt8lKa5vjq9MIq62kGd8Crgay5Vr/XTIBOuXy7LRdQr2vmUCIRnaNc1HWhOte3T0+N1vYkrqrdYJGNQZDkdRN/Ux1/zBcjHWiMvh/TNq+WGKhQJEik2hYgGderrYB8upyBGRJDkIiraipmR63e5Wq0Dua/6XgXmHvWWNs5ei+c96Y+yoZKth2vVq1HhnlUMi8/1V4J+ay7/L+vT9YGKwOA0HRw6OU1Ex7W+KG5K6XMHIi1MafFWr9d+NwQMAUNgFyJghMUufOn2yIaAIWAIvAUCf0+/M5Of+AkMSJbdnh854qJOpkFY7AYvnHMzTz+v0Rq/YyRnoIXa4IeVUGUw499LzzcrGTYTEN5tEmv/LdqsuNgciPp64oPsXzPOXyMXiNOA0oKZnqgS/LUxtDAg8n97V1GeRGC/j6lB3paVTihBgpxVQtng3TZxT58/fveznSEUeHYGidyfge3mGBbMNvWExmayxT+DJ3E8YYLMHtJisyso7vGYEoM88uuVHxiHvKsr7kk+rg2Qo0TT2vYWbuF7IhEW5IFn41jw4r3xDGzzrn+ezNhiCGxjBKpWM8nWVsZXRTiEMvp3giSYi5O4PxxlZ+RT/ko2LtuZpiznuf7lxT4dVuqcNRkFr2ra+NlmM3kpCcNVucHJRBBUvU7D183bDUs4HCv2bhL2qsrNabZ1R66r5tXWVmv9nNgAsz3XXBJ/cUWztwl2uq6Ax7QpEBW0CbRrPtixJz9vd57t+jsMgetIi4bqRSYjJIo8vjMQFHxfqBNNV8ltmoLuyrB+Rp+bXOuL0+Moh7tuabcS10yTVHE/2msbWVdqrwcUL6erOBXdvCrS4ajuimhMRTRmmvMhlaqIyErxifM8lnqlFYksbQZVV+3QmdqFa4Oi6GVZ2UbpMs4KNQBNq9d3oFTdwB0U/Sra2CeVLsnV00/HzfZ3tWYWJ8G1A/lDSpptV4zlGTVplOp25VJeXIvBFgT36n8m0tDPoo1mcg+BuiEu6JduXni/X1KClPDuSGdU2+iH09+jH/52Fvp61FWuQd4nrt6m90cpTd/8JZEjeT5K94iU2Jjdt/6yXD/Rb31apEuX2Br9K22XNvPT2Shp6pjFMos+KrJGapJ6OYiql9K2Su+1Pjh9bJ6NZ7qq8npWgpO60a1Hx54qDktp8Y0qc2fOfDP+cJm/4XNK3oj/QRy1X1b6l0qfE/6Qnm8iPOUy6u08ux1jCBgChoAhsAMRMMJiB75UeyRDwBAwBN4tAppxf1TnYqBgkPMVpQ+5eU3y6n1w0YXpZVestVw8vyzygsHYn08HFxi/f3o6gPmQ1te7RvKDbU9e+LgNnqzwAypPaFz/bdo80uFcDHUylEyM7qgiHldiwOUDfuJ/ngEbkni2WXMNBnPetZQnMYCK+zIbjusdU4J4+P/Ze9NYy7Lrvm+f4c73ze/VPPfIbjZb3ZxEkRRJUwo12JKnmFZsSU7sL0YSBIaNAAEyfPUHB0aABEYCKAkMWYrgSLEhmTZlSi2KlEmTzSbZ7G42e6x5evXGO98z5f+7dVf1qceqriLVXdX1ah/Urnvfuefss/c601rrv/5rMQYMT2M4MHYMKX7D8c8YMNL4znwBBDBC+eR4HMdqYHAMW3Y6QW0c9E+DyYFxSu0Q5sY8KSROGieMTQMomBfjM5lxzjgefTC2RUWOn3VLf2neLfzr027jTyk+/ik1jGbmBIvjMbUe51wsC+j5fvESeM9K4BYMAYpvK1+NUrCERUcRzPlolK0qsvn7uvVXiyx4TOyLeDTOZ+UUXK/G8cmWqlwIv1CmFkWJq37FcJisplG0rlU9pXPJ3m3AQhHtExaZWB1V1amIxZ5YkFPoRKI0MJTaUCHwSMDFov7eV6+moldEb4xy19ffSsRRCJOJeuJg2LOaZ1uZMfaePY9+YO9pCXAN8T7mfSgggndmQVpIgPQmmfq1wYoAigP6vqXf9b4ruAZ57+FY5f14X6WD4myqxowToOgGw2Rbz5g1CBe6N/UYkQs3dw3lz2xSlEKApAoqBx1RVIe6t6u6hwtlfFLap8g164rMD6NGtRouCOyY0/YjsSwSEa44J0PSQk3v8esuIM+ceufup7JjfFpkG2CYZ+tDAiD+oUCJT9VnFpR5szJp1KooCopX158N4+oDAqXEPrqa9kn3hrFpJ/eE2ptqsGj5ju7IeeU+O6CGvkcgyUm1R9XQJQm+YVtj+d5qouin6IXo7fR7TM3SgHJc1r1PDRZ0qFoYbvXNpf2d1fajYlJEc/u2xbSInNJCOQEUYpCMzg27tcPJQLEvxWQc61ESvdmYHX47ijPmiL4MIIOui87LujnCZWqt4perjWI7S4JTT/5S8s1hL/g/L78e/X39TnDRzuW/mo6Z54iBLHcqWOBWMvW/ewl4CXgJeAncZQl4wOIunwB/eC8BLwEvgfeYBH5F48ERTs7b3qQmQv3IPmUmkZM7mHeNE7JkjisIMCKlEAYKTnScGRhYN4oaK9evsMgpS/dkxWONjYEozFDZ+Wlgh6U/wojDoY9xh0FpkXA44zH0jJVhTjwDBDCKLDKMdyAGHg4aokcZH+ADvzMnS5VE/wYOMGco9WZMGoDC70SHlZkjGHPlYt/2WznHg42LuQNUMH4MXJMRkX1E5SEjolgBlFgwFidU+ukxrCA4Y8bI7rooXnL1Y4nb97f3uK2vP+ryMdvDgKF/+uEc42jinP/jab/+w0vgnpQA6Zvk1MsvrHa6pE0Sm2LQqlY347CyR77Cfn+ULOqmmms2a0oJFZyVszDSzdMUANBVFPNJrduQ43BbXsbkF54+eKfS2lQoriunZENPjr2K0H5czuAZFegNtrYHa0EULqlk+AGNb1PjPCgH6AIFuLV9V8MntRv1eyzVCPf+0Dsw78nL9z0x6BLLgvca7wsWoqgBwZeE7vEe4p2xqeuUdyfb8Ykz1MCzO3XvvCdkRv0YBiKW1FDpn7YVYX5Bed3OFEHQ63SKfYWgRn1PlNopVHo33cJhWlE6KAAO1bNIBkkWxnGQN2rRuthUiYCKQateGyt4P9dzrK7nEfK/L5krd/kEm66JjvthtU/BqohVWFsAhXJ/Wa4u3RJR5VEX5NvV9ujrcbX4lNIqLaWjCbF2KMYCeiHXiNWwILCGZzVpRwErWNCd0cd4nhMMxDlH72RB17ydhfES8EIaV3RbjoOOzEDQD5nDNd1TNSvcuFcTOyRWUqg8UdHvTN9nlZJqcqz+VoMgFti+6K3/Vimg6gIqUqWLol/0WubEvc8CqAloASBCcfFMyalGUbU4Obe3CD/+66P+v/ufG//TYDv4vWsa/vUz+ln9+cdq6Kb0ybPnGmgB88WzLK4XmP/LS8BLwEvgfpGAByzulzPt5+kl4CXgJXALCSjSnih+mAoGMhxzNdWuWP75Pa66d+jCSkMBli/IODM2weFplxgqGCwWUWbOdgwOi5iy3OqW6oldjXnBNhgqVoehHF2F86P8rjKKuyKn3UfUMPzYH6edsQzKrAXGZrUsOAaGP8YgxzKHC4X/ACowTF9Xg5ZvLBFjZ9hcLO0UfWJQMjaMTRw6GHKWeokxsa/Ni20NEGHu5aUM6hjwwn6Mh/FybM4Lf2P8MlcWjNCJk3J6HP5GBoAqzDHXOUvdzEcvuvnPHHDrX4StAShCuqljanZu9nLuxbIgZYBfvATuWQlMa05kYi/kTz92oGhUK9lYmbgFRqwpVVQjqMXLYjLkStmyrShmQqCTSiXqKt/82kyzlijl0ugXPnb0pnUg3gXB1HTM5cE4qCsdVU3OylAOrr3KL35Qd+eaUu9QTGNlNM6OqNzGlWajKoZF1u323Utp5tZUPDxVs7QcPFsTalm8k7U33oU5+y7fwxKYghaMkHcP72hSzLDwrjEnpQUC8E4zkH2Slmw3F9uGxXWTpaD2jap9VKMgXO8Nx28mmcCdILisIsSZ0jvVBPBUAxeqqLZrj7JcJIxApWrk5taNnORRPEyzvfozEfDx0ly7NlYM/1BgZkehCrzf/T19B+8ZOci5ztFpcdh/XOfxbwIwCVkiBVShYtrloBMxLYK2MkK9NrvSXyfNUq05Xty8OEvRhrb+03l0Iz3ZLwsk+IHqOahm0qQuDIBFeUFvs3WA0aSDMh37ZrM3x77VcwNIIMAFPREQEQCjXH/tun7EnCgEUHxBjQAW9EKKYbM9C8FABOesaexfqTaSxw4+fuHi4iFlfgoLdFB0ZJsHnyyMH6DjB2o/oXkf1hOjoYLcS499NvnKq38W/y/9jfC/UX2OSc2P6XJSn8fU/okaOupvqZEeywCb68bs//AS8BLwEvASuL8k4AGL++t8+9l6CXgJeAm8nQQ+qR8xPIjqnxTadPt/bY/SP+UuHyayMM655hM4LYiiMlo7DnJz2GMsmSGHw73MnLC6DhzfQAg+bRur82CMAzNn+N3y5VrUJ8YYznuMNcaJYWl5dPm0tE9WRJRjsw9gAqwHjkU6JBwsGGREtkHJp8g4HokLakS5GTDAviyWDsqAiomDcNq3Of8BKfid4xgwAjOC8V4FEa46fYwxQr8G3Fi9C9ZhvJpRaNsz7p2sFI5jYAq/w7xgTKwHwHjTNR9tuv2/uiXAAnkAqjAOa+QR/q4a594DFlfPs1/ucQlMnabjLzx3Lruy0RsoBzz3RkvgxDppWES/CAQUOHkNR616ZdiozfIsyMSsuJNgBfe18ooEbZcH+/TU2q/04Splobq8eV4dJ/kJgSuZalpMiu/mebbY6wfNcRz2XDGqN5vVI0txIy6KsC/HJpG0PA95PnPv31dR7vf45fqeGL5AvvI4ykEDXFOA+7wbywEIOCx5Z/E72+9qsOJtTtJk7mJQUPNje7Zdj/vDcaeSu6bqVYxVZFsFit1BMSsq8g9r20BZ/rWocLmKWhSuVslU4LwjPoVWuooAjJbu5w1915NrvFmtNCbynTI5fihVjmdUvbO3zxSswD+C4//vqj2pVF2u2pwRWNESOBGWdberB1cB6rwIR1ElKw4/uHqpMTfIh536hXMv7esWWfiy0i01GnPD09211sWNs3MtpV16SMBFLuCC5zZ6Ho2AIUAKdD/O81Ud/Or3G/lrYDKgu7GdpZpiW/RSmBpcN5+dSof7l3vVwIh/oe+8Eyl8/Wm1r6mho07SWYlN0ZVW+rwu0lEU5eutxV7t6FNnz+x54EpbbAz0fXRadEn6gDkCe4PF9HzeRQTZwFRek/hGD/5UWl0+ml9+/T/Gf3juhegjw24wL2CehW2oF/dRNeTxr9VglaCv+9RQU8H6Dy8BLwEvgftVAh6wuF/PvJ+3l4CXgJdASQKKsP+U/vyQmtV5GLj64Yac3UuyXuQgG2+qjsWqstNiGE2MGi04xo3SDlhhtR8wmAyAMAeHpSrCyLF3z3VRatM+zaFvoysDHTjUMYKM1YCBZXUbcDhaAVr2pR/G84za59QAHUj7xDoAFyLYMN4sSozfjk37A6xgO6PlcwyAGcAIPg2kYc4YZgADzMsKeF+cHh8j0frAyDOZMD5jXpRTVplcmAvb2t8GUnCMct0K+rFUVIA2ZtjisGSsjOchF1WfdfMfe9XF2jTtcm6YHxF5ln+Y/j+ka+A1sSy+TKd+8RLYDRKYpnbKfucrb2RL8/L1k5BFgdDyFBVXhvIvCoZVmpt8/8pMfhdYCRMmmNCJ6qhIVAS8Wmk2ojVFWStBTKii2/msy/JABXlVoVcFfJUbvBE7OTOLo6rQXdVcKMrakOMrFahxUU5OgFaeHdzbfvES+PNKwJyFfFp6RN7HBrBzraUCBz04Ng0koIZBo14RgOhOCYQ4Lte2XNhOpXHCGa2riVKxVovDem9YoBcoNV0Y1JUcyhXBumrrnK5Vq51qs9KPw6BfFVej3axaDQUv4z/v1fyj7891j95YUX2KK3GtsVypN5QNNRdoIehJKZVo3A2VekKRanfsg2cW24u9A6BRs3s7D7WXes8Nthrfmdu/9ekozj+qZ3V/uF0/+8Y3j652rrQeH3Xri3l2Df84pmOtqgEGWLpPdDOCaW60oL/CSADsoDYE+ijXFcwKC5bhvuV3dFL0RwMs/pa+/19qRzSXpt4fT2lew7iWnqEujYprr7UW+8/maXh+8dDG3P5HL89UG+OatkXPBFSBjQG4YMyM39Z3amMwGWwC6sqxHduz7Ter9aK9fDw73Jgr+kuH82de+Wr885vnw7qOZ/YEc0RP/odq/4/av1JDDncyiIAx+MVLwEvAS8BL4D0kAQ9YvIdOhh+Kl4CXgJfAXZTAX9WxMXjIf4vRdMy1Hs0ntSvixa6L5ysumuedgXGBQQRwgbMfow5DCAc5RpKxATCwDawADKBAN0YVjAYMMEsNRZ+WEmnnvuYYMRDjhLaFbs7xjI1AZJY5UeyYiNH2AYghUstSV2BkYbzhtH9eDaMKpz/9wbDACQMoQuokjg+wYGmn+I5TkPFDfWcfPnEQMn++Y2hhsGGo0Yh0I4KM8UwiMUTPtgYAACAASURBVKf94ohgsbmX2SacBwNIzGnEHC3yzuTC/oyB47A/fSFX5oOhh6wY635XPXrOzXz4vNt4BtkxHrZnv5NqpD2gJgnXgAcspifGf+weCXz+kycmoJ/lm1dBbffLHzly16I3Fc1uz7rJ80CgSUXJwffkRSUTIKFnSdEKo2hRN2mUjXMitLuKRl0YDRNFZEekipkfp3lbRXxPzc64rUY1LlSRg2fB5BnMPO8CALN7Lpj7cCYCHm4062ugxZSBUQ4omDjRjZlxk/3vF0kip4k8VF+mkl9lS7yu8jSBUs+leSWsp0rvViGmXiurlXxJIIarVMNUb+1IKzqqU4NjV2ne4tUkU+HuPCSg4Nq73t/P7/6lNGVXoENxLtEHJ/qmnr8P5elYsR+hq7dHrjk/cL2NpsvS0LUW+q4+Mzo9s9IdCqD4kJ7fhwRloCfO6++P6fdzWqfAH/cI1S7ipd7TR586466cXOpefGVPZdipqbi9WHZX9Vj0YXRkgAXutbcDn9EH0d24TtBXTadE50OHf07tmBo6MmwRdErmRMpT5viQGCGrmk8o9scby8fWnhOY0oyqWW3hwFaqK3UpqqYvziz35gRmEMxEAA5gyuNq6JDo0gAMgCYwe9GdGQu/s560rVy/HOuCvv2EmBYz7aW8s/KAW6s2i9/4+m9VfzIZBR/U7+Xl5/UHQBGpWl/d8Zv/00vAS8BLwEvgPpOAByzusxPup+sl4CXgJbBTAoqsf0rrMNAAITCcMDJarvWB0MVNpVKuL6qGxapCy6xGAimUACvMQOITY6sMGGC8sA4H+Fm1Y2r/Vo0URDjkMWIsR62FmFkklQEdBkRYEWqOg5Od/f+d2qfVOE45FZWljcK4Msc9hhr5LgBaADAwqog6w7kHYEH/GIasM9YFjn3myJz4nYYBhmEIGABl3dgdljrKioDjvKAWxhtqGIvMz+j9MDuISivPEUcFf0OtNweF1d4w2ZSZGNrsupRS/G2gEd/pCwOStFeMf0Pn7lG379deEmBB3Q9LTcUxYKnwybnf4FoQy+LbdOIXL4HdJoH3itNvWieAe1rsiKAvtsSqPJzHB8PxHqWtCpXfPgmFY8hRJiAjn1Ex8L7YFmF/nFbGaTYv6HMuUZoo7aM0IsE3ilbhVIy7UF/c++Zwu2uAzG67bvx8nCsBEvftdfU26ZdI2WTpIXOlndsj4paAxTAROFrTPbyepsVrAiV0d7t51WseilXRaVbj1CkF3Ey7ejoZ5SrUna/zPFB146EADXQZS7d138r8Dt97PD/R5wg++U/V/nv+LorMVZqhm1nZFmAhQozobjMrHZcMK27/o5c6M0u95+X0f0XAxMem4zVWREWshL+odejBgAgt/b1ndqU7GnVr51XY+oCKWBfjftVqOqB/flqNcw+4gO7KOvS5Gy0PaeXLvEfUTB9nDgAZtPKCPoue+5LaYYDx+f3bv610VTMzy909c/s67xOjIqo0kgUBGcgA/fWytkMHRedH5/369JPrkkYwkjE3SFEFoMFYGQ9ABjoydThI94Tevak3VDqzkl8c94KkNuMyhUTtBCwYMzoxeiqgzHUFuHfMyf/pJeAl4CXgJbDLJeABi11+gv30vAS8BLwEbkMCvzQ1Qqz2AYbFBbErqi5emXPxwsCFbYwhnPs4tzFmjCFhjncOw3dL4YShcXJqdGC8QRmHJs5iTnhLCWV/W70Kq39hRjrreV9ZBDHfP6Nmjn/rx9JOMcZJTvrpeMi9bTmBGTsgAgYhbBL6smLYAB+TNBfTcRtgQrQY6zEOkQMMDfYxA3E6rUlUGZFsGHoYixhdGHE/o4axCjhAZJrJyEAIQBjADvu7zKqgb/vbwAwi8ABOWI8RygI4YwvrDUBin2OTMe39a3X3/f8cVgkMEFgnlu+eba2YONeCByxKwvRfvQTeRQmIURFsqa0LnCCqdK+YEpR3VaqqfKi8T0V/lGejNJdvM2wKoVCK+6KuLXpKhE/l17q2XxHTYkFO0XPVMLLUeNzPfvES8BK4QxIQmAGDi3dvT6CD3vdRT8nnklazelBFKi7mmQtHtWy5WguXVJCmOlauqCILTssZnqkEwnYUByeFQQqwELcqDAb6D2c193PxXgFa75Ao7+Zh0IXQc6np9Q/UGkDAldp4wqRYOrLl8mxusHlusTF/cDOvt8cdsSuUxmt8QiwEdC0c9uiX5UXgVfCBLAl/U2mhTgiw+AthnM+reHUnz8NEOy1cObXg0vF1Lhl0M1KgAjBwHfz0TYSCHgu4YjrwzWR3Uj8AOKDzUp/iBY3j9cXDGy+tHF87rFRQTaW0ekzrU7FDTunTdG7ABPRTjoEej36I3nt+0s9V/dN0SXRSdEtADPRsZMh7iEAhJsf7DTCjEVfcQ4354isrx7Nxdy0+JU0WXb68/Nf6g2v/i2pfVfNpDm92Zv16LwEvAS+BXS4BD1js8hPsp+cl4CXgJfB2ElBEPcACxg7pmr41NTbmXO3Qabf8l/+iS64oArB+XvUsiHYiVRJO/XK6J7o38MJSHuGox+kPnfsZNSLEfkvtH03X2/YGVNBHuc8yEECfvKsMjLC0SIyj/BvjwziyXM/0wTYcm9+g6AMiWNSWUdXNsceYYIKwDd8xEjmWgQRWyBsjCqOM8VgKLKtdYXUprBApYMWnp+PEqMNgNOZE2cDkGBjJZdaF9VlmWBhwATDC+Fjoj4XtygwV1jF+SxW17KIZjsE5QZ4YoIAXRL9xvugP4/Q014RYFkTN+cVLwEvg3ZVApuLfmcJrKdrbkYMzk2MzqNbc5SQtFtIsnxHbohgmab9Wia7EFSXpEGKhuhcDbV+VI3RWhXnJj3+uVot47vhI7Hf3fPnevQTeTgKmL0wCJgQ+/EDQ4xWYUmElqNTyYBI5Pi6CWZWmqbkwP9cfFf3+KHH1arzRqMS9amUCOhI0MgYE8eK+MxKYpoPCOQ+bgHOwpPPmGrOFWz7Go7Xjao1go7mw0RXAPFw4IIypnhS15jis1MWcqWToT+iApNfEMU9wCoue7sGyQIv/LBnFcwItsjDOOkocpqAgF+iJfmxmpVfbujhT0y/olCwE2aDb/ey0r5sJgesNoMACV2623TF+EKjSqbVHv92cHb7emB9UVo6tJSoQvqF5Kn1ZQUAOrAgYGBTjZvwn1LgWSc8Ewxh9mmNyPH5Hrz2uhq7JnBkzwAT6IzKE6Qy4wb58AuY01cNJyfXbD308PXz59eh/6K0H//wGA/97WodNgi7vAYsbCMiv8hLwEvASuB8k4AGL++Es+zl6CXgJeAncXAKf1k8YWhjGGBsYHmM39+ETLjm/7WY/VneNEzjnMVQw5ljKBbUNaMCIweFuDAVo6myPk56oMwARpS+ZMAGsODd9WQ0HAAEWYx+Yo94+zZAzw4z1BjbYeCztEn1iPGFoYWkyJyvQTf+WwopPHPX0Q7QYc2SsfALO4PwzUMTYH+yDnMyAMlYEY+edyhiIFmN89AEIQrSZ0fE5FvuXUzwBrLBYHmyTBX0ge0tNZfIlYo0xmqx2yqzstKQPxsUxP+k+W3zH/VHwx/oO24Xx0b8VPURuXAufVvvCdEz+w0vAS+BdkIBS7OTK/8/zaaQCvV3VAr+ovPfHlDbmYF6EidJAJYq07lYqYZqkYSIo46IK+i6MAtfuDZNBvRqui2SR6klT13a4xdqDYbKlbXg2eUfnu3DOfJdeAm8ngSnLgk0mzAi1QOnecD7X87xQ8IcUknRSzmo7joNGtVK9Uq9WeqNEZS6U9k1ghekjHqy485caehT6G/XWWNpocaq14JaOqtBInBdz+/OkOT8MZvb0Tuun2bia7RVToSFnP455zh26HycYp39PrInVwVZ9Rv20k2G8R9tGqhlR1Nu5Sq3nvT0PXKnPH9gKti7NqNLJ4aJzuV0l3ZQWwAAAhJulgjLp8Ky/UUF2WA7o3tcWFdJ2qqmRLxzc+imxOwY67jgI81EYFMo+ODkO4ycY5q+rwfhFF0Zff1PtT9VIWfoJXdUq/iSuXxZ8ZzysfLHaSP4LrRfrL68K+OC46MjIkPptpM/69wJsnpWMHtb8ATOY10rlahHuYz/5K6Mzz/zv9UsC6vfugNsZC/U2vK+qfCL9dy8BLwEvgftMAv4lcJ+dcD9dLwEvAS+BHRL4Rf1NNBRsAGpZRG7hE6+6pV845tofrLmojcMdRoGlSyIy35ztVuQZC8tqSeD4J5rKctCy/Z+pwa4AQLhaU+Gteg0GSBijwNIwWZFqfi+DF1b008AE/sbQwsnPPHDAG/DCOvojCowaDYyN9x7jYJsySEIaJ8ZFwUCAFvYzFgVGFn+zD4ADxinHt9oVNmYbJ0YkAAnbYOSxHUYcwIC9d41NoVXX5sf42I5P+50+y8XM6ZNxMGcMUsZjv5eBivI5srRXVyn7j//zvnvx12CcYAyS3oq6FsgfkIlPrgkPWHBm/OIl8O5KgPttO44CuZPcopyaV8K4qFYrYU0gRE8Pt2Wtryr3k+rwFnOK7HXVOK4kqRKfF4FSzhR9PSAqmdJEdftjJ5BjLMCC55ZfvAS8BO6CBIwVofRQ3Ie8vyfBDXlRyDkc6BYNVbNmUrJgRn9vhXEwKFwUCrCwugCkgPKA450/d+hRBIfQ/haHJx1UTfWBZvQUrreLC/WZfF2OdulN2YPS7q7qj8FEZwKUQpfC8Y+e94d5HmxtXpilr19MBpUTQZTXxr2a66y2+/sevpxHlXxWqaFma61xocLWQ4EX4WCroboY11wz6Ge3WowpvHO768AKAQWu2hiPGrMqjVLJDvc364XSQTUEmtTTJBawUOwXIHNZwMJwkhYqKNDnvw4YM5WHpUQ9ovfOOEujme5aq37quUMrBx67+Eq9NX5Mc0kq9eQFNQJqLguoOTXq1x64/MbyzNrphUcPP3H+yN6HLh8SwAHTF0BEx3RP7nkgf2x+f/6PN86G/3QHPRAdlzRU6Lvo3P6euNXV4H/3EvAS8BLYhRLwgMUuPKl+Sl4CXgJeAm8nAaX8CZXyJ9cnBheGw8fVcOKfc/VDHXfgvzzhKouRG5592bUeJQKYaC/eF5byaSf7gb9xtLMtwAcGOrUcMMCJ0CLNktW+IC8vTAsYAizl1Ej23ewWYw4YeGFpmejXjBfGjVFo4IQBFmUGg4EVzNWADYwqQBhADsZNjQnmSYok1luhb7a3tEtlR6CxJHaOmeMC0jBvDFmMLr4bi4JxAxYwJkvjxCfbsi9jYZwAHhiJGL8AKWxDH/RHygEMSY7NJ/uwfxnY0J+TfRi/zYW+Puj2/apyGNfm3QufBxhh/tSs4HwATNHfq1wbukYyfcb6tOLo9OkXLwEvgXdWAuk4yQYKT72k/OHfC1z4hmpn75WDsxsrGX5ciZcVlb0tkELki1TPIBXkjkIBE/G6VqyPRlmtG40C/b4VxZEitcNABbgtNc07O1Lfm5eAl8DtSoB3vdXSGgmo4H2td3nAemV2y61mWCKwwnSrie4jsOOHjvE2Bb9vdzx+u5tIYJoOCh2XYBVj2LpCZ2rYDdzmhdDtfySrxNUC3RadCtYEui7nC52RfdDrXldDH81VVH0xirNPqLD2wcuvL9cy1aioNMZuuN1oNucHmWpiDAQepNrOqeh2nCWR+k9dOlJ1ottL7MdWXEPoim+7CIxwSv1UEyxeFWihwtfFfhXYfjaoFjMb5+YKFQDvzu/fWl8/u3Aqz4IrS0c2mlkanlJ9jjMCVISrFbAtPiNAY0uskQuD7fqxcy/sf3rzwtwnlcbq95aOrg81h0allpxYOrJ5UQSMzTefPbpy+c2lX1d9lkc0n84b3zj6f+vzW/sfubSgFFqkniKoqYgqxdyJj6SvfPti9ZksmdSmswVd9HNqsFX+hRqghV+8BLwEvAS8BO4zCXjA4j474X66XgJeAl4CkoClN/qr+k5O2W+qPaa27Zb/0k+5Ypy4eLbqGsdxyuPYN0c6UVtmSlkqKBOo1UrAWMOpznY4w8lvizFnqaI4tjETrJYFfeBgwzFuqaXKgEMZIGG9pYBiP2NCUIj6K2qfnvZP31YLg/EAIjAG3ns4/mE+GG0eEOXJ6UQwWJkL+9uc2IfoOQALy9PLWFlvRW7NQcgnfWBcASBwHANcjIlhYAVzKad1MgcHDBUiy0jZhFFMHwAzVoCRtAOs59wwTnIu4+Fgf45px2FKrGOcyILzASjzqs7twB3+B0+5M/8UuWBwQ9/nfHMtcE38VYEV/5L+9TkBUwRc+MVLwEvgHZSA0kLxDMiUGqo/HqercmqqmEV2MEmCIMvdfF5x/Sh0fTk3qcRblQOtolQyupeDcaBSF3J0tijYXatG20onkwVhcKP0IO/giH1XXgJeArcjgWmh7EzgwwSgUDM9hvdzpnudd3qZMUq3t+eqvp0B+G1+FAmgI6Gr/g01AkaOwq6oNgq3cjx3h55IL83uLfphPEn5hPMe3REd7I/UfkUNHYqAEBzx6G1H5NxXH8Xy9uWZ2WRYcWIkUENichWsn16IBBgsCxBIVbA7j2uJQOi8EDthPOzWqoAYt7EwTtgKt6pfMTkuRcOVjkq5nFxYqabM9YqutrBSS4+de3F/tL3aPqxx/rSAk/aVU4uXR71a/8SHT7k9D66eF9S2KGbF62J/1HrrrRV9jnqbjSdUk2Np69Lsr/e3G4dqrZET02LveFg9q/X97lrzM+r/SQEaTKWejIK/c/m1ld9rL/ZPqGD5UhgW6Kxbksfc3oey99dniu/2N4LPlMAadqRI+ER/FagUfuurv+lZFrdxYfhNvAS8BLwEdpMEPGCxm86mn4uXgJeAl8AtJAC7QpvsmTqhMQZwhmMdbbvK8kHXfn/o4nmlgprZdtEizutPYGyo4QjD4W31DgxsKDvIcKiTPgkGBZFmpBrCgONdQx7cn1TDuAKwsKj/smVmfZoTv+zQt/RTzNDSRHFs+oYpgPGDoWjMB7Yz9gPHYx/my1yMZYFzn34BBxjnienfBkawHYAE/dBgSmAkWtom5gCAYWOjPwNaWM93m5Ott0hKS0dl8+GYzAMnBv3/iRrGM8fnmBjIzI85I2djewAG2ZgAScj7a+OwcXMM1nH+kIXO89ORm32t45Z+ccWt/RvW0zcyBKxgjMgKY5hxdgRW/HDIJ736xUvAS+C2JCBQ4u22mzCrBD6MgyIokqxwee7OB0HaHuvpoiLbwyiMukoZNSu2xVDFfLeHo7SjQtxr9Xr8hsp2nxqMkhxgo9cfZ5//5Anv2Lmts+I38hJ4dyVQAi7KQQ0c1MCJyadnULy75+EWvaMXofOgCxLVfzCMXNpaKOLZldy1l4uOakBs6Yyhd31D2iR6MzoTehWBMj+tBtOB+gwZzn0BD28KsNgrECKiLgWOe4EBjkLeAgSc1juxFeL6WPnB8lBp/3J+L3QM0z9vJZDr0j7dYGP6QSecFeOhAssirqdDgRbdajMZCsSYE7Cwff7lvZlSNo01rstifBxVKqtekYUvi2Hxqe//yUPU13jt+IfOLAikSLtXWvGV04tL+tzobTS/IFDmV7X+EKyQUafmssXegi7mn+6rfLzmP2vAywSEKIIVgSKf19xPzqx0a2E9Qd6vqp2Mq+6CwPi5m6B1BNUgZ3R9n+7wVleF/91LwEvAS2CXScADFrvshPrpeAl4CXgJ3EICKP5E2eMcp/Ayn6Rs+oGr7l8QaNFVWqiaDLKqiyqf1Hqi93GaG+0ctoKlSDKHPIfEkMCpDaCBw/1pNQwq6kdwTOoi8M6hjgKOdL4bAGLOfPoxpoU59C0CcRKVqGbsELazWg/U2ZhEKk/HagW6rV+LQLMi0/wNfd9+Zywcx8YGqGG/8d0KX//BdH4/y0Cn88JY/ZiaFUc0kIXfy+muDKgwBonNxWw05IRhxj7IGoP49PQ4pGoyNge/IX+ABeTHPhillh7K+is7R5ibAS50+YhC7r7g0s297th/O+u2v/Y9l6wf03qAD1J5fUeNa8NSW3H+/eIl4CXw55CA2BRvt3chQCNRWqduqxmfE3uim7tc9124qVoWpHpS6YrwZDJOD6iExbJYFpd1g5/Uzb7V7Y23BGis94dJVyyMwfxM3YMVf47zdL/tquvOAgCKh44uBetbg3Bts2+sQDdlAd1vYnnH5zsFLujXsyjecen++B0Sua+9ASysVhm6qwAGKZhrgcCF0O19JKg3Z93Z5nxxXBoqgTfoj+yHjozTHZ2TPtAXO3Lk/6HSLO2NqumHW/ODyvqZt045znuliXIXXtkrxsPQ7Tmx5gQcuPWz806plsSAuC12xa0mjE6IXgxoMcrG0f5Bpx4pFZVYeoFT6qaejnlJ9SVal19fWRGYgu4+K5ACpjXzmATnCEB5UuyLryud1dlRv3pl1Kt+TWNsq4bF+3UVn3prEIV01aIhAGZFwEWgehlXBGIciapDpdSquVxAjYAQATPBd/ubjUsCOfYp/VVNgM6igJIrzfl89slfHF949nerX06Gwad2TO5/1N9fU3tOzQMWtzrz/ncvAS8BL4FdJgEPWOyyE+qn4yXgJeAlcAsJUMiPPLGAFjAgeA9Qv+GQaz2SucFJRWNVB671uDEP+IQCDxBh9RjMAU6kv7EXjGWAoQQ93pgPJ/WdGhlGXzf2BPtaaidzrlt6pbKj/5ozRdvbdtYHY2IfYxYAKBAhZ4CIgRzlFEnGmGB8rIcJwj6WnsHEV3YqsO3vqlGQG6CBfWA2YNQBNGC44eg3RsMknmw6XvqzOdxoLvzOtoApjA25YPSStxfAgBQEGGmcL1gWADYGqEyKeWqxuWCccj5MHuXjcgwYIbAmvqz2MRfWt9zgtaEKrD/uLv4m5xgQhPOEZ5W+/q4a66lx8cz0WP7DS8BL4F2QwNQxnMqB3Gk2qqO8yDPVtlhv1itpJQiaekqsiWERpGm6nefhptgUJ9N0hJNtrO/b2hbAI1td73mH6LtwfnZjl7rWwsW5RjgaZ1G9FgUbW4OaUpPVm43KQCUXhIMV6W988eX06ccO5CWH+24UhZ/T/SsB06lgp6IDTRbqV8iZfv7oU1kxu1KEca14WJocASMWvIMDncASUoCiN6Vy/A9hUnRWW59Nx1FVjvnNjfNzIzn4G2WYCtBARamdinG78aA6YV8I4IBpwaHR58r6ow2JYzDG21noiDSmzOeSjj/eODu/JZBg2FTtDBXI7qrAd23t1GKkcT6qbdAz0eHZh3RRsB8ImAk1tsaFH+z5hOZ+VKPaFKAiJqBqeYRujxTM18JK9mBczSjG7ZTmyg171ddV2ftMtTX+0OxK121fbk/mGFcyF8bZh9pLvS9p/qG2zwRhcFwBG071MornxGTZ3BRcv6OGB2AQ77mcWiNKC+Xfb7dzBfhtvAS8BLwEdokEPGCxS06kn4aXgJeAl8BtSgBjBIWfmg0wFMjDSwonQRIPFW7uw5GLl6uufsIKVGOMYZThuMZQw+ltjAU+cbLjGKeGBI7/l9VwrFsRQqLVMLJw7pvTHKc64Ad9m2FmznWc8PTJNkYBtzRUZSCDEfM7kW5sC2iAo575YASZUVNOycQ+NnbAAEAKAByKWEPlBxhgHAYAMGcbM3OwAuT0A2iA/D4/3c/qcvCbsSgMuLDi2/QPi6PMgmB7246xIRP2/3U1gBEABgw2zgeMFeYJ0INM6AtDjv04L1YrBLaHsUKMyWF5lzkPbH/F7f2bp93q7x3WeQ9Us2To0m3OL/P4nhqgE9fIH077ZZx+8RLwEniXJQBwIUcy9++66lKkk0rbiZtViijV4nbROM2bURBsKnfISCmkKgIrRkVRVCjK/S4PzXe/iyQwZVbEAiViXT+t4ShrhlGwJ65ETeWnWQsD18nSIhOAMTx5bqPzO195I/GpxnbRBeCnYhJAn8Jpj5Me3XGyRFp7/CPp2v73ZTWBFS0BGF9UuAjBHE+owXIlyASdl7atmg/PZ0n4MaV6OlJrj4+JbbAuxsKLYil8YdyvfEhq3bW+6R+QQomZ1KzUmhTBt3fF3wqsQBdmLOjf6MqkOP2BGjrdphgVf9BZba/O7ukuqFj2iWGn1tu8OLsu8ABWhQW/UMsMG4GFWmvohH9H4MJ5aamzAioacS0NxBo5Nbdv+2x9ZhiopsXfC8K8DmtErIp+c24wnD+49YhqVfSo29HbaLi8G14Jain6aktpp0bqY10psGBvM17071qWBq8sHcnPdC6HSpU1HcFbH7+qr9RU+4aaf8/9kHj8Ci8BLwEvgd0rAQ9Y7N5z62fmJeAl4CVwnQRUtwLLCKAAQwGHNH8TVcXnqmuc2O/Gmx1XfwBjB+PI0jbhLMfBb8wKAxlwktNYcKyz3tIrcRxAAAwhUhdhgtCnpVgq13Bgf34HEMAQxKFuqaCsHoMds2zSsT3pkgBU6Js8woAWX1UjTRN9lPP82lyZH0YdTv+TagAXl6b9GFjBuNkGo++31DBOATcAExgf42Qu9GkgiIEuWnXdYuABhlaZfVEGazgusiTCjXEhH/5+Xu0D0/XImPFYP3yyLcc1tgpjgTFjUYDMlX7Oq2Eckr6AbSouqBxwzUdSF8/VXPPhttt+lvNsRcLpl2uEa+U7unYWVMcCefjFS2BXSqBUY8JyclznPrpFSqd3VCYGWog1oYhWNxI4cSkMgmqeFpf0fSZ0wVajXtnK8jxOkswJtOB5y32e+RQ+7+ip2JWdAVbMzdRj1UMB3G4rldgeQIswiParGLRTGrIFRZd35aDMszTrbXVHFyqqlyLQYuBBi115SdzPk+I5j97zKTV0vMmimhVytoeHti+FpxYOZW3VtECXOqkGuIFOSzoodNBVaXUAGucq9VR1hsKLAgMOqMYDtSu6SqV0XCmVrgMr7BhvA1D8qHmhqMEGwMBiOu+6vn9L7W+roaeud660n3nlqyd0rwdPSmvcdnlwUp+5xo8eTVqo/0+NsaJzooMS4PI+NdNPZ1S8+8xDflMtLwAAIABJREFUP/XmUMDEMRH++t0rg+/qObFf8x6IYZEvHtpEv1wSEHJW7I2X9BxZbM73cwqMq7bFy+JWnNHx5wsX1EkSRd/a5ujhD6QPxdXi5XMvRv8xHQcfNRlNP2H7fl0NfdgDFjuE4//0EvAS8BLYzRLwgMVuPrt+bl4CXgJeAtdLAIPrl9WIEAMIIPoeh/RVkGH7O2O3/HOxy/o1WWtEa2HEYRwcU8Mww4BhW0vNROSWpV3CYQbjALbGpFCzGg59nNzGysBxj3EIQIDDn31Yh/FHP8YuMCbFzVIo2awM9GBsLH9BDce9GTSALOZ0NKYEY2IxpsOkSKIan/TDWO24OPhhJvDJ9lawm09SQbEdYzC5GFhTZnewDbJmTvRRLh7OOGxbjs33Y9PjIBOMSPpmXwAT5MbCb6xnfiwG7vCd43He6M9y2TM/wAdAGOQOG2av+PmpC1uHXJEM3dxHFwVYMFfmwDXBvowbw5U+n50ey394Cew6CZAaxya1f2UmaDerRbc/Di+sdiYA490AAXRM7sGxxsb9a88anqtrmW7apDfi2Wnp7thmUnfgZsW97yTgsusukF00IcCKVqNaHSdpQwydOaUZOyzH6ZGK6qRUKsGcUkFVlAuqnWRZpN9wYp4fDJPF8Tj5QbtZu+RBi110MdznU5nWr8DBDnBHQMi1RRH/AiyCPx33XTeK3TGx2z6jH3GaoyOiG5nuV9XTOZYj/iEVr/5TgRWfE0hRv/zaymG9PD4vsEKoX3gr9sSNzkQ5SOdWAIaBFeV+0K+PqaF3svyK2i9rLAIRihUxHfZEUf6m0kN9U7Up6lqPXoueuRNcQR9Ep/ym2kCgTFOpnRTwUgwEeHxJ/Twq8OIJrd8rNslYf0dRnI0lk/OL9eSkAI5XxaiYFfuCQJo1Ffveq/RQZzQG9HT6htlSC/UmWzqaPzOznP/2YCtC7yyzlt/U3+iuDZ2zbZ8W6kaXi1/nJeAl4CWwOyXgAYvdeV79rLwEvAS8BH5IAoqQHylSnloIOKaJmjLGRe4qCwtu4RNVl3bWlR6IbTAOACD4tMj/Y/qOUwznGO8P2AwYHawzsOH7U0MDIxAHOYaWsSYMNOA3y9Nr7yFjLTBuc8CXjbQbRT0bu4M+MLToA2c+x8GYxKHHWC2llLE1OIaBEmwHawEGAsYT27MfjkG2BxSgyCLrMKDYnn2JPLP6HXY8xm0slPJ4yzU0yt/LEdwcl+OZPBgzY8DoxOAErMB5hJxZ2LZ8PDNu+Q0ZIAsbA+cIkIJi2qToMvZG4cKa+o0GbvbjMtj/mVgqSjxzlZ1h551rZY+uHcbiFy+BXSUBKzh8aO9sVU7biPQ4Klqdir2gDEt5pM9C0Z/FP/uDF7O//xcfN2D0XZHBzYAGHcwAC+5x7k977jEOAyXzuwGqvCuC8J2+2xIIdHFXVMR9sRqH7SQtVlS/Ylksi/o4yY/XK0rwkrtmluaLYl2s1etVOTILORTDbDjO8lYjvPiF584lv/D0Qa5Lv3gJ3MsSQN9Cx0NnArS4ukhzwoF+7On0X66cyD8yYSFc1fnQxdCfCCaxZY80zouhCkhffGXPp+X4f1CFpZ1AC902ExVMhbR/ZBGhe3N/GdvYdNjb7Yh9ARkI4kGXs2UooKAV19MHBDIErYXBk3EtOa9aGl+59NrKp8WK+KzYDzcaLbourIdLKqJ9fu30Yja70sm0/weVGqor4EMAhlsQ+HFKr8uhvqNL743i/IAKfdNfJkCjp2M3YVdoG9OhAUlIZdrTPif7G8GbkuUhfb+u5od+p34cgBEpUb+s5lkWt3sl+O28BLwEvATucQl4wOIeP4F++F4CXgJeAj+iBAAUfkENxzcsAQywrlv6uVkXzY1c/+XEBfNntY4USzRSJWHQsZ0BHBgbGEQYcHziQDs57ZOURhg2E6q3mtWFALzA+U0/5foKON4xxqyQtBlL5mzn0xzzBhbYNgZ6mPPemA6Mk2PgpMdwsjoW+jpx4huogNEDEMB2FCe0FFn0D63eCo0zdpurMUwMEAC0sfoc9F8GJMrAix2TbayuhDFVWMexWc/+HJ9PDGhLIcW5YoysN+YKYzSZmOOS7fndABlkjrHJeIlkQy5sC0CTuMr8d1z94MfceF395szN0gAgE87VMbUvMEC/eAnsQgkEDx1diutVxYBmOa01SrKaakeMFYXuxLZItjtDZa9w/X/+R690Tl/YIuWS3WvvqDhuwYCAOWEsivJxf3RX2Ds6at/ZvSQBA+iUaiyP40hMyvCIcIjHAhcq81O+rHoph5M0V4kUpYkKgrRSCTsKDQ/1WyWqhCt5UXTFxBgJ3Fj/9pltX4j7Xjr5fqzXSWDKrkBXQn81JvEVPeuXY2ljraW8M7snf3TYCb6jGhZPBNHEaf7+qQ5l7Fbrk/RPsQpKP7p+dl5FpitKdnQrUsTbnhB0StOdd3ZE8MjO4+/szN4LlsYTPZfAnL26tzv19ihQjYlOfXYoLkR0gHRNjdnhF1ScWwyM4LfFhviIgJcP7uhUOmRwRPU49vbWm51KLWlo+6KdBb/bXBjUBEJkAiRIK0pQDCAJtgN67YtqFOqmvt1xfRJchMzRS6lJgW4KALSh9FtvjAbBgrTesr5sw0D2BFOh73vAwt/PXgJeAl4C94kEPGBxn5xoP00vAS8BL4GpBHCCYwBZeiDeA3U38+GKSze23NLnDrioijEBoIFzHCc5BgKR/jixyYt7bPob6wy8YBso30ZNx/GNkx2j66QaBhYOdgwnfrPC2uxvVQeNqcAn0cxWl4GhM5Zy6iPWWQomc87zyfEsVRTF/Dju1TleBRZYJhFf022ZJ8CEjYFt+W4gB4YXf5ePxdg4FnOAjWAAQ9l5uHMd/Zmj00CTsiFqKWms5oQBFzY3i+gzGViNikkamGljbmxv+3IerfYIRiFzRv4YvHwuuaD6nBudf8SF9UV35B/NudP/hLkxV+ZtDJm3Ig+nAvQfXgL3ugSU2ibc7Azlfw3jRqMyq7Q3c3LWziqqvLHdG1XllB3px0SR6HJGuSty2p5TqqgewIHAhTseXT4FNDxAca9feO+B8aseBe+0FaV+Oi42xcpwnCzqxVHRdV5XOHisiyzKimKcjZUiKspXYt0MSokzr6jzeDjOK3kx+sFwlKAPlNk+d3Vmb8NQsvei8yyku3qK3msH5x4gDRTX8GcnupPACl3nLqqJfBq7N5oLxbyqLPSkYf3+VCdCLyKQA90InRf9EUQ7Vr2Gjmo4LI+6NafUSO/EXOmfxfRh9DrarcAK9kEP/g9qABbofh+Z3AShRhrlD1ZqqaMg9qhfObPnxFp/8fDGB4/+xNnTG+fnuirM/ZHLry9/sL/VvJrGSk1gzNWB6LuKhNc2zs6vqeD2vOpWPLZ5fu7ZPQ9ceX5+/9ZJ9Y88CBLCFvia9tsnmXxbrIxnqo3xjFgW6JbGvmZsAByke3pKrVmfVfascfC6vv97tc/tECLnigCcUGBT4NNC7ZCO/9NLwEvAS2CXSsADFrv0xPppeQl4CXgJ3EQC1KYAOLBofjm8g66rHZxz7cdnXTzTc1GMYx8LhRREGE2AFPzNO4PfcHjTB38bw4L10LWJnsKowPHNNhgwFHqmtgXmD1R36PcYiRh/Bh6Yo51hAwTY+Mypz/bm1N/JtGAfc9JjhLIPY8YIMhDEnPX8ZkwMgAoMT0txZf3waUaiHYt1gAP8bTR9jsV8DAhhm53jZh3zNSCkzBwpb2uOSD7t3WzbloEcvmPkIduy89JAEANaTJ5mHDKGH0z3pZ4FTJu6i9ufdu0PtFyyVXFhAxkDQpmhzPg4DteMX7wEdo0EACtG4ywajtK4P0rma9X4wGCYHhYocaxZrwxUzLrQ38lcO74wP9sIev1xXWDFtlgX1LYYyTk6ereYFrtGyH4i7zkJTIu5yycbVHWNN4VCTNIaaqmrdoXAuvyKflzI81wuW97/xXKQBycSl9fFrhjJeRsPRqmAvHBNNYh5971nAIsyQ0nsj+CVk1eCmVYtUB2ayXnQZzBlKU3+9uDFe+7yvNMDQldCL4V5QFFn3QhS8KR9xRXlB4zcm7VW8Whj1jWDMDita/+FdByfVP2Gh5XRiCCOn1CthlaaRMONc/PPy8l/SJ9u1EPl+rGXM9oTZnMZlOAeKzOPb4e6ga7HdvNiNMCmXRabYlipZkPVmLg8t3c7EKtivdYepQsHtvZH1WyftltePLw5jKvZYn+rMUjGcaMqlVBAjEsGVZelqsMh1ghNDJLhhZf3xQItVmb3dH9Gfx8SOPGGRrmufv4NMtXfi6qN8V0BFn2lnPobktVMVMkXVMMCHfPP1I6pwVp5QE2FPoJwsN1Oh91i0QX5yg2KfpDi6mfUXlHDNvGLl4CXgJeAl8B9IAEPWNwHJ9lP0UvAS8BLoCQBwACc+zjribLfcJW5plv919SxGLjqoee17hE1jAOMJgwDtjfnPF0Zq8DSGAFSQPuGxXBODYc4+wAa4OyGyo3BRfokAAwMMIwy1hmAUHbY4zC3It+2jTEgOH65TkQ5PYuxEayA9Z9qWyuWTaFxYycwb+YGA4Sx71yMsWBhcvauLLMmMLoAKmxc1nc5/dTOOXEcxmjrDYCxOdqnsSYMeDFwwsZTBivKoIalyLJ15ZRcyPxJtZfUuAYYPymiXnPxUuzGl2U4ZpGrHZ1xo1NEvlmqLqtTcgMx+VVeAvemBAQ6BPOz9Vi4RDPPioO9QXJczApFkAc4cJtiXQBkzg6TbO9sq/YD/bYs9kUiR+3ZRq2yefzQwrYHLe7Nc+9HLe9gHI50rZ9Tyqd9YhE1kyQ7mObFHq2r5C4fBGGYuKyYVTr7VPfIUpDnLb1UX5a3cjHMghP1Wv1Ks1a9oFoWg/daLYvf+OLL0XMvnYvkYK5p7Lxjo/E4DevVStZsVgZ6OaZrm31SrPm6L/f3zYC+hU70VyZi0IUBu0IVJyb1K5QSqlFruiRL47nNi+3DcrwXqk3x6Znl3j5VeUmHnfp2Y27gOlfa2+df3BeJXVAfq27Fj1qvQvy9iUo4AQNcsKn/0J/LiwWQsM4YsG935tDhASzQuwUQFL8/s9Id7n3ocqKxf0/jWxXgkjcX+gcr9QQGVay5o8dW4ko6P7t3e0vrz2puC2JinBd48ZHulTbsq+9qzrnAiYc01hXmmoziTHJ5TnJ5n8CJL+1/+PJ57fsz1LNQaqlM4M1/Eob5ga1LM5Uz3ztwav7A1ktLhze+W2uPvyQAAz32pFpH/UXatnr2ew/M11qbYrn0vpaO+k8Xk5Jq1y3lVFmebXh/379+9l4CXgL3iQQ8YHGfnGg/TS8BLwEvgakE/po+Lc0RTusZ13rfyC39fNVVlqoualOMG0MCpzYGAQ486OWWaslYFXSHU88KWwNEUL8CIIAaGETwsy1OcYAMLA/AAZzp9Mlys0gxq/FgjnurecH2VlQbwMUACuvLDBiOS65bcun+htovqVFwGqCFPo9P92U8xqSw2hTlMRm4YEAF5qyxIoxVwdzebjFWRrkvY0MYKGPprjhOue4F/TLmG41p5zq23Ql48Lelt2J+MF/on/PONQCYtOSipmSl2MKlz1Xc8PWBu3iKcwiow75sxzXzv91inv5nL4F7RgJiSwT1SlwPWm5e6fyPjsbJMWW90TMlmB+OUzlxQrGYiihJ0vluT/n843AQBHlLUeitKCpOC7gYqb5FJqdn4iO175nT7gd6VQKKZQ5yARW5fLM9OfXHAitGYeCGAivacvTXVUC4yENX1e+6PVxDDtxCvzeiKKoKzOvWKvGM0krNdPoj6At3PD3ajU6kWBXhmYtb1fXNQV1zmomiYF73a5DlRa66NPpaDLq90ZbSWw3qtTgRuyrV/cs72LMt7rM7g5RCmjJ6F/oNumRXK9rVhoon6GpOhsGZcT94rr9VrQy25p/KsuAJpXmqKx1SQ2mTNnsbzWrncjtpLfVhFURywBeq66AsasoqFRTn9GmpUW8kWfQy9Ou62Aau2kxUkDqJlErqSp4HY9WPeLuzcUu/jfpcEXjymMZxWOOYa84N/0prsbcsZsUZHadWa41XBRZcCaLioLYBDIGBQbqlGWmaK2JBfLe12O/tjy+fV32LYt/Dl18VUBFr/0sCKNZf+eoD5zT3g+r7E0Ua5p01VbFYK57avDD7C7rH/unBxy+cVL+PS55z9dbocTFSGq2F/ujCy3uPbF+eid74xtFTKsYdPPG575/S+guS6/gHX31gtr/RPDjqNR6vz4Tz9ZnF57cunhSjZfj+EgJETQwCom6HYXKfXdF+ul4CXgJeArtXArd88e3eqfuZeQl4CXgJ3JcSII0DQANR9NDah67xeMVlSgmUj1WEMzLQAVABRwTphwAJcF6Tlxb6NkY+vHcaDAy2w8kNo4LILgABqNs4yAFAOI7VgJhEPE4l/3Zsg6vsj6vpp6DsA1rQH7UcMPZs3zIQQLfm/IdRAGjC78+qfXw6VsZCjlyrqcF2BmQY24N+DFQww9aAB0thZWmajCVR3t6AFGNqsK8BHaVUXNfYGRyPcZRzFluKq6moJh8GSJTlZr+X1/Gd8wyYgqzpi3MFWwJWCQaqyVTRdeHrbvjmHgxvFy2yPecX+SB/rhX68ouXwK6QAOliLlzu1JMsa8l5uU+O1yUxKNqKIF1pNKo1OWerURi1KlHQl/dJkejhQTlNzucuuKgIXDk+Xb03GLdq1ShXwW7u7YnT0y9eAveIBILRKInzLK/q+g6rsRJEFcr4khVrivNe1H2gd1Q4VLx3XxHf7TgsMvywSglVk9tyXQBAMhqlVQEbAi3CEKDgqcOz70oh+tuVp5ge0eW1bi1N8zndoItpns4LYFkU2qII+bwQ6FLUVCxcDlWlthIYXwR9ATadJM3QKxLPtrhdSe+a7Uxf+ppm9N9NZqU1tXbhKtKUGnPF1+ozUXDh5aV2b2NhVnUfmgrpOKR6DVKX8pFAgUOqxzAebtf0X6Wj1EnrWgfwkCXD+LTKT5cBCwJD9suJTw0JpVwrAEgKMROkblMrIytUBHtT6ZpOKv1SPNiuiblQJhTfVObUaKNeBGmkYETPktJKIEDWXu5F1XqytnV5pqlxtlVQu6tjDavNcVXFsp/QXNHHYR2j76HXc/+i621pnAcFZsy05vsdgRLo/4tKE9XXeKtKITW/76HLLw82G5p4lOp3VRd3n9TMagIejp9/ee+xFdXEqLVG+8M4f4DjCYQp5g9sR4c/cN6d/u7Bh5Nh/ZfHeZB/418+9a8kr8sq3L2ivgkw0lhIX1VUJVSlqArer6ZX7zUiBQFGk4Ae1a+4q8+bXXMX+Il4CXgJeAncAxLwgMU9cJL8EL0EvAS8BN5BCVhKJiLLcPzLlb4eu2g2c8UQBzWRVhgxE+NFDSaBMS0ADwAv2A8DA+c7jnBL8YRjHFABI4f+MTAACHCcm/O+DDTcqAg1fdI/jf2XpnOnD/tOH8YS4OedEVeAHYAUABG/pvamGrmKOR7Od/rBIgRssTEYiLIzPdP08NfVprBUWDeaC9ubhUXfzMPAA36z45SLarO+TPsvMy34rQyW2G87qzqynvNglq7VB7HxA0BgRJMi639V4zzzNwDUG65+YuR6Lyau+YDNjXHTh6Xxsn78p5fAPSsBwIrL672qQmGbpLrpDUaHwiA4rIjzBUWOzyogu1mJwkGaZu1mozqWU3eUyYclJ2hbKaHmlD5qqO3k9YlwdKZaN1KfmRy2Pj3FPXtV3HcDz0lvVq3GMCXWoiBYEFCxlo+Tal4Eib6TKk2Xft7XCy5T+qhanhaJUA29cwO5//NQKdRmVbBbmf4r2JFX9Yi7tACYnDq/2RAAsSDAQiBFdlzjPqxaG3v7w3FbAMV6HMnxqjodip9fU92ObrUavjkYFRd1L/dVtwZdAn3HL/ePBNDd0IGuLzihp3hbGPTc/mK/IK7N/la72d1oKlmTmxXDwApQHwJoaC/2q/2t+rLAiqAxM+yrsPSf1iujiW65IzXUKW0vB37mBEw04kqWqu7FrFIrTWpmZOM4SUfRpbiWrQ+71ccqTWVjSyMxPSwW5odOiqWFQpdno6Nq6JjfFWhyYHZvp7l4aPOkjnVajIZXBB4szK5047iedJTiaa+0ZYJ+0OvYl/cY9zDf0YcJNkJvXtV2qwIvWLcYBdm25j9JmHXoifPNwXb9/zj3okSUBR/Wum+o6TFSrIkd8j6BD+imk9SKAiu2iyxsa9+oOT8IBHgsSU77VAtkQVryfjFWAF0Iarpqb4jxFVUb2BwbSgelYucFOqgt/6++fIk/fNHtH7om/AovAS8BL4FdKwEPWOzaU+sn5iXgJeAlcEMJmEPeimUrFdS8DJEsdWGLuhI494nWwlDA6MD4AKjAoMB44W8MJJzjfMe4AMTA8AGc+KgaRgjGDcYPBiEGFo5wS3dkA9vJIsCItPQSjIXv7Mt6mAGMi3EQEUa/9GmOfgMPYHkAbnBswBPAiw9Nx8N6xgqgwrH5G+DFCnob8FEGLRirsSlsfJYaqhwGd6O5IBMWQAKzPpmTsTaMlWFAA3PD+QO4cFrt2HT/nawOtuP87CzaXX6nl9NMGeMDmcIuoV/yJJ9Ue0gNhk3DZV05pWLOuRmyZabIdCj+w0vg3pSAoqgpwBsqqrouZ2tb6W1ayms/R+7+RjVuV6tRhd+6/dG8nLQuHebV3iCdr1bCSIW4Nxq1aCQn6KyKdc/Uq1Gsm3IggKOvPnlGvSfS4tybZ8aP+k5KYFp4e6R7YCML8jml5i+iIIJtUVU0c10AXlVxzbGcqStiUSiK2g3JsA/DQte8OBnBUJwL8kiFxTCt/JsvQ6q8e8tWZxiNxmlzMEpWNKdlgY2H1I7ovp4pcjk8g0BMqnCfgIvZOIovK9nVeUVu5/VaNEgShZrHUTYcJZba8u5NxB/5TkrAdFec/m8tusDzNFCRadcZdqJvhZX6U6rx0AZgyPpS98SSEHPBKa1SsnBwszK7L2wp7RH1J6gDkauOQ2f1jeVvCIz4gFg8++lYjIpGfXawGcf5vECDVnNmuK2C1uNqM66OutWBClpvDLv1N6v5+IzqSixWGumFpF/ZFGDxszcRiOl56MO2oNu94MLiVY3liICJRIW0RzN7Ol8TsPJ4a6l3TMCKiocX6MPsT2ol9kfHQwasQ0+2dKCwNtAz0ZFXmJs+J4FKSufUPPHh08+sn1n4E9WuaIhl8cdaTzqs50f9avviayvD40+ffkX7LGrbeREsAskjEANDtUGKMxrHCQEbj2kfGqlaCUxiXKKvBGJ4uM0sTbqqo9PaEQXwqLb5hBqsGJjgntl4kwvEr/YS8BLwEthNEvCAxW46m34uXgJeAl4Ct5YAznFL93S1DkSyWbjRRZkXP4cRR7ThMTW+09bUiMTHoPieGgABfRhAAZiBkWOFsOmTqH2c9DtTGO10gJdZFwYGYEgBRtDfoenxODbHZRuMKAwVIsp4h+G4t2LTGFeAJm9Mx0gtDfpiTh9Um0SLqU0ixab96OMao4Rty4Ww+Y3F7CY7PvKjL+Zq9ThuNBeAFcYHSGLsEPrbeQzmhpxfno4J+f2+2l9Xg/VCHRAcoiZ7+uBvm3cZCMKoZB6MZydIwnkCrDHwCFkxRsk03HaNRw64AaKb/G6Rs8yP8+0XL4H3vAQEStxsjBOQUOBCVeyIZlyJFmouOCxg4uCwP1rMK5FS3BRVFePeo5umNtOubY6TrJqmaSMKSXwTXlZO/CLJisZ2d7Sszl7XvmmjFgcCM0iLk3uWxXv+8vADfEsCuWo4jPWSGIs9lLpIcEQRNBXRPKu3htYHsYALvUTyoereKmY6GCuBzYJSLBW6f/TyySsq1E09i0C1XMK7mVJpuzfSKFyrP0iXsyI/LPbIfqW3WtF9HEZxJCdosaSaM2OBGc3hKGtkWVYRSFGhTk2tGqfjNAt1Dw+Yw/S9+UPXiUAef+3sPgmgD6EPXlvGSoTWk8YVxm7v8vH8UJ71VIMh3ydWhNtebYtRELqFQ5tJc75fEWuhAIwQQDASIyKUE/5BARYNsQk+IqaDXifRpPyCtnmyNTc8EzeSmKraM/s6a2IhpKoDsV9Mg9QVabXSHB/S916jOlzPk3CQ59Ev/xjifkLgygtK3/SsUjFt1Jrj4oGPnjyq4y8IKJjXJwAKeitgBDop+iR6ntVjs0NyHwCA8PmKmtWUY1908XalkTy6cnztDaV4Oi+WBXr6xJ+kORw99dyhfPnI+u8rLdXrmu9PZUm8JCbFPKnmlo6uFwIvXhXZ6YieN4yBwJmybrwo0GIzrtWLuFpTf2PJ8BouQRFxzhlghU8J9WNcIH4XLwEvAS+Be1ECHrC4F8+aH7OXgJeAl8CPLwEc6AAROK5R/kO3+a3YLf5M7LKBpXbCYY3jG4MGp/bJ6XfSKlH4ju0wcnCIm/ObT3OS22/llE824puxLNgXmjpGFWCIRb6xHouFcWA44dhn7DAoOCaggUWCMS6+42RnfwAMwAorGs72bIPz0sAJ5ml1HvjNimgbSGFzsrlYWimOsbPgtrEsjBFBBBv9YxSXQQ9jjSATxsaYMQSJNGNuBsjAVIEBwjHZjvPBtsyZMRvLhe8mV2OcGKuFuVr6KGRBFB19mSzQA+Zdui2GjaaTdxgnY6E/wCjmWablM2a/eAncaxKY3AeKrJ4Uklde++VhXhzTykPjJG8Mx/0DcRjGqepayJEZVHpJqhQXmb7nYRQOxbxYHCXKhRO4roCLkdLIVJRSZyyGRapmzKx7TSZ+vPevBHjOD/VWWguK4owuYN0bTimhihO5rnNBdJnSRW3p76FyQ20qLVpVnsNIzAVxEtxlMS+UrsXFAvXC1Y3eXU2HpntTQwrqaZ4viQG1wt2otE/LYlKsCKjoyGNcKVTFQhSRUKDFXjlKa7qHWwIhU32mQZKuCYjhnQiLM4GBcv9eFvfNzNElCXpBP4NrmuTQAAAgAElEQVSJSw2vqwW3tUYpnCozK4Ogv5m8KMZDrdYcxXEtnZvd00lVdyFUYepUKZcygRRvZmm4un5W/v0iEOgQ7VETOaDo6p6Z6KViZKzW5wZD1Y44o21WizSSTlXMqvbFhjTRgfZvRWn0/mRQ2dtda50VE+EpgSA/zokYa7+DAkvQ0TcEULQEXsB4Rpd7fqrHWW04nP8ABuiE6MromdTagGFNEAvrABP4JIgIvfwnp9s8o3fjHhXjXj/30r5LYoLA0r2qg6oOlOpvLD7/xfe99uG/9p0XxaaYiyrpoVrTHRZIM9tZbdcF6pzRPQgQQlATwTm2TIOegnoYV7aUGuoHYWXwSDa6jkjBfpwvf4/+OFeI38dLwEvAS+AelMBNEyTeg3PxQ/YS8BLwEvASuD0J4OjGmY7TvuHGFxT3pSwQySUMGKN+YzFhxOMcx2GNc54IK6wHPjFqzKriXYLhw984zHFyG7vCmBc2sp2WWBkYAEDBkCTMH2CC4xijwoAGnAoYTzAPiAKjP5zuk+KZ03FyfIwafmPsAAYYXYABbMMxLDWTGa44Mo11UY7eYl15LsiBdYxxZ5RX2YhiTMjCaknYvA1AMLYJBjNprJg7sn1JDePvk2ovqiF/jlMGhJDNJGJcjaV8XORQTmFlUaNszzHomzERZUdkG+sHrvHgvBudy108z9/Ij2uDa8SzK6ZC9h/3rASuPafktVRwddgWM8LJgblJChz9Xa1VokQFtYkqr9DGSdpU9HXUblXl/CwCOWoXtG5JkdvNZr06nmlVYxXdVr2LaHY4Tu3Zcc8KyA/8/pLA1ClPuqdNOfpPjtP0+5LAtwRKvKCXx+sqOi8UQtHjckAWCirXvdIWuygUUNcR6Heu2YguCMhbBQbgfXO3nPy/85U3YtWtCFRUeygQcizwpaYMbrO5vKgaaz4UwJIkaSJQck5O0jiIgqEYFyM5dlVHIDs2HqUPax5tgRdV3c+3Ven4/rpSdvVs0QfR0XDWT9gQiRgWgy2lCasVG7Mryczcvu1Xqo2xAkeCy0oDtdlaGCTVZrI27lVPiU2wlmfBq2e+d/A5AQ1bYlZ8Q874UGyCUCCE1W5zAiaKwXZjMOzU6wI2otWTC91Rr5bU2mMpX8WcAI4Z6llon5VRt/aUtt9Svz+O4FeVCGr9yqnFh09/59AljYXaEgAU6JjorZam9Wl9R+9Fl0YPhJYIe/qkGilDCZwBrCDwiH3RQwF3JmKayquqmhQfevBjb54VKPE1ARhf0PrPqH2U2hQqyn3o5T956GXdZ38g8Abm8JcGnfrvbl6Y/ePxoMp9RnongI4yu2Oiz4I3CtiJgzB6JNItSeHt0oJeanp/eb3/7iXgJeAl4CWwSyXgGRa79MT6aXkJeAl4CdxEAqb9W/0DmWyLiq6v1ZwSI2gf3gvmpMZZjjPdUhud13fo3y+o/Zya1YHgE2f420U9ldNDcWz+5liwKlis2LOleXpO6yjGh0GJkULDeGIdYAQGlS1lBgFABpFiGEJWQ8JqVBjAgMMeMIToMQwxDDQDEBhXuXj1TsuRcdLv0ek+VhC7NJzJVwM6kA1AELIsp2nid1JWcSz6MObEk/pOFBljslRbxp6wguQAMABEyMZACzsecuK75dQ31gcgBPvQF/sbiwJZ7XPy1wisiMhfUJqI9fFjWc87BeL/9hK4ixLgPqBYcFvFeetiRawoMrulIto1ARU1pbnphiooLD8RxbiFQwQ1RY/vVbqY/nCQKmA7aLXqlZ6izeUXVbKPKO7LH5o1apVCjk5/f9zFE+sP/eNJQCBDrjRIfd0PF7OsGFUqQUd1XdYF0K0Ih6gWQTCnS31W/sK6nIZrejWsCruTk7dQyppgW/dPV7/f1WLVS/NNpyxVcZZmjf4gaoopoWCGYkXOZ+EVxciNs5poUXCg2mKFDPWCG+QuqAjkmIki11CkRiLQMhOjRKjGpMAw70Ufvf3jXVL32l7ojQSI4KSfRPrnChlRiiO3fjbqDzvZmtIefUDXzpO63mMBDgIpFPc/OxxFy70iGcYvCGhYWDy08VfkmA/EtpgRWBHIMa+aFm/Fg6q/Pf2NxkDaZiGQgzRQUVxNZ1TfQfeWqEvNJBb7YFvMilmuvElqNucoDPPIbQoUHRLwQTmr5OpXmqr2cvfXxLT4E/19StoguvpHpte1BdEQ9II+zbUOk5YAHIpxw6Iw/Rg9Fx2U8byqdny6D+P6igCahb0PXjncvdIeX3hlzwOa/xGtx4Y4rTm4y28sH//ab3/oz449feabYlZ0Lr22skfyeUJgDHbEp6YyLwf9TNi9Yka9mo5686qas6ymVabaTnT1qwE2/h69zUvDb+Yl4CXgJXDvS8ADFvf+OfQz8BLwEvAS+FEkgDGC051ofqyqoaLrmy7tDFxQwzqApm31K3Bwszyj9lk1wAUrxk10mtVvKBecNmCiDFDsBEnoH2OJhe8YRl9Xw0nPGIh4w6nONsasADiBWYHxhBFl9RuMhWHpmeiPuWGYsQ6wxdIfkWKJyC5Li8V2HMvqQTAeHDCMnf3L1pIBGnwyBow8fmcc5TRXNtey04PtWUxOGFxWMJxIPAMPMFIBWmyO1N0gXy+GpI3HCmLTH3NDZuVj2fEx7ujbFivUjaG6MN2HvpBxxxXjoQs1pOEbAB5WH8SYHT4lVEmQ/us9J4FrHg95MVsqzrugVE9LYlAo6rpYlbO2JcersIhiIM+m8n2H8RhHp1LeCLlQkGeu3B95Q/kuQvlhenla9LMwH4VhVAO00OY8o7yT8xaXhep8sEWZscbf1+SmGiD33IW1GwYs4GFQqUSFWEQDnRyxD9ySrvQoyIrjAu5U+8EJyAhSl4dDOfpHYiVcSpK8I0BPYMd1APcdFweARac/bvX7+UK7WZ3T/T0SCFFXurbtYpRG8t/OKo1boMI1ghrzWbEpwljFxrV+Q3Mdyx+auLyo6yJs6WVnta3u+Dz8Ae+4BNBtcPKzXPfggWnRvRJmg23xHwon9k3RCiPXF1DxhgCGh8TQWdTnhgq77K/U0/cpBVJ188LccLBdb25fnhHocX3yCpz3cuZvifEQC+SgSPUgjOtHKtVMJILCRXE2ELNCYMXkeCzohvt+BImw/aTAN4/XYaf2ffU3L9bH0frM6MsCLv6CfkB/RM9GbyVQBoCC7+xngUjowuh+BP3QJ8FJ6KNsxzsORi7boJ/y/bzSZAVHnzoDs6O6fnrh2wJwOpofNsSCQJyf7a03n3jxS4+8qb+ZGcFGBAlx/N9RI+gItsTVWnpXG9/3STBKTKdKOZlKfEyFovXYHJwrHyAgIfjFS8BLwEvgfpGAByzulzPt5+kl4CXgJXBVAhZ9X0p/INstvZK57rcvuvYj/I4RY6wJAIBfUgO8wHA5NTUaMEIw+nCmlxczJiwVlB2PfvhugAAGDNvApICWToQbx8RhjiFJw8DCYAKg4Di8s4yJwDHpg99pBlwwL8aJEUaxcNbz9zE1jCyOCQX+qel3+mEBvLAxWtRXeS58Z3xWgBAnvqVbMpbFTkOKvw0Y4hhmlAH0AP7ApGDexryAtQEIwd/0D7BAZBtGpNHgDeigX4za8jHYz1JdGaOCfljH38gOtgfyYH9kTDXRr7jhqRMu61Zc57mdaa6sP8bvFy+Be1ECBp5Gcn7EFP/U50CAg54veax0UKpVEdVURHio9E7r5LpXRv+9cmTG4yypRSJm6MmQ9AdJS7HaTUWkK++MUkgFwWg4TIdKKZW1GlY65l4Uz7s3ZoEU9kwsA752PjiwvQcCbcv3mwI/HtB458/TNJVTIqZFquufAtxiDwVJJYi+rXoP/bwIFCserOF0VZGLgf5bFZB3UQyMvkq9jCnc/c6P6vZ73OoMg9E4K/rDtB7HYUP3YbjdH5HXcCOKg1UBK3UBLmSVGYp9UStUc0P3ulgVenFGwbYKcPfFsAr1Ytd0gkktq7tZQPz2Z+63/PNI4Ftf/c3ig5/428aURRcj/eW1ZdQLls6+0Lg4u9cdasyNL4oNIdAiXwwipRHMw+Vht7Y87lPWJSi2LszGl19fJs3Yd1SH4lNkMHrLxz7p8jUxMx4o8npf8PaMtqv3ksgplZKr1FIBDPWG1u/cBz2YYJUycIEuazqqBcFcJwaOK3DkkNJC9bMsnF04uDWncZPSCb0Rh/+X1XgWo2sCPtA/QS/oh+ib6NgADix8Zz+ABYJ9CKzhO/tPUphS50kMkdOqZ9FSTY8DF19duSC5fECgzYPTotror2WmNAEy6J7o7Maevl5vVkVu1bDIA1GgBCxqs2uvBOaMHowez1x8kMD0RPkPLwEvAS+B3SwBD1js5rPr5+Yl4CXgJYBWL8tBiyn3OL+JcuL5fxUg6D0/cAf/ftvNffiY/ib6Cac222DQEZGP8x+jDqOGSCso4RguGA4s5ZRHZee9GSIYWRyf7TBY6Nsc+RT/w1DiuDSMJxzrOPKtqLYZThaBxac51hmjzQUjhu+MD+OG4oMnp/0zB4wdDCXACo7BXBiLgRHMBUMRw4zfOb4ZiBY2ZwWu2ZaFfW1+ZUccv5X/Nocd6+ifcT6mBgvE6nRgKDJmY5Ywvo+rWdFuZGbMEhszfTFmS/HFONkPubDeFvsb+VrBbs4hx1afRd0l201XWWE7AzkMkLH8xaXu/FcvgXtKApPoaaWC6igKe7+eiXiIcqLE07CoNOuBgq1z1d/NqlpXUfmKvNqICgqnZlka1OuVgRy4iRy6Ub0W9QRcDARcrCkdVLYwa0Sze0oe7/pgp2CFPTd5lvI8stR/5onieWOp53jeWHvXx+cP8JYEAC7kqB+LMdRRPYiRQDuxENwFUYpalShMgfjERNK/oq/7Zqj7SHUhMgs+uGui7A8Trpduf5RcEBtqXeChIrsLYS8U11atCt6FSgmlgU90F923ifygkUCMA5rjgt7eSTWKr5BJJy5yrs+7Vo/jrgnx/j0wz53Tav9R7cGyGIRdDdfP7Hvsta9V51oL43jPA6sLYlPUGnODc2JFKB1Upbl+bj5XTYYwHVYGAglWlerokUpzrHRQgcvGqpH0FgjR1ncVxA5JVXZ1ySM3FBNDrAtAj51gxWSLqR5WHtZtUtCCGdge+anFl1aOrWfLx9ZIoYpubemd0A+PqwEYMCJ0Y2NQcJ9YLTuADnRPGsE/31azVKywMNBF58M476sY+baAkSfU9vTWW7WN83OxgIsZzfeYtkGvJeAIeVNLjmMxFmNKl+eIvTJKh/1KJtJvIYZFaTmp79Tl8GDFdRLzf3gJeAl4CexuCXjAYnefXz87LwEvAS+BnRIwh5A52WVGDGK3/ezY1fZtuMYDRHFhYABQ4NwnCovoKory/WU1nBQYLwAZ/I7D3aK9jH1gKZbMKcUxccJjoOAUKBeLZh3GEyADhgz9GqjCJ/uW6z+UWQRWQ4P9cNwzbsZPZBr7sP8xNdJNQW8n5RIGF2Owuhf0D+OAueBMszRPjKMcaWbgg5mcBhwYk0SbX6OqAybYdozRHP9sg1wBJaxuBowKgB8DgwBwGA9GJtFvVuOCfiz91CQf//QY9p2+OTc2L0AH24axWEoAzp0xVahfQaqtp13j4ZbrvqRaJg1zKNKfgTM7WRf85hcvgXtJAlzDyk4edHVzrqt49uEsSxaVOqYt3KI6HGcD6lMozHooICKSY7NLHQtFbV8ZjYtEwIQyyzilfwq2FYndVSqc7XotTuZn6nhUckX/+2jP6dUwBSqCTm+kwuQxz9qWZNaU7GJF5s/IgZyl47yrp1M1DsO+nppdOZqtvk6Z5eZlegfvsClowXs6J7WSPkkH1dA503skEBkhB1y6yojJJu/z7G4V2y6LRdfZWAjFpcFg/KY+dYuHK7pdj+v6igRizEGf0ODrun8rAJbT9+Iixbfr1egk9TnG45S5WlDBHZS6P9RdlAB6KgyAP1L7mNqJyVhEkQijymeyJFjeutRS2rDKiVp7lM3v36qqYPQ4rqRrqsmw7/xL+3oCHKoCHNC1HldNh3zx0Kb2zZ3SMZ1TaqYoS+JIxbS/r22UfnASCHKNiqd1a6pvYUE/O8VgOjXvF+419EF0NdKEvu0yAUVUVF4skM0X/+jhV973mVe/M79ve3+lkfycoJEVpUz7vuKXvjudL0E86MawqifvMjV0aRr6J+CABQoBZDAGxgwAga44UF8/IbbI++b2deaac8MrvY3mVztXWnWxSo6oLgfPDPanP0AO6oUAgDysVg6osTkBiAr0ERtqMpGdpOWJHNBzyzr2rUTif/cS8BLwEvASuIcl4AGLe/jk+aF7CXgJeAn8GBJA0cdowlEOWKBI4yx2zQflKLpq6qhhlODAJ/LKovc/r+8YLxgLOJf4nb7eKt79lkPdnPkYWlYY2pzkrMMYo19Lw2Q1EnCw41A3MAXAYKfVYgW7ber0ixOCPkgtheMfw5PtMMZIOUX0HI5/o8CX++RY7GPOMfbDyMIoM+fZtbg4rWOMjJu5T5w2aoA2ZlkZwGDGWJm9gWw5FnJnPYABY7JaESbr8nisHzs3dnwDKjAay7x5xoRhyDpkYwAF45wYmNN5MQdAE87Padf/fkt1LPa60SX65RwbkMNYfshq1Dq/eAncKxK4dn/0BuOGct0rlYXbBJyg4K4clkoPFdSiMB4pFrsvB4yAzqJXq8cNOTzdKElV1DfP5dw8I6DjgrbdiOMY8IJ7CrDCA3rTK8HACsm5oroIM0SxC+lZSqkTkOYbo6RYkdNsRs7vbdUKGYqtwuPlAs48QCD9YYyLyXPUA0F39habAhBjsS2MqTcSO8GS3Nh1PnkXvRfAiv0rM7kAi2B5vpltbA8vqA5NICCxJsAlUB2aZV1/kahTzGFVt/Ci7ueGHNIU4R7WKvEa97621TMg3MqL1ECzOyt0f7S7IgGlhcqVFgqGBfobbIKrgAUXN/UT0vGJdOiGKiq9oNoT63LEv1mtJ0Nd/P2Ns/N7BAjsF5tCmdKUUixSdfqV7njvg6vbct5nSonUVdHpnmo7FIOt+mtbl2bfEIhwTs+5IwIqYEqgm/KMu9WCDkez2nG32n7yu45RkwYYKEXVvtf+w/FX9z1yOZ3ft/X9mZUuRcRPSKMbqHaGGEfXMGHGgh6N/oj+T8AO48ROoO4bD2ruD0ALdGP0fxZ0TdZX1F8ctnNV5XA9ARUVFRZ/mXoeGgsgw/NqFP/+aTX0SXTRnXolz/6eduhmabIHc2SSXuutGcPO4LhvBVu99Zv/5iXgJeAl4CWwSyXgAYtdemL9tLwEvAS8BG4iAYwLc+bjDMdoSF3vxdRFM1YrwRgROLupc/D/s/cmQJZd533fudvbep+efUBgsIMECW4SaVKUKJESaUuUZEm2ynZJVmIlcSmOnLiccqrs2FWOXeWUUpFluVxJKVZF8hKKUkRbijZSpAgS3EmIC/YBMOgZzNrd0+vb75b/7837Bnd6poEBiAFmus+tOfNe33fvuef87/Z93/9b8MDCKwqvrLvVzEBv0QEYmsxTrEpiYAznb47JPlajwnQQIywY6ta6EVfzrrV0U1XCAQWKcTMXIwAgRFCSUECJ3jihBmnBWFDKSEFltTAsggNMjGChf+bNnFGsLFKB/a0IONuMUkiMx27EzdbPrZ5glgIKbKwuBYoaJAZKIqQLCqKRFhahwfuaviwCxDDjd0t3RfQG431iPHfOmx3f5sDxUTLBHiX9NrWem7h/ToXXY7f+NeZjx0YxBF8rvs4x/eIRuFkRGD3XRFKsNWrxMdWkmOmnw0zERdmoJQdqNdk2i3JZBnZtF0ySGz+PCtk5S54VIjfcoiIuzikt1IZSR8nzNs+mJ+o+CuDKq0H5tUplEtJzRMY8GZEbimCZ05NyOi+LA3og3UFuobCUSTALBqoV8qTIjRV51a7KQnVev3f0t0WleXxfo7tNJEX1SNWUi6N3iAiK12gk134YCK0/+vPT5USrRl2KZV1rFA5vKETqVpWaUZ0Nl4ZRMCFS4lTeU/hF4FqKnKJ4uAKqirYigDZEVyS6yAo9B3i3++vt2uHfCVtaOjrkrkuLcgcSaTGhq2SikKTU32juGRXGxmkncAuiuRMZ4i8rXCSie7M121sQedFXyqhk3+0X1qJafl5G+1I1JZaUNuqj7ZVWc+P81F6liPqv1ddlaaheAkwcW2z5ur5QF8Icfbbb9Uc0xvd015rPnvjGLU+uHZw+qXoTq9P7Nu/Ls+ic6mc83ZrpfV21J77cmuu+V50gG+LEQr/IiESfIDvfrwZRQDqmj4wPxvMBuZ/aH2yPjLgqDOpJPe3N37p6pn2h1RUOs8IKOfwH1IjYQI7lPrMo6+rYFa1SumzYX0z73Tu2FNxmO2RWzsGAGiTbTdqv9wh4BDwCHoGdhYAnLHbW+fSz8Qh4BDwCL4WAedljIMcYfTECIttMXfM2wrw/o/b9Y+UAQzpGfNI1YQz/UTWIgCfVIChIr0QfVrAQJcYiCqqpkowYYWxGNvCJ0sIxzNvKIheqHstVL6yqksM2lkMbpRMiAoWIcVGXgk+ULggWlLDn1CAhjLhg/lsjLYyAwFBPn1YMvDqXajorm4+tAyMWqwEx/vPSh21HpApkEAvjRgmzIuNElXBc1vGOZiw2nqpnmaXfog8jloz0wBONfTmfVhwcHI2wQflFAYVwguyZd/l67MJ64dYespRhnBeuDSIyKgXat07J/+0RuHEQeBGjaiGD7CjdzTAt+pvd4SCKwudkpAxbjYQ0UFNpVjT0QNB9VTa0errfT2uKAliKk+gp5fUvZIzZSEJ3qjdIF+Wpvb45SPMPv/Wwj664/PQHvX6aiLBo4OUu8qcho9l+YXef/j4wcpl1Jd6z2KY6WI31GlBaruCUolf0jC67SgiigIwylzG5oBC3j7J4be6vF7l3bmjj4A+/40j+uSeX0unJ+lAX3PRgkNZELPY6vTRrd9OOoqNuUYyI7t9gSROJlDNKBb2CUNfbWtZN13VJKsKnXG82koFqYvhowtfmcrtRjsK1jZxIfYaLyyglUe7ytK86FNmoPhuxx2UeIlMhn11mO2FzRSpsiJwYxEm+T6mXJmut4aausp7qXeAQsjx7eH1C0RiBoi02nvzs3bFqPHya4tv6zYz4HBn5ERmP9dvZZzD2f9c1gofcplouQUtkyeTa6dnTGtP+1ednkYFrRREcq7eG67e+7fQbk+awEdfzvn5nDDjqIDsiR98KImr0RV05GxeyrOkSyM38RqrTk0qN1brzLzy3fOyhOz+/uTSF/Il+wLx4/1rEyFXvM92L9bjWKKIkWcgG3aMX00KNFuRjUr0iOyOb+sUj4BHwCHgEdgkCnrDYJSfaT9Mj4BHYvQhUCm4Dgnnco0BYzQYl3f2mzP+niFDA+E34Nl5VKCVWLA+lBOMcUQEYvDF0G+FhBbTZvurRb6BzHBQtS7Fk40AxM09a9rUoAiMz+KySCuxnx2I9ylU1WgNlkugA+sTjC9KCbVC8UPIsQsGiIujPSATGZ+mlOMbvq6HYoXBWPemsYHW1Bgb70Q8kAESCYUX/1agQyAlwoz++H1NDOYQEYjvWf0qNOhaWOgsSwgiTquHISAzW8R0lDoUOrzfOEZgzD8PSIl8YI9tCRKCMUteDVFBLrvvkAad6hwx6vL8RJN6IMwbFf9zUCIyeJ4qOyGVU39i3Z+JYluaTSu00lNf1jDLfHKzHUaqNljbag1BkhurxuqUojFwQuaEM6E+Lt1iRd3ZH+w9FcniyYsvlcGxh2UFUCKuGolj2NxvxvXESHxVJNNnppjNZnu1R9ERThZGHF1OUB7mMy/cK92kZpwrt1Kwl4aqiXx4V6ZHLiGzvh5v6wvODv74ItLsK4ZluDkV0tXUdne0P0tn+IKt3e6rcq3eprqkijoI81XVYi8t+rMLbaVqe17ZP1BvJKYVYrA71XBi/a6/vYH3vNxICPF+QY3kafVLtQwwOwiIbDpyM5q04qStSoo48ZRENyENWE2wk+8lIT0RFKaJiTuQF8hcyJ9EJGNqfEhEwHUTl2xSB8eibP/Tkwvln9v7Gs185+gkRCe/T7z827o9aaz+ptp1tBmKF416LA4mlb4UQQdZsqJbGf6lPxbYFk43p/htm5jsdFcueVUTIvo2lqV5zqv+F5kx/RWMlYhe5mbHg8GMyMsQDWNnC3/yGrEo7pfYHIh3SuKYq473aMyJFjo7HS9SzyZbbyZOifoA+m8rT4dEik0j+AmGBzEr6Ls4T+FhkTGU4/qtHwCPgEfAI7EQEPGGxE8+qn5NHwCPgEdgeARQRIiMw6OPFj0I/dL3nWq5/kr9RCDBiQ1iYsRsFiYYxHIWFVEPkj8D4boZwohi2kguMwggM3jdVA5+REVZbAWXG3km2jyk2VUN9lWBgLFaED7KC3LuQIJAMNnbGUE3dZMSARWhY+iMULgz0bEsfbxnjZOMygsL+tmgSM+rbGNnXjm1REIYL5APpmowoul3fOR+jwrQMVAuh+W9S4zjV+hVVJc+OZXiBA1EV9EX0y1E1SCX63IqlpeWCKIGYQrledvGcFNOw7vK2kVAcm/PNWC1yZDxE/+ERuPkQGBcVHuUNV5FdogA2lW38GZETt040ay0Z2utKANVIatFiFAeLNeW7n5LXtgiOTC7bqlsRLrc7WQdDulrx9IkL1efSzQfIdRixDMdBsx6HKqJNke15pc/ao6xbtcEwq2O0U8qeGZfmpdZPCe/Jfqos70E4yBrxHhFAdzTKfJ8rwxPC+szoAT3INhVlMfB1Qq7DydpBXRJlodRQQ9WzuKDIqa6ICe7TeREVekcG67PTjZaiL+K1tV6ktGQ91a+YrifBinLAnVNk1UYQR9n6Zn9E8G9JjTVC6UZMh7WDTt/rNpVxHQsM+tQ6Q94h79mc0tNR+Nll/Z4rJ2aQi6vRvZARyM2WZrOvNEgrsq0vyUCfRhcJC+RC+iKtEkQEstiUyIzvqV+r5r0AACAASURBVE8M3vGGt5x5UCTHs0999u59IhKQtZBDcVR5MRKcVKY4mlzLgmOKvJBGcqA5HY1kVY2x35gYFFN723cPu0msehxhc6aXTs53Vw5NnvtaFJWkvXpY2/5IZd6QJaQsJYqC9x7ECf0idyJ3I3PT/wOaz8NLx+fbnbUmOgHjQIZE9n2xyAh+y8RZdwbdzVvTXlvRLZdxEhA/C2rPqF1L7Y9rwchv4xHwCHgEPAI3AQKesLgJTpIfokfAI+AReBURQIHAqI7ygxcWipJi37sb8j1ekZbQl78YBnMUJzOYmxca27I/nvx4V/2K2g+pfUANZcVSOpmRnGFXjXpmdMcoTjQHRnMUHytUjVJTXaqpmKrkhRELvMOYC6QFCs1bx/1ZTQuOjXJZXdjHojSMrKBvmyvjQTFDMeI4jBHFlG0hNWy7anom+jOvN/qy7aokg83lAf0OAWDRJewHFqxDqWW8fAcTSBgjWwxHS+1kUSIWRQEJBVnBOUW53BodYaQJn/SNIn0RxyI/47KNTTcY2QhpFmnCNcLfVmBRX/3iEbixEbiawVEjrt6LubI5RWeXNpyMm8uKBKjJkM591JPHv1JouI1WPYn0GcvoyfNgWUbOpc121pYDKKljhvtaE+Xf/OA9nrCoXArCPVBBc1VbjfRMo1CzC0Q4UGD7kIzFdyopz7yIiLqMyQNFrygKI6HeQKByAi6Oo8M6F41uP3u228uKWi2eC8Oi22omPMv94hF4SQQowK2NRh7fuubOUhel1axN61rbo8iL2UE/q4dxGHY7ww3lhLrAtTXMnerRFP1hmpv390sex2+w4xDg3D+nBmGAXDZayjx16aCrKIteGNcR/y5bkDlHzh9RXJyfv201nD24IdG5NLsKMhZyLjLc96tZbQg6WhNx0d5/x4XkxDfesNZdbar+SsDvbGtLNeUnfZl8aZEGRMdeMagtYySqAVmU7czhJpBEnmwsTq2lw3hGhbGz/mYj1NsxUcqrt07vmzg5ubc91DzYx4iB4/oORm9T+y21/0/tb6ohHxKFjPPTqM6Z5nFY/Z19/tHDA0WPoBsQZQKpgXyObHs1pyZ2HekBiq5YHnbWp1R0e7zppRkxF4sc9u/dLSfa/+kR8Ah4BHYyAp6w2Mln18/NI+AR8AhcicDvatX/oGZeY3iXoZxIEZIeULSXXDhjBbJJD2X1KXhfYDyyPL4oDZ9Qe7uaGcer75Rq+iXzREOBQ4H6jBrh4xjC362GMobCgsHePNlsH2ZQrRtBv3i38cnx8OxinBQiRGlC6WNsVULBFBxT2iyM3YqCWwopcGCMjIvoB46D5sS4+LR0TkYWWGg6nxZVYeRHNcKD45nnHMegQRiALV59kBILau9RQzGEwOA3I3Lo3xRWU/iMuGAO9MFYIXysrofVvqgSFbYPSu+jahRDlCtbd8YNF/tu+Q857zSuCSOSwJRrxi8egZ2AgD2XhiqqLTu5MlDk5QUZLdenJuqnREi8oZFELd004aYMm7KrD5XWaEUG91y2zo6M6usKuRheWOv6dFBbrgYiWD720PFCkRVgLCNYoCw75YSCUQ6p9napehZD1Q9QSpKis9lVvh6FsKgWSI2EWxTpFnHRTPN8XvvPNRrxZBKH0zI8Q8BGvpbFTrj1ru8cqHWi66Q4u7TpDsxPrg/SLBwO5YCh96hqU5xXjrdkupYo51i8oeieNIoipYkq9a6LetzPXL/Xd4S+9xsRgXGUBdcJMunjau9knKpzoicTATqy8Yu9VmrV6vAhDGTYL5bmblk7v/+O5aQ+OcgURUYKJhbSKuE4QhQCRn0M7shVOMMgo75NURmH7v6e41945BNv/N18GP2c1llhbeRMZDRzvIHMsAVZ0ZxcLKrharAiMyLfQRZQX8KciMTdBXE2jCY2lyZbIiycIj1OtpcnStXXmDp47/nbNE1LbYoMyZgZL7Il8igkBWmzkDl5NkMiMNZ19Xu6v1mPlhf23KZC34t5GpHqiuMSgfFS5AoYd5WzbTkb9B+opIKyuSEXQxKhP/jFI+AR8Ah4BHYRAp6w2EUn20/VI+AR8AgIAauvgGEeQzoKCAqFPLpUWnZ4/h4Xz2AwR4EjksLC2wEPYzaeXygNKGN/Sw1lhXVmDN9qyKuG0tMHBnCiAf6NGu+gf6H242p/WY1oBvMKQ2mqGtv5znGsXgR9sQ3jRBki1y5/EzKPcmNeZXw3ooJ9bKkSAChfeH8xBwz1YHNIDQUJhY0+UdggeVguGuQuLvRdjQThO+O0aJOv6vu7xuvYHvz5HWUUooU+jQgBS4gK8yar1v3YLmrFImGYA55w1MVAUUSZvVqEBzgyNup7MI7cDc/d5oK0cGGN4/M75wEMaNVIm4sz9otH4AZGYJv0LaR6sfsh0DY5kRgyXG6qbchIE6suRdyox51OP51WIe5chnMiBQathtxQlTsmicKVpdVOT2mPyp//8H2esLj6NSACqIhEBrVE7syoVkUoC1mYxIEwLPVTkYuk6Csxyaw+p5Syh9RcK3roiD0K5ikWIo/4syp6rmiWINEO7f4wW1QUjPeAv4HvuRtlaOMC7TnEBe8/3dMd3a9pTReboqgCpYxySS3Je700JdXb+QvtUd0KT1bcKGfwdRsHsg+y00Nq96pN6hnlinToSE9Ua066IL6idEQswmIQxfnZMC4eV1QCci3yshWZRiZFVsawj3yGPMc7iM+Bvm3OHV5LJue6S+vnp4hAMMLCInqRbatRF4BjKU+RS01u3Spjsx1yHDIr47ko512UPUeR0CIXFrTFA9kgUQRJohSvZSdpZPXeZuPuibneokiMh9RIiwrhYlHFyMH3qaEv4MSDnIq8fLFWXKmC9mGZti9MNEVW4Mhk71vkySU1ZHfrizFWF/Ha2bHO6vmoyK6aOerT2vgxjiOCyROLW9Hzf3sEPAIegR2MwNVecjt4un5qHgGPgEdg1yOAId5SBgGGFYtuubUvbLpsJVaKIBQMlAuULZQD+4RssO8oV/eMf7e6DWbEs8+qwZx+SLNE6P1H5a32ebUH9R1ljoLYeKyxWKSFjY0+zFjFuFG8LMIBpY30SZ9Xw5MMhQrjP5+EotM389hquGd8VU8tSxtlZMO39DvHQrF8ZHxMtFUjZexzPOTLCnezD2O0WhHkMTYFC2XNxoJya5Eg4I1nHvjigWe1RGzstv9lLn7j/dHuUCDx6APDv6NGjRH6uuRVN94WHBkb/fM5dEUWqHZJ4bon+q77FNhD+lTJGHDgmvGLR+CmRmBslByRoJAXkBb6PronlLoIAybPhAsykp9Zb/cXZUg/r42XZHBflLf/oqIC+vcc3ZuLrPAFP7e/EkIRQIWe7ZnwCjv9YSimoqGolGmtL6Mg6Cot1IEgCo6EIU7MKoSsmIt+P72g732tmxTmt6qLPanCLUR8qN5IvvW5d1Nfh37w1x+BMXFRkr5N1x2RUcgKyAbtXi/rqih8X5EYKc8AT1Zc//Nxox+BKAuNEaP6Z9U+zniJqqD4dtrvuvxyI/qovI6aHHqCY6r/sDzo1I4pQuFLWmfpm5CZMOgjn0FGfEUNudLql+EM0omS4sCtbzu1WGumT0F+yOCvtFIj8Rl5DjkMUmLrAukAEYGz0XZ2HIv0ZV/kyKqDKgeAZDiuKa5R11oEhjJghcPV5+emFR2hlEwhciApRpHXiTph7AtqyNsUv8YhCHkWeZV7a6HIw2+XRbAhwqIvwgInneoCiUP9NuTJqy1Laa/71bS7+aYX6mxf2uw/6RsF0cHS16/YBkC/2iPgEfAI7FQEfITFTj2zfl4eAY+AR+DqCKAAYbSDZECR4hPlS9mcv5y59lMd17rvnAtn2QbvKhYUJBQjlC3z1MK4hxf/D6qhmLFczfPJjOYY1SnyTHj8YSmD9PnDaqRBotA0f2NkxysMBcgKRls6JYucsDoLjBuigdRG7Ic3G+tQoigMiGKEogVhACFgZIH1Z7UfzPjI3Bg/x2YdChlpoVCSGDfjtPzGbEeztFU2b4tGAE++M+dPqTFPcGcc9LE1dRbzID+wRZTo6xXLyGN0vLZqwGPcEDMor6QAYPyQSS/kLH5hrBYJQuQMtTSecEWv5fJO5DqPgKFFyzC+anqtqynNVxujX+cRuBkQGEVIibQoZawsxpEXKjc/pGXKhT9UHYYwzUTm6VZV9EUxN92klWND6BVzlEe30283w9yv6xhViDzfPz/R3zs7sS6v9lVFR7SVcmsjjBysQ6kUUVkikkKkUNrO8lSO75mMyk3VE2iOnOCDIFRBAadsPpmiKjoqzp0qtY/GXK9GmF3XOfjOdwYCRlrsjNn4WbwGCPCgIUoV5xfaEQiLXFEWhWoqEG0RRFFbL4RTekwhI07KsD+9fm46Ut2G75uc75w4Ovc8aaGQl5CfLJoWGXVBDQcfSDPkU2TvprYND9y1dDSuZ4+dffIAcuC+YS853V6e/Lr6vjPPoj2SCj/8Hcwd8uWvqlWjjJFbkbORa1c0ho+IKGkpSuSCMvedjGq5MmEVyJBEm+AEYxEakBPMC7kfWXJEAKqNHInUB+NHhgRD5HWcfagLgn5gRAO4IqtethRZ9ql+e+0WMUQiNq5QI5Bp6eNaC45/B3D5XT0CHgGPgEfgRkPAExY32hnx4/EIeAQ8AtcXgTeq+wU1lA6UABQnNISey3uZi8UTrH+x7uaxsY8WlBG2w+PKaimgQFj9BksbhEK0nVGJ/iEAvlcNZQ2Sg7+JKsDIzn78TZ/0g+KD0R+FDyWSfVhntSQw+qMAYahHcSKE3wgV1kE0WBon0lthSbT3HdvR6MsiKmzcpmixj3ncUYAcBZT5V+tiGPFRra9BhAJEDkob+ZAhKyA6+M6YmIsRLni4sTAOlquRPWxbJR4scqO6Pb9DLKEEVscJfpAZ1fc8Y2UMYMk4513/6ZobnF5xi79rRb8vFmG/OC7WLahxzfjFI7BTEDDyj0iLaBxp4cbFukty4GsZE5ntQEb40b25TaqpESaerHjh0oD4mZ1qdqdatfZgmJ0VOXFc6Z6OKCXUnIqdz4iAyJI4HoZBqUCMcJTijyiMLMvb9UR1znNI3XJKURZKCVXmqnVhBPFOuf78PDwCHoEbDwGeM8ia1Bf7stpPXYqy6HVkS1f0g8LD9ND6VtyYaOhzQlJbt7MycVsYlqq9U+5RhMFCoLpI2peXCLUneI8QXYC8jWz6oBpkABESyGMY+u+cv3WlNXd4va3IhEJtqt+pza6dmfnYqUcPv3fQrn1YERCvFK2PaEeTLRmTpVpFJv6gyIqzOn45ubczKhou8mSxMdU/oPXzOuZAn8j/jH0UfaiG3EpaKOROIpvRDZjnIfrRkZ7XfsjByN+W3pSxI4viPHRFXi1+VATLlFJBaZ5XnSbEyufAz6eDeqWXgd/PI+AR8AjcvAh4wuLmPXd+5B4Bj4BH4GUhUH5qZISmLgO5afGMQplCsUAJQZmaccf/6Sl39y9jXH9Yje353dIbobBAMrAe4zjGfFO8qqqGaVfViAEUHAgIUiGh0BFpgaLDsa1OhuXkZWwoQhjXjQDgO2PEOM84rDj2W8djQamyuhEc56gaOW/fMe7DyA4jGMxrzCI3ULIYI55nREKQpsrSUf2ovqO4kU+4SiAY0VGdL2QKf5P+irRUEAnUlMD4z/78xruXsfJ5tfRZ1X6ruFZJEsMWfEZ5idXAzFJXWURJdX8jJcCR5WnXe/5+t/Sf8ZqDxGA9OIEvuNAvyvUjunamgh8cKeF+8QjctAiQ/sWICU1iRF5apMV2tS9u2sm+DgMH31//xJPiHopepzfcJMoijIKOvq+JiJiMAteQ3a9s1KJNFTIv8yxvitRQip6oLWPVam+Q6s98ueyVG61mUChXSbHRyYqZKQtuex0m5Q/pEfAI7HgEMIa/830/g4yE7Mu74ads0oPOhozqqZvce6hVFsWH9Fwihd1dMs5fSAfxY6r94Gqt4VH9jQMQsiUpoZD3MNoj5z6vhiPLXxn3iYzFNiNHIKL4VDMiUhMz4rLGdP99rZneF2YObnz1W394/69lw/jntd3WemnXek5IdYVchzOKOeywr2TeQPXLyvVac5gqymO2u97MJvZ0NySlNkS7RCophIyKDEmKKmR2HsTImBAeyODghbx6Mu3Hf752duaQok2Qna8WSXFVskKk0DAIw7cokqWux/3WOf2WVnxijKlPB3WtZ9xv5xHwCHgEdhACnrDYQSfTT8Uj4BHwCLwEAigrvzdWQFCiUCDIR4uxmt+6rvNo263+2Wfd3AcmlEwXpQOFC6UKgzgKmNV/QPnB0F2NMLAUSQzDjO5WcwIDOv2g5KDsUHAakoB98Oi3VEmQFmzLeiIT2AdSwyIvMNDTB8SCRQpAYpgXrhUZZKykmoK0IEKAcZsxn20tQoR54cH17nGfz+qT/hiTFd8mhRIFGenPlD4jDIysME2L/eiT8UHuEFLPfMCqGqFRVd6sLyMX7NMICo5B/0ZyVI/Nb2BH39UoFyNbLJ0X+4A7/fD9IdUqOeLC+jm38kmICo5lJBHXBJhZOqzfH+OlD794BG5uBMakhT2fRqndxmmh7B6+qp/ni0VY3NyIvLqjV4RKMdmqDUQyLE626qqh7SZURLvfbMWkhQoUOcGztyZDVUMkxbo8lTuKpEj1vSZDYMeFQV/lLqgp0tdvqnBR5tul4np1R+578wh4BHY5AsiXyKDIbqT03FPkErvEKEQqup3nqas1JnFCsbRGc4qqCGXoXzx7bP9j9clBPntoY7/qUODoYalIkV+RpZD5SF2KTGxpjkymHj0T1ZYkOXcDV8b1ieGHFbXw2cn57vH1c1OnRYYgl75cuw1yHXPi2PSPM5ClW9XXspvUxRpP9zfjWtZQGqojg24tbU710zAuiYhGT2D7+9U4PnKsOftQpwJy54wkyq9kg3hW6awEV4izC45ROOxYzTvIjqsuSrvVV+2KTpFWy8pd2pRjHR33dwWbsV2ffr1HwCPgEfAI7BwEzNC0c2bkZ+IR8Ah4BDwCV0Vg7CGP8oRBGo8vDPK8B/BcwtCPQjDr+s8eULZxS8lEHQiUK/5G4TFjPMfAAM6+RhaYMbwav8736t/sjxcaRIQpfvRryoh5bqHgMSYIAn5jvChCRDpgoGc966pGfdah4KCcYainXyI6IA9su0vpYLTOSBQiRT6rhoL1h+OxMWbGyDG/oUaNCfqrRlMw7+qcOQa/sw8eae9UgwzBww3ip0pM8N3qZxghYUZU/TRaqhEqbFuN7rDUUhyTeRsxwX70Y9vbcfi0HMCcM+GSPeee/Ucoli+c+4vn8yJ5dRFfrpV5XTvbFUu0sfpPj8BNgwCkBfUrxveJkao2fntmVT9vmrm93gMFW6WFSmenGm1FUiyrHMgzk83asgqXLydJeF5OtGd7fVmnynJTD6Ver5/lm52BS/MijmtxONVM1uIoOJWmRWc4zPoqiO6LnL/eJ9Uf3yOwCxAYpxxCPmWx2mzy7chcOuy5QvV19NyqIoGsJKLVPb/y/NzEsc/fGfXbdVKLUr8B4sNkOgz/b1dDVqMD5CwIAGRZnm/IliyWPgo5+QGlmfpgc7qXqpdXWkeM/iFFcO7hGMjGyHYsyNhrSSM93ZgarIu0qE3Ode8U2TJPbQ01i4Ze0HbIsCzMA1mYPpkH/e0rXfCmQad+8vwz+85pLeQGaVqZH2TH1W1NZan0UcVTiqxY664th0VxBR8BOYLeQbTyqk8HNT4D/sMj4BHwCOwyBDxhsctOuJ+uR8AjsOsRwGsMJepbahjkSQ+FMoQxGwVtrzv/O4Vb+h08zJ5QI9USigMKFkoU2y2oYSC3PB1mcK9qclVjuxn5IQ5MeUKRYSyQBJZ2CuM5CgpFCjGQ2zEhFlC4IFusVgO/WcRANbLAojOs3oYRBVUDvpEMXAzMgdB8UkfhFYebF+vwROMTjO4c/w0OZsQ0cqLqqW3jZe4og0RXoBxaqqpq5AT7VQshVkkLxrXVy9uiV4wkYV/GSvSHaXrV49g4wZMF0ulJNbC9mGP45C8lbvPPUaA5J1bUkGuBa4J5c43QD+fJLx6BHYfAmLgwwtXmVyVYd9ycX4sJgetjzyymqxu9jZWN3kmlevr2MM0fUXssd8VxPVUWVVD7maIoH5Hz8vlWs/bMRCP5aqMeHWvUk6fUjtdq4VmllkqthshrMW5/DI+AR2DXI2CRpV8XEiY/jSSyYa+ttumyYX9ZkV84pSDfITP9kCItfmDQqV1I+4nS2wXUeSCKmAW5F1nVSAlkN2Qui5bg961LS318WhELMuY36zr2gjZA3qvKrtd6opDtTNZEPra6aYpyCw4rlVOgNkr7Gib5pCIuAj2fkXXZDpmRcSIDI3/zHXmdOh+/qYZc2dPcVzorrUD1N95Va6Y1kR0Paj3OTvRLpMnWpaNiRZv5cNDurJy/NRv0cBqqLhz/V9Q+qbaghmzrF4+AR8Aj4BHYhQi83NDCXQiRn7JHwCPgEdhRCGCEhgzAII8HFR5SeEw9pYaBHW+mdbf2uVl38Gcw2P+Z2k+qoWyhyKE0obCwH3+bx1jV+3+rsb1q1LfC1BAIKCWQBRS5pj/z/mIcFz3XXvBGI+cvv3M8FCD6ZJtqmqet0Q9GZJixH6WnSm6g/FmECf2izP1tNQovghHkCCmlIDIgIxgv0QijNDJqLBaxYX2xL6QACimplv6SGgqjERxbsdkOq2q0RZX8sbmAPefnlvE4OC+Wb5hVlu+YbSyShvPN/uD9q+7Zf/IhfYLJghoh+0RT4Bn3NTXm++tqEBdEWvjFI7BjEajUttga5cScr5oiaseC8epNrDx5dr1/aO/kBaV8Kuq1cD0K3UoURXo2ljIEBoWIiguNRnGw2UiSLM3PDAf5YtgITigCY7Gv6ApFZ2Scm1dvSL4nj4BHwCPwogggEyEDfVTNikWHSl2ktFCxi2tNFd9OkO9s+cHxl6+JrPjIyW8ceeq+73/mpCIXKNyNIwzOP9UFGczIDNab7FjdZo/eOke1Yjqq5SsiFv5U3zHqI8O9qrabtF9788qpuTPN6UFZa6X9Ig9y1R2akQQJkUIaVJx+IG6QD7+qhlyMHEzECLI4svy7Z4+sf7DfqSfDbtK5cHJPt79Zv0PrmSuyNJ+QNqNFdUCWht3NR9tLp9+fpymlii4DSH98QY36GM+x+bht3cb/7RHwCHgEPAK7AIFX9aW3C/DyU/QIeAQ8Ajc7ApZfFiUDwzp5aqnbwPsAT7Hb1Tbdyme/5IpsTpoZiglREBjtUVRQUFA8MOxhDMeIj1F7u3RGZty3lEQWGWGEBUZ9jOsoQ29WQ7nBa4s+0WIwtvM73l1GaDBWGsdknRm0TLGpkgPVSAiLYtAulwgPxmH9cTzmyOeCGvU+CIEnioGaDkY8WDomm5uRJ/wNgWBpsqwQNjgZ0WDH5rP6vRoBwv6Wa9jSUFlqJyNcmDfn0opr81nFwfoz4odPyCjm+qR79G98Tp/U7SBtFYop557fuBbA/iE1zgP4Q474xSOwoxEY16jwxvFX6SwbCXR2uT04emT2gh6SQxneVMeiXJftbzktsnkREqMoMZEVNaUVWRmk2QWlk1pRRIaSSuWDX/jI/T5v+at0Pnw3HgGPwDUhgDyHLITsR82JkDRQpIVSJMAoyiJpThRRXNuapeKQJLB70kFySHUc/iQug28p0oDUUB9UI0LB6l4gD9KQ36wm2taBtSShfr9Wnm3N9mY2zk8/nQ0ji641BxZzlmFfIiEw8BMVgYxuhIhFSmw7cREUZxUd8Y3lhT2z1BFStEVHdTiOqwA4RAv9IUsil0NWUFcOefHHxnMCg+PaL1Hh7vl9Ry88sbww/3XVw5gOgpr6C3i+Ezltcv9oHEWetjqr59+apQOln73ilYvc/K/GGC3o08uf2549/4NHwCPgEdj5CHjCYuefYz9Dj4BHwCNwCQHVIuiWn3K5Pgf6xIBN6DoKAd5beN5DGlxwvWP3utP/54PuDf8dRMV3q1ktCZQiSAwzpFfTGo10ETVbZwZ9M/Cj+KAAVesvoMxgfEc5tILbKEccF8URwz0kgPWLgmRh6ShmFiLP+qoCZ15r1VRKVWLBCgfyO3NCoSLtFIok/ZrnGOmRUNBQooxEoZ9qTYmt6a9QFq1/iASLFDFyBJyqiymurKMv5scxDSdL7wROZsBjO4tuYT9bj4JoJEZVsWV+jJ9z/Mfu/Ee/S59E1nDuIWLIu0y0C2H8jJdrA6KGvoa6VpyuGb94BDwCHoFrRmAcHVGqqPnw7tvm11Rwu5dmRV0J0msiK1SMOwjkzdtVkW1Xq0VBlufd1Y1uf3Wjn2pfnwbkmpH2G3oEPAKvEgLITcign1fDMH8ppdGgu+mipK4a3GEYTSQDfUE+suUWGejdxvmpTaWGWlZqJfn7FE+LtHhAGyBvbV1eNPWg0ixtFFn4qGpjRCJAfn48DggI5EOr14bMjAx9Wg0ZmnpryPREgDA25NmrRXBUx3JIx3nv6pmZVhQX7vAbzx0Uh4Dsx/iIrEA2JOqZiAr0A5OjqWsRS2LdV2TRilbWkmY6HyXZWlzPDk3Mdz+b9pIjirj4gHBBnieSYq3M89VBe2OjSNO3XoWsYLPfVsOBCbmc8+CdCK68dvwaj4BHwCOwaxDwhMWuOdV+oh4Bj4BH4BICVsT041qD0fpH1DCaEzmBwoOisN8d+8VAhAUFCDGCsw8GJJQiU4JQJFiHQsQ25i3GeuoeQE6wP/tAYvDO4RMjuUVVYNzn2BjLMaqjHHEsPPutYCBGdlMaMa4TlYFB346PId8iKWxuVe+3rZEVFpnAfiwodvSPMmg1MAjlRyFjfqM8vWoY/FmqKaEs8sGKVYOFFVFkDJaayZQ8I1Wq6asgCNjfCmezjaV3su2qabUYg623bU0pNQWaMTA/UlShvDI31v2Z2h+o/RfjeRBRwTkigoXxQk5RSsoI1AAAIABJREFUePzjEBRjcssrjOMT7z88Ah6Bl4/AmLjgWZp97KHjg8EwC9Is3wjDoJhq1IuV9W6w2RkGtSQqICte/hFu/D1E2rzYIKvvg6tuN44AuvEn6kfoEbiJEVBx5+Kd7/sZ5FnSpBJpiow8Woosdf32qiIsRqJglay4NOMsjWZEMjRaM/3ZMM6RgYnOrS7IXERcWA24K9ASWfF8b6Ox8Oif3newt954jwz+yNZWsw3516KakRmppYFcjMPNB9SQZW1syHQQL6R24rlKQ3amD8iIUboq9T+XDWK3cmrWTe3bnJrav3mgyMOuCnAjQ9I30SEcE4IEeRyHFpbbFRm3R9vtV72NXGTNnIpv3zc535kWYdMScXPHhZNztWFXZTgkRZZZNui3104NOpvvu2LSF1cQkcIYOR6pSH2E3TZA+dUeAY+AR2C3IOAJi91ypv08PQIeAY/AGAEZokeeq/rMZZAmWuKYGooPnll4UhH6jXJyrzv+j7/h7vhneDuh+BAeb0QBf1sdBQzaKDUoQKxDyWE7FA/L34viYREBRibgrcX2HItPPMXw7HrruA/2QQlD+aKh6N2jxrvLiAWL5jAiwN5r9jdjgBCwY1pYPYQKhnwUUyNRrBghiiHjwSuMdFgYk8jju1VBNUO+kTEoc+Bg0RXVVFOMw0gI9oNIoE8rlK2vl42x+rcpbWxbfW/TD8euppOywuiMgwWyCAIK5RsFMHafDlDAqVUB7kSw4DlHH6QV4HOWa4Od7VoZ9+U/PAIeAY/AtgjIKB9sV3PCDPYqom2RE/ZZ9TS+lK98q4H/ZjfYv8T4iUKxdH8WWeevNI+AR+D1QWBbQ7lM7m7QWXNhFLm4MTFQkNhlcqHIhvrS8b13HrxnMY/ifBDExb/VFH5UjRScLDjnbLdsiDz47cXje59R+x7VhKAGGs8F5DfkVWRr5EYWZFrkY+RW6mXgYIO8x9hxBLLnCcZ/asAhzxpJgtyPU5At/D4v0sGdfvzQjMiKu0U6PD5/6+qkUkNBdiBDIysio9MCjXNKkRkb2TAedlebk5vLE6pDHi42pgbTSl+lAtzhXu17oTHVf6SvJLMa+oclSU9FcfL2KEmCbHCFHwwrqLH3oNoT4+N5wqJykvxXj4BHwCOwGxHwhMVuPOt+zh4Bj4BH4AUE8Kb/b8fKDNEVGLpRgIgqOOSe++cXRFh8Wt9/Rg0FCCMTRn7z8MIQj8fVUTWLKIC4QCGyaAeM/5bCiCNb/QkMVWxnyhh9HVbDmM84IDjoC6UFhQmyguNbZEW1CDbrjJwwTYj+2Y9x0A+Ge1OAWIcBn8gJlDyOxXeLArFi3hA4pthZlIOldqoeh3lBdNCHpb0ygoLtbXxGZhDRQD5gi9zg+CiWhmGVnNiaEqpaL8SiPQwTfgM7lFfmjJL7nBopAyCD8KwjuRNKM+eYsZIGijmCL8oo14RfPAIeAY/Ay0YA0oKdthIXVzHY2/NzV0RwXUOEhUXJmW7Gu4J1uwKfl32h+R08AtcJgXGUBTLU/zWWoX5Sn5eICaU0cspl55IsO1OfmDqn7xAHpFVlqXXWmh9ShMSX6hPDN+hv7mfkL1uQo5G3zKnE1iO/nlGkw9Lpxw/Oby5O1fU9Js2UFpyJrrbQ9/eo3a+GQw/yLhEWOM9wDORKGn+P0jJVFo6PDIwsiDw6WjRud+7p/bPT65uHVD+jJ+KCPlmQH39V7c0a03Q+jCZFTKxvLE0tDTu1e2sT6YTSP83FtfyWpDksu6utJ4IgPdGaWQxWTx/cKHN3Mhv23t7vrKsWSH9UE2TLgp7xoNoX1ZBTTX/Yup3/2yPgEfAIeAR2EQKesNhFJ9tP1SPgEfAIXAUBFAQ8v0gLBQHAgvKFIkNExQfcZ5KPuR9I0S5QeiArjo63swgCakxgVDElDCM829FQ+izlErtVvWkxlqO83aVGWDvNoh0wtOMNxt94dlWjM+iPaAAIAsZgqZpQrCyywgz+KIGsg6ywaA76Y34Y9CEJUNYYF8ewBWUJ8gDigv45jqWyqqZ5quwy+sqYjWBgDJbmif3B5+tqKJREnuBFxjEYD/P93kpnRnZU+7eaFKyr4sh3Ix8YN+OE+OE7nncofxzvSffNH2aupA3gXD+thkINNvzNWB5We7B6UP99dyDwjee5va9Y7Fq2Hy55wG/d8u1v4Hb0y25GYFxoe5SeTwb6Yrtoi92M0UvM3Qho3juWbtHSDHpvY3/heAReOwSQoxbU/oUaMu371Ujl5PJ04Pobq6Q5uj1pNM+GVOIJXhDJyjzc11ltzal4NZHGEALIyMii9Insyn1erWtBvrgzis7oKo3StIiKpxTtgAx3rQuOPzicmByL7M1xiMZA7kQWpL8qSUIqUOQ9ZNYPqo1SpGoMrrfedBNz3ZaKcddFWpxQyif6AQP0BG1XzuZp1Om3GxfCsLxl+uDmfNaPa921ZrMxOchEcqzFtbRIe+W06lnsaUw2ji09pwpFaery4UDHyNUue5whvyKP41yDw5InK671zPvtPAIeAY/ADkfAExY7/AT76XkEPAIegRdDYFyEG82B3LEoVRjwMV5TKBBv+7oS9064vP/nLmrgxTVS2LSgGFn6J4z/eG9BGJBqCSUNIziGftZBMBCFYcRGtS4DfaEwodRxXJQo+sWwjuJC9APvKot4YHv6I/IBwmNriiRL/VRNAYXyhkKEssaxGZeRFIyPPjAO0a/VkrBwerY38qDaJ+OoEgj8zWJzM1LDCBTmxvbgS3//Ue1jav9oPC5L7WTzMcMVfZqXrfW9NTUUv5siym9EbrAtyihECBh+y+XdxF34Y3CwuhycY5RQsKC4IddAwTVhk/GfuweBKuEg8oLrx+rCWEF7+7xkTNA+3vt791wi1zpTe3bxLNuR9SiuFYjqdteQEsqe79xfVieKLlifQACNn90WsXfZMG72lFmvBFO/j0fgeiGgKItctSyQhUiZ+lE15FeTf0VaDF3ab7uimL9LbIU5zTCctoiMyY3FqXcfuHP5uApRX1DhbRxDjITEIQh5kDoQVpeir6iFjbSflCqwvao0S4/pt7/4MubGswF52GRUnGJwOMILAZmc8SGTWw04joucjgyIE81n1CBkRlEkRR641dMzX1FKp3Lm0MbJemv4tiAskV3fLyn2rIpsP6lIjNt7m41DirJItH2u9FDl9N52GNWzE3lWrmb9QdjfLBvZINvTW1/6yKBdvqHI9GqA2KGgxQsL0SePqv2uGjIrDjx+8Qh4BDwCHgGPwAgBT1j4C8Ej4BHwCHgEfl8Q/KwaeW+JMkD5gUCw2g8PuOd/+ZPu6D/E0H1UzYpTYzhBCcNzC0O4GfeNyLBaFiggWyMfQL0aJUBaKJQl0hPRL+HteHOxH95dVXcsjPv0bfUr7HiWKqmaaoTt6A9CBeM8Y+E7DeWNcVuaJo5Bn+ZFbv2hBFrKJfvd0mNVCYaqwcmMuzZG5obye4fa76kReUJhb0gZ9qvW7TCvdsPMsGI96zimkRg2HvqmT9ajrDInalOcULuYCuvcv4PIIIqDeaN8Q1RAJHHOwQXSgmvBL7sYAZEVRlRwbdG4drmuuE54Bhj5VmjbUb59T1zs4gtmy9THURaj55SM7Pb8LXd7tMU4gqn6zrvMasc9NE4bxbMbkp2FZ7VF7UH+sN7ep9tGO/mr0SPgEfjOERiTFrwPkdOQFStL6bJ+1/XXLyTh3P4TUVKDILgU8ati2bXuenNuKslXZfhHPoMg4B2K7MU9jHMOUcWpohqOnX9638Mqen3X+vlpakLgzIKzybUuRlTY9jxncOqhJgSpnKhZRqQtzxOeIxa9hawIgQJpAUny96wDkSc/tvTc/JMiK7554O7Fr03va3+/JNVUxEot7ccHFAEyp896f7MxGHZraxOz3SO9dn1z6ZGDT07uWZ4o8vVbhp3ijt5GcGjQzlwUB/J9uoKs+KaO9+/Vjqt9ZYyLj6641rPut/MIeAQ8ArsAga0vuF0wZT9Fj4BHwCPgEagiII96aldgmMTTCUUKjyyMkhhHLobFn/4/9iuGG8Ml21i6J4xSRGGgjKEgYfBG2WBfPLqsbgNKHMqTFZ7m8GasMSICAgGvr/eoYaDBkM7xzHPNjKhmzEfxsnoW9EE4uZEmjIftq7Un+E7YPOQHfaAMQsiwzhYM+4yf341oMNKi6nFuJEGVrKAPm4tFZxjRwW9sa/i9U9/JOwxJcbsaRbCZ81ZvdSMoqkQMc7Z0VVUiBYIHDJgn3yEnOE+M6bxc5truyV/AeLigxjnlN84T55pzznmNxteC4eE/dxECRFV86pFzcac3TPrDrD5M8/pgmE1mWXGwKMp9ajNFOfIU5d7hXuWarUY+7SK0/FRfDAGRE/YsrHr97nbQ7B3Cc9tqFV0iMMZkBe8AsOP5zPuSZ7q924xQtzpLXofb7VeUn/9rgQAyFzLVr6sh715aSGvU31yd621c2KfvEAKjAAIRFO3mdH9NaZPq7ZXWSa2u5lvkvYmzCPLgn4gAeFZG/5PHv37b1NljB25TGqZf1LqXQ1Zw2O0iHZH1PqyGcwzPGktHNUr/pIW54Zxkddcuy9Ok8d+3uTz5j6O4oPg32+UKjji1dm7mk2eePHjs3FMH+ivPzxYXTuzZXDs73e+s1pN8WLy5yNJ39DfK71k/Fx5aeT5UJIrICkVtjBeeZ8inRBn/uRpkBZEVFP6+7Pi2g4ijS5j7Lx4Bj4BHwCOwuxDwERa763z72XoEPAIege0Q+Lh++GtqeDyRWxfjPwZ9lKv73HD5pFv79Ffc3A9997gDFCRLXWGFuIlgoFEvAW9/M9IbcWFFsU0pMfKBLtkGLza8zjDkk4/XaliYJ6kZ6Kteqig5HAeyAaKg6o1q22OYR0FkvBAdfFqkgnmQWyooIyyqxiBL/XQ1L7arzaXaB2O1CA72RxHF4430WpALYIXHHZ53KMP8bkQFuBhZYRgx1yqJwtwW1CxSxAxh4IHRi3Oz6BY/ivca0RVH1VBOzQgGgYN3Hf1yDfhlFyEgI6kRge7YieWokcTN/iBrTbZq5ok5rezcrVoURXhXxlE4U4SuCIOA+5TrkPutLbKDa630kRa76OJ56any3DTjelExyF+x505NZzROrcZ8jcS2FIRGSvDb6B3yI++/11XuH/ACP96nVp2WZ7b1ZdF39i70qdle+nr0W3gEXikCyIdEKzyo9tPVTops6Ibttb1xrXGiPjnbDELXndrX/qIIi7fWmkobNYhxCDq65cBGXj6qaIovPfXQnZP9jcZ/o9oX7788W9I1D7cqE1d3Qo4mgsKeM6R14tkBkWE124j6JW0oaZlIC4r8PVogX+Kacj2VwQG1oVJbUarjjjjJnp49uLFXUSHrmxda3TDM9gz700EYDuu9zezI4jPRkTgJXU+uMPkQsoI0U5eGhcxAVAV4QlxQy22UqlTEhH+OXfMp9xt6BDwCHoHdgYD3ztkd59nP0iPgEfAIvCgC8qz/rDbAcM17AdXC0r/ggb/fFf0jbuGXHnB5D+UCwwmGFwzfeGph3OQT4zmKB8YZwt9RlPAio7EPnxhg8DbDCIPBHgUF5YnvGO7vUsN7+81qFv1QTX1hxnyULosCIUIA4oJjWuHvKmnAONmWMdKXGY+MbLBIDj4tegIF1XKF27uyqhTaOGwb+9xKbtjfHNsiQb49xoB1eLxxLCssXiUjtPpSAW/rh9/NgAWWGI5/TQ1PNXAFA6JVICIwIoeuf+aUe+xnwRPveH7jnNIH59iiNb4+vgY4pl92DwJc281GLZ5dXunuXdsc7FGExZ52Lz0wSPM3hoF7mwwNb+r0sls73fSOTi+NRGg0FHVBMwKS+3xEpFUMtLsHQT/T7RDgecfzhec574vtjGo7GUHmzNx5LhMtaA3DId+5d6wW02X3zziFlpH9PK+tWfRF9Z2zkzH0c/MIvG4IjI3o3Hs4geDUQfrSS0sphiHt91xn+ext/fbqV/Nh75OKtjgpwuLbzZneytzhdZx8iGC1heci9StOigSYOndsf3ft7Mx3q3bF214hWfFi2BhZwTZvUiOitypDIgOa/I7MaJHFoz4Zz7BXc6pXsaz2p1rVUC2LW/bcsvY39tyyMhHG3ZVs0J3orG42Ns6XqnuRTraX1490VwduY1HFu9ckfraD3rAXKED70jBJd/Vnaugc4EBkSurJitftEvcH9gh4BDwCNzQCPsLihj49fnAeAY+AR+A1ReAhHQ3DNsbvd6lBMqCoYVyJ3Mqn3ug631xx0+9hHQZ2DPxmkGGgGMQhDiAH8KLCewpl6OL+F9dbOiIMMShTGF84DsYb9qVP3k1WRLoahcExzHCPsYZxEK1AHl4rqG2RCvRn9ThQNCE/OA7GISMt6I/FCADzCCa1FWQCxlwbR5UwqKazYvzVSBDrs5qH1wgPMEAppJgiOGDIIsLCSIOthAj7VYuAo/JZwW1Ih6fV/kgNjzjGjGGQcYMJfXI+Hncrf4T3HOeTc2Z1Oyy9COeabTn3ftklCIwjK7j+uN/2yG2yIO3TMM1ajXo4l6b5rWVRzpIGLs30f1k8X4vDdrdfFq1Gsj9s6t4Igo1sUPRrSTQThoHl17dnxi5B0k/zRRDgGcMzjOc/z7tdVYB7XAuGdxlkBe+fEWGuZUb3G+8B3kvgQ/pDjHaj96P2yxVpMTLvVUgLf6F5BDwCrxMCGNNVgJt326fVkL1+VO0XbTilrPHpsOc2z52oDyfqF47cn6/tPbo+pdRQhxSRgJPI82pEHRu5Pycy4NH+Zr25emYmK/IQ+Y3nI8/JL6kRDbugxnOC58ertfAMItoYooCaG8ikPIOQl4m04Pgmm+rFH6i4eHghG8TxoFvbLwIGWXFdAnAtSrJGY3K9m/bKyXyY7R/22vNEm1DXo8hyCdkSZy9KyhbJwfcvqOFUZLI5875qGqhXa8K+H4+AR8Aj4BG4uRHwhMXNff786D0CHgGPwKuGgDzsj5WfGqVlItIBJWJB7U41q0mx6Z75h3X31k8uK0kvihfqCAZ0izbAGM5+VRIBIzoKkXnbohixHUoR/VYjOjD8owySK5dt6N/SOpmBnfkasYACSZQBxAhkh0V08G7DGGskg0V2QFaw2DGNSEB5IjqBlEzMhUKIKIqGg4XvW38WUm8pr1DAOAbHrKbqsPHbmFEWmTfHQWmkWLmlsWJbjFZsY2mf+I3twcUIEPBG8cXLb0ENpfOEGoQE68EbXBjzihuc+rI79vd+QN+JfEHxtYLp5GR+oxoYnOHcM0i/7HwEKmmguFYLGU8P5UURi5jYq8874zickKFi8kJvMF1LYtdqxqnYiUkRGuv6/UCShcMsj12WpxvDYd6em2kedEHYUpoorl8ifowA3PlgvoozHKdMosdqlNWlFBk3W9qkcfFtnls8ezDGjd4Du6H49pissGc7ZMWtanXdQ5xf3hO3i7jo6d7Ts7qc0CfvTN4jvH872j/16dVexZvLd+UR+A4RGBfgxsAOoYAseYmwGHUtBqLI8/cOur17l45n//fhN5XHZyXJBpFSql6URdmP+mXIfd3eevOTz3zp9sHG+ak79b5F3uR9zLPh/eOhQiBcjwX5kjFVF45LQ3ZEFh7V0FAKKEWPJPNFETQ1g55qWvxxGBYuG5YPhFH6bGNq+IwiSt5fFOE8REWepa6QILHN8j9pPVHcOPk8p4asX3XsuR5z9X16BDwCHgGPwE2OgCcsbvIT6IfvEfAIeAReZQQ+qv5+QY1CgRjCUVxQ0lBwHnarD97muk9EbuL+gQsjjPRmTIdgwGA+MsaoYRiHQMAwflQNYzm/YZQxQw7b0wfGLH7nncTx8P6iEDVKnhEARjJYFAJaEUZ2KwDM+mp9CjP6mfZkJMbW3N/abXR8vF0hLohaMK9X5sGYjZQxwoLxW8osohaYE/tbNAlKmHmuWUQExIN5HB/Rd/CxWhIocPSD0lqNxrDj0X+VhKF/8ILcgIx4UA1FEGUYTC/mKS6yBXfuP7zH5W3mAFYowqSg4nfOLcfnuJxzv+wCBCpkBddOPYrCmgynB2QwDWtJ2Eqzcr7dHe7N8nxymBbTaVoUeVa4OI76jWZ4VIaL7kan/3S3n55VPYuDeVEuNRrZxkQjCVSynftolNbGG1uv7WLS+ahGVfHM4BlhhcxHEVUUsGa7F6sBwdFuUEKD55wRt1Yv5RIJc20o3ZRbcS55Zk/q/tqnCR+VPXNSRs29+h4GZTmrv+tlUG5EQYDxTu+TsqP7kHeBeRzzzvCLR8AjcIMgMCYtcJJBRv1NtZ/bOrQyL+cXnwn/9uOfSv7BO39i2GpMlbcoyiIRDc2zkHv9lFJBLV04uefbndXWXYquIFqDSFsiMbZbIBE4LtGy12tBruQdbjXhhhrnvn67vrl+bvLY9P71WKmuDriojPWcmkgHbvaZLxY/m/YH+/MsU62KAeFjjI1nGHK9LaR+4pmGbP3l8e/8vRveA9frXPl+PQIeAY/ArkHAExa75lT7iXoEPAIegZdGQJ72JxRlgSEbI/d71SAEUD7wkiUH7oQ7/9Guu/2fodyQygJvMQxsGPAxSKGUYaSnD2o14MXP3xhf+J31KEU0DOcY+jnWKNR8/Dt9so/VmjACwNJD8Ul/71DDmE9BaYoLEmWBQoentxEgjNvIDH29RBoYGYByxfHxDGfskA6ME69YxmAEB79bwUI7PvuxHWPhfco27I+XGvtZKD9jZA7gBGYop7Yf2LIeXCyahHGa4gihYH2Ncv2qMSdLRcUYIZfw4B0ZodUgJWI3PHfWPfe/ggeKMP2zH8e2c8q4JjjnHNAvuwYBrhOuv5ZyPTWUzknREW5flpe6hsp9qk0xncfhHtW1aOR5WaRlkZVZWcTDZJAWWT1w4ZHGVNyX0WKxVYtTERqL/WG20qjHSRSG3CMrFOH2pMWLX08iICxfOM8Tnh/c/9V0eKMIMm3HPV417txMhh6LjGOuPLtuprG/ogdCJbqCd8FhBVWI6Cvv0D12e6B7TU/zVClkMt1vKmZbzgdxpJRspYjm4FgYjkgLroE19bOqe8hHK72is+B38gi8+ggoLRSdIsthfP+dsSz1I9UjYbNP+8HUyW/Gf12Zoibv/b5sozlT9qKkvBDF7nEV5T6giAQ5AWVTpIQSKYC8SyrWrQvHseLYRCZXSYCXOzn6sYhdS9FkMjB98Zzm+QyhMqo7JHJiVZJzLR+k55/7arDWudB89q73DM+lfVe0V4I5ze89a2cHc9lQXV9efMPGifPML6mRDgvZGMyQW31Uxcs9e357j4BHwCOwixHwhMUuPvl+6h4Bj4BHYBsE/r7W/4oaBnKKYGMMR+FBaeq5jS8Frv/csmvecVBRFhjUWY9hBcP4b6lRO4HoBBQWvhNpYd7DHBIDHYZ79rOIAjOiYkQnxRPKFAZ/IjjMC9m2pQ9L+cQnRnka39mGMZsCRr+WOgqjPeOwAuAcA+WKufEdRcq8wzDsE7WAMsl3FvMQ5rsVHGZsEB2kYqKWBuv5Tl80wt7xjuO4Nlarj1ElYMaHuFRk2+ZMX4yJfSwdFGlDwJpIDUgI0naBG+cC8uJeRVU86B7760suX4cwYoGksDEf13c8BDFac679srsQ4DrmWuX+a8uIyvWkmhXuNuWA0PpyejDImiIzYl2EsSvDIlPtzO4gS8VfFK7MI+0zpZoWx9Moz5M4ihWVkR/YOymbbOlEgHAd2j21u5C9xtmOI11GhGwSh800KwLhNh24YHbkgR+4gVobOLO82Op1fzMZfOy5yvPsZhr3NZ7Jq242ImV03kJFIU2MIizKsla4YLrMinrpyk3dRW0xFuIm3GyQB6N3nM6/3g8KdQpdTT9wbbTH9Sx2PMnznYDt9/UIvA4I8EymHgN2FKKI/251DNjvi8x936lHYre8ELmpfcXHRVQ82l4OhvvvLEoV2I4HnWGRp+liEMXmYHO1aZgzD8+D74SwMHm5mg61SliwvqFwSt7deghFe/O0v5wNB3IiCob9zf69T3+xmD7xjQZODvdTQFvPMEVVaOsrK4UTzYv+ADakLv3qWB7oK0LF16t4HS5Wf0iPgEfAI3AzI+AJi5v57PmxewQ8Ah6B64CAPO6HirJAGftpNcgGIiWo53BReeqfrrvswsD15DvavCsUaYEyRSNkHQM7Sg85uS3lER5dlkaJEaO08P7B2G6/oTBBJPBp6ZZQqDD2Mwbz1DUlCwMYhh5+twgO1CdLrcRveHZh1Gd/Fva1iApLGcU+fIccMdKFOUBCQJzcq0bkBv1YiiqrEcHfEAXVgt+W9snIAfq1aAkbc1Vpq86HMWLUYx1jgexgX8YPEWEYQz5Y8WzGwhggNBh3IE35U+75f/let/Z5CnKzztJR8cmciEZB+f1tzjUH9cuuQaBaH2F0PYqDkLk8mpGJNNLNJwNrgMEUs4VKbrqhCnFPh3E4LOQWLkIiTHPXbGTFMK6HhwfDfFGG1rV6LZq9sNY9sX/PhK5RmWb8si0C4zRQo0gKFSxX/QK3v1aLSmG+X8agPcJZqTecPlw/CoNOPYkX9Uc7zXKerzyXeMaRKupmMGQzRsZdJZ53+tXBfRXmeQHzNKs2oXRpcH2KrBg91ycVxaTz7WIVpo1UF0bcX9gUUPW8LJeL3J1L4oD3Bu9Pns+7hejZ6deFn9/OQgDZ83NqC2rIhz9VnR52fNWgdp0V5YJaiX5Sv3231q1uLofnJeHNRrXglplDZTOJ3IeuAgvPeN6jyHmXdas/TMbk2Xp6/GxFNjc5dzuUeS5VSQ+eReZYozRVZSsb9puFqocnzYnHRVbsHXY2g7TfqSkx5B0qpH1Hnxlf8h+6GlfhHtcG1IBjXHzitIQM68mKnXXt+9l4BDwCHoHXDAFPWLxmUPsDeQQ8Ah6BmwqBj2u0b1ejADaFnS2lR+6iZuIGZ/a6eKbpcP4t65mLIlN+vlfbUlQarzGMVHhxY1Q8klYIAAAgAElEQVRHmbI0TyhaRC1gUL9Njb8tgoPj8RtGeBYM7vxeTZdkhjpLl0E0h0VPEGmBQsfxKWzNWDg2Y4GssGLeRhRg6IcYOKpGJAlKHdEHeIY9oIYiSN9GMlh6KUt9ZTUqUDCtqLWlbKImhUVGEKlh71xLBTOe4ujDxmNztYgTjH0ofzanBX3/PjXwAjuIITBjbntV9TFymw+/zT37TxjPB8bzQSkd5VNX41zSHxEunGO/7C4ELJ0Z90UkQ/hGHPJR9mVQxWmyjGOKbLuB1k3o4lYwRVAqiEL5ngLuyYbCKIpaLR6qzcmQMakK3L2piVqj20spKWyk3s1gTH/Nz/yYrOD+h6zYpxoiczJc3y56YlMEkfKDB3cpVVASxnpmBm4oEqOtEzYTlm4pDOMNGcHbYRhCIuXUtLjRSYtx4W2eXSMi9kYf76t0QYwIC563urEO6v45IqKPm6OlqItpERRNrWspmuaCzq/IQReWgVLzla6m7e/QtpluxFzn2dIU8g7wi0fAI3BjIcBzjTSmT6hRUBoZ87L0UAy3EoBAtPEbiE5gKfLiq7r3JSuKpi7leFOWXYVXQXxQC2JNDxHeCW/UH2v6RL5DnjVZmWdMV9t9U8+QWW1zSD/09B1nn3FtuVKRDgHHRJa8mr0n0X6p+lbWx+LpPBuuDTbX3iuC4ja3tnwsTwf3KAREo7OsqC/5Sv89Hec5NWTnb6ohVyP7mxPOjXX2/Gg8Ah4Bj4BH4KZAwBMWN8Vp8oP0CHgEPAKvLQLyvO8pyuL/1VF/Qg1DN1EG96tlrv1I6nrPnnJF7zYX75l0USyFJLKC1xg1H1FDeTuqhpaDwmRe/hj/efewHsP7Z9SszgQ1KUhPMzLoqUEKoHxZLQtAqGpNVtvBIiwgJjDu0B9jhnhYUHv/eD3KnHms0i99WS0N0iSxP9tALjAPPMRIvWQRHrY987FIDdahtLIPx2VujJd0S0YyWH0Jxs9i6Z6qc7HvRswwTrzTOA7H51xQU+Q9lWODD2OkbgDz/qZSdQXu0Z9g7ERRkKqA8TMe8HhMDaWXKIv/xDm2AfnPXYXAC+SjrnMZyFsiI7h2MV6MLK3y9J5QOpuyzF2aB2VaKvNTGUaz/WEuAsNNdXrlQRcUq8odsS8Jg8NRFK3MzybTytXf19XG/RgqnU3h61hccV2N0sA1G0ldxqIZGa5vV4TK0TgJeypgrnzm5W2KqohEWJAOqqO/9+j8zCvt1oJ2PClyqKnz0p5s1fKV9W4m0iK/CUgAS8/3khavHXIXjmqSyHgoQk/51PQuoFaF6MC9Mk0GsVI/1ZJ4j1JDrejcynu5jIbDrCaCQjRUMdmsxzJaBm3ts6w+VnUfjd6d/l7aIVeHn8ZOQsCebUTzUq/B6pj91ZeaZJGlf2ftzHOuNbs3SxoTZVRr7JHEKB+AtM9zX0TBYiw/gLLI4zxLN6OkNgjDqKENRGQrSsOVkSrh3JIOuufZtsiGp+qTc8rmFFHgW4RI/jzPD5EgtyrD3JQ+kQEvWziY3kNFf3Plvb2NlRn1p/0gKco7XqJsEnXS7lOjLgXR2Cy/r4YcjTME+sKuqFn0UufZ/+4R8Ah4BDwC3xkCnrD4zvDze3sEPAIegR2LgAzaXxZpQT0IDJAY8jFwXzR+rz4kv/6fzV22oizrSgmVTZ5ycQNjOMb1v6BGCiOUOYLI8RrD49+IBzyvMLKj2BAdwW8Y0/mb30h5xPGOqmHkolULb5vhy4gQ3mUY9rG1YqznOPz9JTUiPoiSYBsIAMZoKZwYn5EQzNNyxbMdUR6kwWJ7FvpmnPSDAQnPMfb9ohpebIwXkgIihLFaWhzWMU5LacWnfR93PfqgLyNaUHohfKw4OeMBG/6mXzA+oUYEB3NBEV13vefX3cI/18jOGuFCkfSLdUcuNqJOiKx4gnNbPbj/vqsQ4H7gmuQ6mpdH97qMpecVS7EpY3mqXDXUr2hlWZnUk2hZV/O6jBrTukDjUF+0rRLaOLn5y8LeiOu1JNwrw8hSHIct0hipT+6j3WKcftkXzvREraZHZk3REpPCaxrclBLoDTJoK32QO1TIoC3v22XZnBTZEsrrvkh0098ppkjBL2FbnvhpvR519+2Z6C6tdOwZ9rLH8RruYM/vgqiQqy0iXV7D4Vz3Q5VDlaIX98d7YkOEREdMxJyiafpJLVzXeZ8dpCIAlV6t10szapcIIKVVCzu6vXju10Veqbi9m4vjgPeJ3VPXfeD+AB4Bj8D2CKgGw9V+HEU9qCA3DzdkZWRbZM9ffiks82Hf9TdWRUhke5K6Hhc8NLrtFl4BeTp8R3N6nuI2FJUY5sOBK+QZoJRNzTCpZSqEsdpdW7592N24S4TFOW10RKTD6TBOfk/v79NFNninSJADzek9QVxrDuJGq6X39EguFUcxCv1QREVLhIfrb66KpJDYqnUiS6wu3XbD53nEXB9EfhjPmegKZEp+81EVL3Xi/e8eAY+AR8AjcM0IeMLimqHyG3oEPAIegV2JwDc0awz3GLzx2H+rWsPVD/RcPFFz+Wbq0qKvbNxKxdRAGcKARkFfiApCw0krZUoMhlL6wQiDcZ7tMJyi4GF4/5YaCh99yMNrtB39YHTnu8Wm24ngeOyPkQeigr8tIgHjPmQBn6yDxIAIMfIAL1gjOXgXQpSwPUYmyAr6sny/EBCmhHFsjP7sg3cZaZlIyUTfLJYOxPIMMzYWjm9GXLapzsW+W1oryAlSNzE+9icv8M+pgYMVKj86/h1yA6+2h1UM/afc2d9EkTSCxvZnXmDLHMGXc+qX3YkA1xrXAPcf99ZRSAZ5ehdhWfQGeZmqnsKmDBtYLmZkZO2m8rpM82JPmAXKDBVmjXqse0EVL4pyQhdytLrZW76w2V/fM9VYnWjV1mpJk3vOeY/wq19gdbFAiqwIxUYkSg+UJEmYKOuGalfkcyIyWlFZNjEdhYpwETnkWnGgFELRrIzXTmURzsmWdWJyok5B9JoIDUuLd8NezeMIkN1Uh6FUuq9MJAWRdyeU7+Upfd/Qm+FwGIQHZUxMu/20oHYJIRVKrRY3kqipc614DAU1FWUtK/IZhWiQDnFSJBX3qdWeuWHPsx+YR2A3IyAyoyfS4uvCAEcAZLj/We19an9xO1xEDrhhv+MgDeASFEWhEmQKdNRznwSNIiecyAmIBGRl+QbFhGCo7lT+ZtWbuFCkqQgDvapJR6q+tO/dbtD7H+14KqI96k+RGa4xM+9EXGizXKQImajYSux3T8F8eX6xl4v5q66IxBj3x7uGKAr0AOTjP1RDxuR9j4zKd5/+aTffBH7uHgGPgEfgOiDgCYvrAKrv0iPgEfAI7BQE5In/mKIsMMj/V2oY5/H2f9itf3Hezb4vdMl+kRbZlEuCmhuuRy6eWpJ2RKoiFDa2x/iPAd1IB5QbwsUtooDtMKYTDQBJAWHANg+rWSom9sdgA9lg0QuWOskMORwHYyxGHrZHqeKYfCfNFOQDSh+ECcQA61nH8egL0mSUrkWNaAmOM842PBoPxIFFexAxgnJGOibqVlwsdv1CJIiRFlo16t9IEv7mt1HKHP4YL/bdIjzuHI+T4+PtRhoo+mDMLNSgYEwXo1hka3YL//SH3fH/hTB95oHySBoqFsgMvoMv8/63nNPKsf3XXYSAjMd4uXP9cS1hCJUDeHlABgsZykMRccFtKrWdyXaS6WJP8jxvplmhaAAlgEpcvxaoVGjpGiIwLsjYUu8OhlGelUWtEcetRlLMTTe5liHn7N7ZRehe21RFOIQyQk/1BtktYaDc42Uwmxf5hPDOVX15XbjKizaf1TlQvYOyJ5JoTXakgNoWesR0a/VkQnbuvcJ7bXa6mf36J54c/vyH79tNhMC1Af06bSWirlAap0w1Kjo6TxtFXrZFUvT09qh1+ulELjZC91wUy406SaJUrBOnt5WmWapoC9WvGEUzKUdM0NDbolok93WakT+sR8AjcI0IIO/hRIKciTz3qBq1wt6pRn010p6abHaxy4tRDa7ER2DAY0ILb18tQ5ENrq8nyeiviyLmRZ5h9L9F/247NOpPjCIzRID01pZEiJCJEJHxYoSFyA8iOS5GXGy/EEWMzPm/qT03Hj874JBk0cIj2VWkjY+sfDEk/W8eAY+AR8Aj8LIR8ITFy4bM7+AR8Ah4BHYXAjJwf0qkBfUrMHJiEL/ddR7fdMPFvpu4t4YnthucveDi2f0uj1sqwj2huhYYLvEwNQ8syAOUOfogmgJSgKgFPqnNQA5gq4OBIgYJgOHe0lEZUVGt/2Df+cSAT/8shKZbPQnIFggUlEU7vtWvQLkyg5D1ZcQE/RiBwZgtmgPiAGWU8RBtAoHD7/TF9hhrOQ7vV9uHvizCwoiXqsesKXkWaUHtDepMsJ6i2qTYsqLZjBeShJQDLZetDl3nWM09/y8hYyAsPqj2xxxw9PvFeTNmokK+xLkc/+Y/di8ClpaM65jr9zBFP2UKIWIiHYqk0F03IQ9wVeMupmQoj2Tv6MuiMpCpoz9IC1JLUJS7q+LPg4lmMphqJSt56fLBMHf1WuS9LLe/tkpFrcQigaYUZiFP2RGpmojAyIfDYCrLioYiXIisGKUHCpNQz1NXT1VDRNtNJEoJpc9MxEYuL/1EtSyGh/ZN5TKQlxjKd+8lfcPNXOESpWInwskkCVpRFMzrHmvVYjdMVWibovZpmq8pNZTy0hNHI9oqCEVYhIHoDAqud7WPvRd49vOu9ItHwCNw4yPAfYvMiWOICl+PZMz/rPZutY+NPz+iT9KQsnxbbd+4cPaVs4PMGK19ZVzAiKBQaB7kRDYgOPLiISBJLMpiy0GV73UkryLr/2s1ioojc/IMYm/+5l1jTj3Iu+U26bKunI9f4xHwCHgEPAIegZeBgCcsXgZYflOPgEfAI7BbEZCh+1+JtICAgESgkPMht/bphmvdN+3q+wNV6ktc0VbseU2pYjCuSxmKEqubYMZ2iySwtEakUcKoDimBwd0M/JAcKHkoRxAIGOnYziIcjFyw/O1GFBgRQQorojNY2IZ9UaqIMGChH4vQsFNqfZvHWPV38142Q6x5kDMv0i0Z+WBpoDAuVomVajSF1eKozoVtmSM1JiA/UAwZP7Ux3qYGXhwLnFbVIDMOu1y5BNa/FLmFXzrj0k0UZEt59YC+o2Di6YdHHFEsz+oc/oZN1n/uXgTGURYQfJB6GFS43qZl17i9DNxmVKhQfUjd7TJQ9EQnEjtBHgnl3j/XH2ZNFYh29STelL1jQUb35TR16zKeb4rYyHr94fDWQ7O5Twd19evr7tvmAxmqlVtL9UBkpR4OcwWrlC15vPKMUkHVYtLl+kEGbXG+PXnmQ2LUldEjjWE64rCps1EfaKcsTZNBGjYnmzWeszd8aqhddsepFEnAe2xF5/uMoibuUEqvmiri9hR1UVebFTcRN2rxShwFfTk86/QGq/qedtNyqHsvSxIRhXqzjkyHPiXULrt8/HRvcgSQ75D1aOYo81V9Rzb8IzWIAIpWm9PMXxvPF4cTSy/66kIwIj6MpBjJ8rz/kV9/bTwOopJNFmVcyMt/okZENAsyA+8Zmk9R9+qeHd+bR8Aj4BHwCGyDgCcs/KXhEfAIeAQ8AteKAMrLv1AjJdKyW/7EMZccSN3+vzLhkj0iFqZS131WSddvVax5c9NF86RpQtm5XQ1FzepTYJQ3IgFjPsZ2FCfqUFjKJvMCx+hDFAYKEoZVIyX428gFxm/RCaZQmXEfYz/GfytijfmnGu1gkRHWH8ewHL4oaGxrRQhNSePdSQQIyihj41jMz1zgjKBgvZEb1fGaMmukCH9bYVUwwOudNFD8Dh4cj09+s8Lbp1zv6YE79x9EHH2WSA+UTQgOSytFuioUZbAH738DSH7xCIwR4Jrj+uC+gdhS9vxyUdzEhlIRtVVlQXbyoiujap5EUUeGjtuUl18UhiiNohxkWT6UofxMWhYrchVfd4HqWpRB79iJ5ezH36X73y9XReCeo3vL0+c3BkoHpaQfpTJ+FINcCTuyfEQwyqM1aAyyUcHmPEniNFfghYiLjgzefTEbgWpe9PsDtzrZSlTtvFbMTjWaIo94xhhB6pG/MRDIRS6p/ksx0Hle0dk5IY5pThFLIjJ00wXBfhEUSSCySoRGS7VIAv09yU9R5M4pBZuqyiiNlApZaDr+froxzqkfhUfgRRHYJsqAd2xf9S1435ocaGlTkR+JAv5343cxZIbJwj80/u1z+sSh5/1qpGb6wPiT9R8a94nch6MOCylW36Jmcuhv6Tsy5bvG+5mszDrqmhGZy3fkS5PLT+g7ji6jiD61rREU/pk0Btt/eAQ8Ah4Bj8D1RcArONcXX9+7R8Aj4BHYUQgoygKl5++rEWXRdVMPvNEd+YUJt+cDynrfrqtaoFKZhHVX3xe6oCZCYx6yAIOakRQY9lHSUJBI/cRvVqwPBQvlCAM9ihMh6WaMM8ONKXzguvUdhhJFlAILKZOOqqH8WToq6696TizigXUcE0LA0kRZ2DvjQnljPcQBx7E6FBYFwnEu+sK+kEqK7xZJUa25YXNgnaVxoV9LH4DxErz45HdIH/qnZgVExDHXX7jLPfXfy9T8+5Z6iyLdhOpDXoAvaaXw2mbc/7uiK/Du84tH4DIEVM+C6wdPStotIixmZTh1URS9UQTGm+UlXg/KMpXR/O5aEveUrmZD3uGqwuA26rXkGW1zKk2Lx5M4eE4G2fYv/vhbRgW3/bI9An/w9VMTne7wDbqx35YV5buVq2NPf5jPK72WQtXchNICJeTrqKmutvDWP3dK/5dxEjVUr/u8vp6aaNaenJluPjXRiNdVtPmEDN54zF41FZeiXfzpeB0QUJou3gfzui9uFymxT6f0ARFVB0RgNHW+9ujNEOleUiqoYE7EYFecRSFSMFQk05Nyhn5K6b8W4jha0G+k8+vqPPo6Ja/DefSH9Ai8WgiItKh2ZZHBJu8iGyNjIjMTZUE6T6IgIA/2qd2r9hU1nFB4tiDfIRciK/KMoB/rk32J4GD919RwiIHQoH4GNd2I0uWdgbMCjd+RVY3M4HNEVKiNFp/yyZDwnx4Bj4BHwCPwWiLgIyxeS7T9sTwCHgGPwE2OAIZvkRa/oWl8WG3atZ844NKVutv4ZuJad8Sq5qec66oU2D/Zcc3bjrgMO3z0rItrh/VllIedFWpEA/CJEQaFC8UMJYkdMNTTUJgwgJpChzJnBn4jMKpRDXzHOkcaJBQ1UwAhKqymhNXCsDNhpAGf1iy1E9uwPd5wRGhAHKAwQtqwrSmLKI5VT1iL2rAICyMoLBWV9W9zQVlEKbVoEuZOQWT6t1QveME9pjRQB1z38UnX/nYhsoJtwNVIGRRU+mQ9Simfn/BkhZ1q/7kNAtxz3GcD+XMfUGqoiazMF6PQPSNz6l2FimwrIdSGDKtd2c/PUh00LIN1ERXLwyxfyrKsPRyGw0Ga+bRE13CJJUmY1evxprBeVRqt4XCQKzNQuRGUsRO+0yKMptO0rPUHWYMC3XrQzCpfUL+RxPojLJPEdRV9sViLwr4eKH0IJBnAOXLgU3Fdwwl47TbhWcx77azOKynUAmrfFoVIQBdspkWxV3UugiQMNhVNEVADpohdXyTFaUUwrTndbzq/3JujcysC5IpoC09GvXYn0x/JI/CdIrDF6G+OL/beHIrQQNbE6QbnFHPI4eGOgw8yIFEQ1HtDFkZ+RsblOWORECbD4rSCQxDrkS/Z9uHx9qzjfT/qX2PyROh3emL9/h4Bj4BHwCNw3RDwhMV1g9Z37BHwCHgEdiYCMoD/sUgLSIYfcGV62q19ccXNfl/D9Z6/zdX2JS5R8EW2LLPa8aFr3qMUMoMZFxzYo0LcVgib0Pin1DCwo0xh8IfIIDx9QQ1vMtZTiwGF7JJype9GBlRTOVmRa4uQwMhzhxoKmxElbG/RE1VPsupJQnG0SBDzFEepQ4HkGIwNxZHtIBUgMVhQIq1guEWEoARart9qWquthXEtKoQoEIgVxs6xUDwtPRTbPOmyzZrrP9tyK58u3TP/wAgNcCT1FrUtKKhNKimUVX7/DOeqOkH/3SNQRYB6Fvq7UKTFyKNSqYeG8vSepSBnnge5aifoz6CQpbWl31Ro253TukKO4GsysK4XeX5ORMaiyIqe+vJpIq7h8spV60MEQzoYZh0RFudktN4vD/w4jMNzQRnx/JkMo3JDv6cqwN2IoziXaSkdZtS5yNPJRtJRBEyQlUWqJ0xfGaHYx2rfXMMI/CavIQLcT6pTEVGkfq/upeepQaLEaqEiKGIRfjXVwh0GYqsUeSFeozgXRfEgjBSp6MpNMkWN3wWv4ZD9oTwCHoHXA4ExobFVRmQoyIS2IFsiH2+7iPjgd2TCSySn+i613kgK/65+PU6wP6ZHwCPgEfAIvGwEfEqolw2Z38Ej4BHwCHgEQECkxXv18dNq97t7//Xdrn5k1kWqY9F7tnDNOxoulKGtcU9X0Rapm7ivcKFs8lGCsmWRA3iTYWxHuYLMIDT9NjWM9RjgWCxllBEJkAeQG4TNQwhABlgYPN/5jX4hHGiQFhbFwXaQAJAg1l811VQ1AsLqRRihsqB9SLPEQmi9HYd6HvQBgcE6C6W3XMBsb+9aI0ost7DV7GA8KKSQFTZ3yBv6I1LkUaXbWnSD4290Z//jvDvxSxATf1kNYoL9wI55gh9zfkztt0VWfHE8Xv/hEXhJBMbpobj+cGZpypt/Xulo9ujiTUVUTFABWFfyKGpI9nLqKnRV6EJRAgWpJbIx+fGSx9ntG3zsoeOh0muJACqOCNL7hln5PZu9wWQUhh152otoLZTTPEzzrJhOaiHnYUN1Q7qFcu2pnsj5Rj16pl6vPzw9mTyt0Iw1EUadcUqoy1J4GM7eC//1ueLGERE82yG2KVo/qWilgyIsbhFxcVgvg8MqYq8yMEVXURVNpfrivjrD+dY2Z7TNmu4/iGfeBQOfEur1OY/+qB4Bj4BHwCPgEfAIeAQ8Aq8PAp6weH1w90f1CHgEPAI7AgGRFn9JE4Fk+Cl3z6/eKqKi5YKk7qJ66dLl3NUPxy5oZjJ0Fi4+uOEaByEKCGcnBdKdaufUSA9FmDoGfYztEAxvG/9N1AFGG34j8oLtMeCwL1ENEAMQFBj3eaexLesx3GPMZz0LxjzWQwpYSiYIDtYdVyMiw4poQ1LQF/2yMDZy/tInxieIAouaYDwQMOQcpq4Hxl7LJWyh/lbbgr7Me84KaROxwXcIB+Zo/TF2xoUx+Ly78CexO///zLuz/560VODAGBgvWELiGNHxu/p+wkdWjM+c/3hFCIi8GBWnV079uiIA6iIsEhlcExlQZUcNhvIOHypSIE2znPvJkxUvE+Xf++rJZGOzPxcn8e0iLt4i0udOERYqcB7OyM1+XhEtU/1+WlPIC/UOuLf7ql/RqdWTE0rP9djUROPY1GT9tNatRVHI84nnha9h8TLPw/XcfExYcB/xfB9FAYrkg+y+R/cQhPuU7qm+CnGf0E01oexQkyp4f0bn20ho3kO8g0aEoE/3dT3Plu/bI+AR8Ah4BDwCHgGPgEfgRkPAvDxvtHH58XgEPAIeAY/AzYEAxa0x7n/eHfu7D7t08Ywrej2Xb66JrBBN0W+4oAhd/3TksqWmG25YwW0iEjDMPKRmdSUgG6gP8V1qFKB+RM2MNhAFGEcx3piRnv05NqQEffAdAsIiKPi0OhjsYxENGP05Lsagb6pBNLCt1dTgWBArRnYwZgodEg3C8milLyM3+M1Ss1jUBn3SbLH8whzHUkFRc4PvjI2xkhoK0oJGruKz7sxvbLrH/1ZbZAVzYywQRJAUp8efbAcun1fj2JwTv3gEXjECipbgfkqHad5TFMWmDKukl1iSwXWZ76qvsCmygvvHkxWvAOUff9etabuXrrQ7g+d0w369oQLm6ma5N0hP9wfpSTFBy4qo2BDWZ1v1+NRks9atJ/FqLQ6eaNRrIimCDaWCGoqs4H7//9k7Czi5quuPvze+Hnd3JSHBKVCsOAUKFCtaoNAibSnQYqW4O0WKuxSXBoeEQJAIBOIQt91sstnd2dH3/r/fMC//YbIysy6/+fR0dmfuu+++773vbTi/e87hc8cRSesxGh3SFASSAkPiPko+l1GDJBE1MQ8RFEwNtdzjcS1Huqi1EKgqOKeYTrbn3wfn7xaFcaVvaYoJUp8iIAIiIAIiIAIiIAKtmoBqWLTq6dHgREAERKB1E8BO/k2IsngGozwHFjS+P326MfLOfeFiCRpFyCbj7oxC3OGA4etRYVhRZOteBYd71VDD03UVUkbR2f9L2OqkQ4f1GFhYkM53Rl30hH0DY60L7iKmc39Asg2/oyOIzh0n6oCwKBDQweOIBc6uY7blZyxmyHdGLzCaYyRsRPL8TkqoVAcRBYL1MEZ68GfWxHBqRnRJjol/SymIOC9HsEjUB4BRqOBnjjBDZxQ/Y1SFk/rJKZbN3ynMlBpWLGCsfXi4sfDCYiNeNg+fMcqDYgUZUayguEGHFo2CB/t4hnOSMhb9KAL1JcD7gGvWKcrJNcx166Q2M1S3or5oDaNLUY6FCJayaMxi4Mqc/AJvv2Ao0jMUsUJ+v3tdnmkOQHRLoKggUBIOxxBtYZf7PJ7VPr9rfY7PtwlSBZ+fvOedejlybNd/OprkSIoWiLTgvDi1jThnnC+K7fw7Esbkcw6dCBn+bWCKPz7D2ZZ/t6rLad8k41WnIiACIiACIiACIiACItBaCCglVGuZCY1DBERABNowAYgWdOb/A+Y1PJ1GG31PixmdduuJuhXDUSw6ZuSPyTcqF6wwzJjbCAxzGS5/zPD08Rq+fCcqYV3i2P8vHssIAwoUdOQw3RLTLjHCgM55tqPjlDUbGB3hpHtyHKp08jjpkhyqjohA5xF3i1OEoGOIAgQFB0ZTUABIfbEt+6aA4uT25/k5Hh7LiBCOkUDHD6YAACAASURBVMc7BbidyMXUv690OG0pfphyAooTHCcFCif9FAWVYiOyfqhROqXE+O7EOfid6arIgWKNE7HB+hQUSYbBFsF4zddCrGBfeomACLQBAg9Nme/Oz/V583P9RW6X0be8Mtw3FLPyAl53FaIrBmDnfTd8vwEphELhULTc63XPLyoMbAqwYrMHtS1+em7w+RJVjYPWOeHJ1FB8/ju1lhyBm39HnFpJ/DvIZzuf4/zb4qQ05NzaSgfVOudWoxIBERABERABERABEWg6AhIsmo6tehYBERCBDkcAwsV+uOhfwoqMPqeMNTrvM8Tw9cw1PF1cRnjFEqSI6mp48tyGt1vA8HaGuNElYrg6rTXcHjr86aShA45OfDrz+Rn/TtHBQ2GBDh5+x2gLJ0UUBQtGWDgRF2xPx09qlANFBAoNjpDBn53dq4yScGphOFESqbvInVoWTs0IntfZEUsxw0kb5URScM4pdKT+fU3d+ezsiKaDio4p1vLgZ0yB5TbiFd+gVsVko/i1XkbJm7wuJ+qD30+G8TiKEhRcyIhiykcQKqbwxHqJgAg0nACczOyEz52+yXt5JZzGTk2ahp8gpQcW4Q74PW6k2coLR+J4ntm5fp8nDMGiF2tZIBVUCSIuTI/LDAcC3rV5OT4bqYP4fOFzgM+QRLFtObUbdVqapDOsKyctIPvn3xvOI8VoRxDnXCZEClgiOlDz2iRToU5FQAREQAREQAREQARaOQEJFq18gjQ8ERABEWhrBCBaHIcxj4P1MAZetKMRGFhoBAZsMAL9uxtWON+o+rHEyB2aY1hxj+HrXmG4vZ0Nd7cqwx2go4ZiBJ1wdMZRYGD0ACMfBqU4dViwlCmanPRPX+Hn3ZLHOcKCIyTw7xydQE7hU/bNKAZGK1C4YP2H0TA6jygGOH8XeQzTeHA8TuQFnUiOI4ntndQ4jsCRGsXhfOZMH6+Nu2md1FA8loIEhQg6plYYwfl5xoa3xxhLrnwNKaB2xmcUJFjrg2IM62ZQZJmUfOe4KVrMhVjxtHMSvYuACDScQFKwYPTU3rBtYR8n7lFGP/0kEm6VpgeO5QadmIW4SzZW+m3D9LlN04N0UN4cv8cP8SKSk+N1F+UFmDsqCHEjEVGRtIgc2g3C3uwHJ0ULR9R2/makC9wSKpp9ZnRCERABERABERABERCB1kRANSxa02xoLCIgAiLQPgg8i8s4FDbaWHaDx+hz6jjDXcTogXVGeE0I/rh8w9fFZ8SCcMDDb+MucBuuKtvw9vYbnlz461wUDigYMHXTTjD+reJnTAtFhyGjMOjMZw0IChdDk9goIlDooNBA5z5Fg9Qipk7qJ4oprAHBHOLc3cr+nILbdCTxXDyWYgUFEMc5yXf24eyAddJTpeeOT00L5URe8ByOIML2HN+nsKBhW2VGyas9jWU3uY2yz9iO9TsouDB6hONiPnMnmoNjIoMlMNa1eC157XoTARFoXAIUGCkKroHx2bJj8t5jKjregxQwGq2+AAtxX/3kl/EBvYvCECncsbhl+v1eoyjfb8dR7bysImT37l7g1ORJPHMkVjTuhDdlb0kRjKdIXTPO3470dyOlfWJYDRXEmvLa1LcIiIAIiIAIiIAIiIAINDYBRVg0NlH1JwIiIAIiYCDKgmmWuDv5V7Bcw3TnGoP+3tXosm8/w47FDFegh1ExP2zkj3IbVpXfiAcZbRBCNEaO4R/iRY2L9Yi8oFhAZz2FCTr4+TtFAkZH0OnjCBQULwYlP+POY7alY58ppJy84U5bvlNQYDFvRk7MgG0HoxDB81AgYNon7qLmz474wBwxTB/l1MtwCmk7URf4KtHWSRfFYxkBwvFSROHPHJMTRTLdCK+cbZR/3cv47iSXEStjJAVFCtakoIOUURW8dkaYOLU9KM6wLzpS34G9j+gK/qyXCIhAIxJIcRYzbIJpofjaHkaxglFavFf5jOBzazWssqHiQbqDOu1yakoxt6WZHNqNuADUlQiIgAiIgAiIgAiIgAiIQIsSkGDRovh1chEQARFovwQgWlAc2AW2A4xiQzej1/GDjaI9RhlWmccwA6aRM3i1EV7bz/D1ChpVC6qM/HFRFO3OQ9QFalsEqvA9nfcUP36EjYdRWKAz3ylQ6ogLFCcoJlA04HcUDOhQZJQCdyU7qTf4OV9Oqij+TMFjZmJ8P4kWFD0oFlDQoEhAUYJpqDgOCgZOrYvUPp1ds85nHPcsGK+fAgojOShYUMD42Jh94EKkf6LTk85Qjm8kjOLDYNgHMIo9fPEaGA3C4+gs5fm/gE2HWMHP9BIBEWhkAtWIB7yve8PGwBjp9QOMz7QhyXuUwgXveUZdJGpKpA5JYkIjT5C6EwEREAEREAEREAEREAERaNcEJFi06+nVxYmACIhAyxOAcNEdo/gzjEID3P29exm9T+1iFO00wnDllhrR4k6Gt2vUiG4sN+xonhEt9RkFk2xEWaw1qn6wjPyxm43AkKjh8hUhXdRz6OEEGJ39NIoI3PHspGfiGfg5HYYUHCgU0LHoOBD5d4+WmpaDxzPFy1IYHY/DYU6BbwokjH6gE9IRL9inUxDcAUzRgemcKJawRgZTyVAsYSRHDPU6Kg27KscILu5jrHsCpbZvZU58ppihw5NCBJ2dFEXIaA5sIowpn3gtFFT4Wge7DUIFx6qXCIhAMxJIihh8dvB5QNGSAiNrylBkpBBKQYNC5yewxTAKlVteEi2acbJ0KhEQAREQAREQAREQAREQgTZNQIJFm54+DV4EREAE2gYBiBZ0xLMwNqMtWDvCNgrGDja6HxkwfH26GqYZQWRFd4gW64zcEUwRlQMxA1EYaFc2NWgU7hQ2AkNRoDtQafj7UBigqMC/YYyIYOQCBQQ6CClM8GcKEhQd2NYRMFILnTKKgiIHv6NgwT7WwhihwX7okOwDcwQLnos/sx2PcQQS9sNjKGLwnPfClsFYNHsy7FsjvHqgEVyw3ih9H4JHZICx+rFlRmQ9j6OTk+IGhRAKF9y1TWeoU5+DIgbPy3ExqmIqxAqKFnqJgAg0M4Fqoi5431OsoPDI5xCNz4bPYHx+MN0cnwUUM1WDoJnnS6cTAREQAREQAREQAREQARFouwQkWLTdudPIRUAERKBNEYBowXzwLCj9WxjrUHQ1/H3nGHnj94cIYRq5QwsNE5pA7rBucOhDXIhXoZ6Fz7DDUURgxAxPZ8uIrFuLY/yGr29npIyyUeeCggSjLJy0T3xnyhYKAnxnxAMdi6m1JpxC2PwbSOGB70y15NSl4DErYYzQoPjBPvkZhQxeA493IjU4B/yd372ZuCYeG49ONqxNuUbVj9hxHSswgj9WGps+jRlrn7GN+CYW36b4QaGCQgdFiFSh5EP8TmGH0R4UNBhVsgJiBeto6CUCItBCBGqoM8FnA4VGpovaF8Yoi9EwRmX9F8Z0dhQf+azZEtmliIsWmkSdVgREQAREQAREQAREQAREoNUTkGDR6qdIAxQBERCB9kUAwgWFhP1gB8OqDC9qWbvzhxqunGLDQgSCv08Xo+dv84zYJtsI9Hcj8sJjeArixsZpFUbhJBeKdCMiwvIZnl7rjcJxcAwGvKiHscxwe+g45A5npmrhDmc6B5mmxSmeTZHAeVHQ4O+OkEFnItvR+BnfneK6/JniAR2RjBRxCmdT0OAOavZTAn1lsVG1ZLLhzu2ENFfrDcvqZ4SXFyPNVcDY/JXL2PC/NYi04Bj54vjo0GS6KgoRS2CMPKFzk234+RuwKRAqeF69REAEWjEBiBl8DoyADYNRvGCRbj4f+KxZBPsSNheWiLjgS6JFK55QDU0EREAEREAEREAEREAERKDFCEiwaDH0OrEIiIAIdFwCyYLcR4CAk0qF6ZsY1fALGB1/dPIxJVMUAgbc+736GJ5uG4zCySGkiyoyCibGIGi4jJyhmxGhMQq1LapQ8yLPcBUVG54AC1UzEoKRF0zhxL91jGrgOdi3E0nBCaA4wegICgROwWwneiI1eoNtKCSwPYUGR0SwjPCaqUZo6c5GbHOpYVXivPZ6w9d7lBGvqDBCK3wQWEqN5XdFjaqFUGYS6Z0ogLCv1cl39jcN1g/GehYUR2gvqbA2p0gvEWg7BCBc8P5m3Z4jYbznmeKN7xRPX4a9D6Fii2jRdq5MIxUBERABERABERABERABERCB5iEgwaJ5OOssIiACIiACNRCAeMEC0wNh3JHMwtPbwBjdMAi2Auakd2L0AQWHkTCmWOHPdAYWGoU75Bm9ju0HASNo+AeWGTmDSg1XXk/D5WYUBAtgM6KBggDFCqZvoVPRESjYD6Mm6ESkyOH8zKgLigkUF5w2P6WPiscgLNheI7QIUSHhPkZ0A+pulKO9z234EEASK3OjBodpFL8aMUqnzDIq5zGKgvnuKXSwP6bGWpocCwtzU2ThDuxlEClm410vERCBNkoAooVT84bRZEx/x9Ryx8IojF4NwYLPMr1EQAREQAREQAREQAREQAREQASqISDBQstCBERABESgVRCAcMHaFnTmnwF7HbZ38vdVeKfTj84+ChmMUuCOZdZ/4O/czbwcdS7GG132DRlFOxQagYEhWMTwD0Ax7y4bIVywDY9h/xRA+Dv/BtKRSHPSRpEFRQqKFnynaMHzMsJiE9I8FRpWsMSo+qHU8HYainoUbogVESMezkHaqnIjutlvRFaVGBumlBu25TGKX14MYYOpniiSsE4Ga1L0TY7hfbwfAnuAv0OoYK0KvURABNoggaRIwWcK09LxHt8IY5QWny+TYENhjCB7B/YURAs+X/QSAREQAREQAREQAREQAREQARFIIyDBQktCBERABESg1RCAaMFIhr1g42BMCeUUvabYQGc/oxTo/Gc0BEUFOgQZncF282BMBWUa+eMto9+53Q076DHyJyA+orvLcOeshbkMXy86FPnqAaMYwWMYgcHoB6aOYpQF/z6y/3IjUvojojVGGHZZpRFaGzTszRAnunqNyoVVhjuQg9obHiNeifRPK/NRCNwyYiXrjKU3rTEia+iQdGphcEc1RRdGhPAzCiBMCcWc9h9ArJDzMjkpehOB1kygmsLbTtFtPkd4bzNCzEn/xu+Ylo7PKL4oyn4H+ycEC0ZV6SUCIiACIiACIiACIiACIiACIpBGQIKFloQIiIAIiECrIwDhgg6/QTCKC51hdAYy4oIpnihO8O/XD7BtYYxcYOooRlugCPeWotn43NPV6LLXYqPrr/qjpkSB4e/nNgL9IkZw8UKjx+FIGVXQEzUokEaq1wjDqtgEYQIChhuORBciJVaH8NbJiG00UZ8ihoLgm/G7xwjOyzcCw1D8u9I2XB6kmPKZqKuxzqj4tsLY/KnXKHmDURmzYEOSY6E4QaclIyqYGsrZeb0UQgUFDL1EQARaOYEUocJJ98RnEiMndoVRpGCxbaZ14/0+H/YtjOnuvk8+qxhhsXvyOXUbBAs+J7a80vrfigbas36OXiIgAiIgAiIgAiIgAiIgAiLQ7glIsGj3U6wLFAEREIG2TwACBmtPjIHtBBsFo/OPAkVPGAt3U7xgLYhfwYIw7nTmO6MkGElRapjuoYiuCEBk2Gi4OyGSw1VuuHMhJFidIVS4jK57dzEqFpQb/s5Bo/sxI4zwShtREhGj/FvT8HVzGYH+SPm00Wvk9IsakU0xHJtj+Ht4jE1Tg8bqh581IiUcF0UKFsxeB2MkyBIYnZefw76HQMHx6CUCItDKCaRFUvDfy4y+Yiq5HWEUKcYm3/msYbQEU9cxlR3bfQ2jOMmoMEZXUXQ9GEaR4wMYoyxiECG2UEiej+dxauvwOz73+Ep9blQrXKT21crRangiIAIiIAIiIAIiIAIiIAIiUCsBCRZaICIgAiIgAm2GAIQLRlcwvQqNDkOKGHTq0aHHaAXueGZaKRblZh55pndiBAaLeTvt+LePKaAY9cDUUuyzGEZHIMWNkNF5z0IU8C408sZ7DDNuG6EVMdSksAw7imM8ASOyttzY+MECI1rSDe2ZzmkmjFEhzjm4q5pOyWU0CBXcda2XCIhAKyeQFulAMYLG6InxsD1hpyU/c+rpMHUdnz03wlCzJiFUTodRtOTzha/tYNvDWIT7GdhSmJ0mWDiRGzwfn0U81qmt40RjOGIGj1XERStfSxqeCIiACIiACIiACIiACIhA/QhIsKgfNx0lAiIgAiLQCghAwKBzcB/Y/jDWiFgPY954ihB0MrJOBOte0LlI0cJxAPJ3Fu2m0YnINE38m8g23C3NXdIwF/qHUPGT85Cf83zcMU0nJZ2TFCJYxJtCB3dT/w/2HgQK9q+XCIhAGyGQIlRQzOwHYzon3vN8rlySfKcY6rxW4gcKnbzXP4I9nvy9AmLClogI9MtnyXkw1tvhs+YRGAVVI02woNjJtnw5wgSfVxwPn1MUKNiG7xQw+EyScJEyIfpRBERABERABERABERABESgfRCQYNE+5lFXIQIiIAIdmgCEC0ZScAf02UlnH39nBAWFC6aN4jvTslBcYMQFnX0UNugIpFPSyc3CNC4ULeg4ZFs6DFmYm20palCg4M5pvrOeBtNO0YF4L+xbCBX8XS8REIE2RACignOf857eAXYCbD/YRzCmehuRcjkUKN6EvQH7Kvk8qKqlJgVT1j0PY9TVDNhbaLuldg3O7fxbnGIEn0OBSDRuGrYN0cPMdblMD8yKWZYXPzCaKx637FL84oiifP5IuGhD601DFQEREAEREAEREAEREAERqJ1A6k4xsRIBERABERCBtkqAIgR3Ld8Co7hAkWIcjNEVrG1BpyMFC0ZgMDqCKZz4GdNG8XPmnOeLaVu4O5qpnFh7gimmGKXBCAoKFvysP4xRFnNhFC8obGyCcQx6iUCLEbj6yS+dmgfm8IFd7UXLNtiXnrD9ltRBjnOc6YT4c0dOK5RkQaGC9zYFid1gFDZHww6B8d/ITlTWh8nnwrt4pzG6ioJoXTVpOB/bwiigMlKCkRHVpYdLRFLEYlaXuGUVBkNROxqNV7pcrhyP1+X2uMwiE4V2oi5rncdjxvBRvCoUNbxet9u27Cjeg7ieRMRFTYtPNS5a7LbUiUVABERABERABERABERABLIkIMEiS2BqLgIiIAIi0PoIILKBjjqmZKIZiLigaPE2jGJEqnjBFC507DGdC4+h0MA0LayJwdeK5GcUP1gcdwGMzkQW200VKSheeHBeihV6iUCTE4AYUdM5+G85muX3eRL/rivK9xvhSMzbuTDHevWL5aGi/IABJ7i5YVPQ6top12L6o44qVuDandRLg4BqZxjfmVJuMozCBIXHEhifDy/DKEzyecHPGI1VqzBA/inppfgcosDJPplOjsduJVhAfPDYtuGpCkeNaNwqKq8IF7lMw+0yXUY4FtuQ6/f28bhduW6POw+RFX6PO15smhgLzGWaQURk2D6IFlwDyXE3+XrUCURABERABERABERABERABESgqQhIsGgqsupXBERABESgWQjYtu0UunZ2l9NpRyGBv5eapsn0K/M4GAgZFB+GQ2hgpMQH+J1iRplTFDtZ1LsIvzNygu0ZhbEIvzvFc1OvSWJFs8ywTkICiJSoFgSEDKYv4w7+IJzcfsM08y3b9sGJDYe36SkrD5WGwvEIdu5HyyvDkWWrN9lriss7XMHmpFDBf/fmwU6BHUpmvP9hFBP4M0XJZ5Nt1uKdYgUFhp8VyM5iRbLfCTA+R5hu7sPU+hZOPzHLzrUsq3NFMNoLmaD6W5bdvSIc7R1HHqhILB4O+qJ9c3O8cQRUhF1usxziRGeIGT/YhrUmP8cfxTPQj7mtghjFLjt05EwWc6OmIiACIiACIiACIiACIiACrZSABItWOjEalgiIgAiIwM8JwClXHRKnOC13MlOMoDlCQiJdC4+DaJH4OSk8UKxIvBxhIuV3Oie37IBOChuaChFoVQSSqZ8oyNFYd6Gn2+WKu90uphwqrArF8jweVxEc3zlWpf3j5orwxljc2lQRjDj1EniPtGvRIiXKgdfMVE+MdGB9CqZoOgzWDXY/jELFFBjZLYQx3RMLZPOZUVfKp9rWBYWkI2G9YYzYeg1GcWTLi2mplq7a6CtACEUoGitAGqiehml3wVwVVlVFelkWRSjTi/lEBJgdC/h9UVfciBm21Tk3J5DncXlQ48JYb9nmZr/bw/MxYizC9FAdNYKmtgnRdyIgAiIgAiIgAiIgAiIgAm2DgASLtjFPGqUIiIAIiED1BBynK4vR8mc67ShaJArR0nnHwyBaWBAt2EYvEWgvBBJpoGBRpAcqxBr3IWXQEq/bdMPR3Rm/e6NW3IsCzZ1RpXkjUkQ5UUJ04HsgekRT61u0FygpQgUviUImOQ2ADYPtDRsLy4ExfRxTNc2BTYWxiDWFnJ+JFE7th5Ti2I7ow/63tE1p56CkIHI4bAPMqYmzlUiEyAhrc0UIU2YGopFYP8xhXzywuuF51c3rNUsxd1WImDGRLcpnG1G31+0yrLgVsKxwfq7f0x/ihi8n4Fnhcrsq8XMEqaM4z0oN1coWdC0p3ThSrilnXTl/u352BTVFWLWyy9RwREAEREAEREAEREAERKBRCEiwaBSM6kQEREAERKCpCcCBV9sp4J+1KUjQ6UiHj+MA4g70xN86fM/3OPpp1zvLm3oe1H+rILBlXWM0EOnMqOky83weVw5SCw2KxqwhyAdVgQiLYji8XdFYnPcG8wXRIc+fE2nU4ESNtxfRIk2o4L3eFcYaFRNhO8FWwyhW0Jn/Fewl2PswCgoULqp9LiT7dZ4nfCc7p46FE+FV3aKgcMr6OCzO/TWM9XG2emGuTBTb9oRjcTfiwAYYEWu8bdh5KKbdGREzXcIxK2Ladj5SQMXCkbgdc8dtRNP0rAxFq4I+T7Awzx/Lz/WaiKipgFjRkIiQVrGw2+sgUgUH3HfOHzMnnSHXK9eLI6pvEZzay/3ZXudV1yUCIiACIiACIiACItA0BCRYNA1X9SoCIiACItAyBByno7NLlY6fLfUnJFa0zKTorA0nkOLkZGd0eHJtM9URazLQuocisS54HwMHeKcwyh9AsBiFXfcU8fg967LQKcrURywgzdouVclIi/bi6Oa/a8lkdxjTMVGgoGjAtExLYC/A3oFRpFiNqAiyyORlJyMs+FxxorlqO45j2BdG0YTtZ5B/epqmNz9eYBTm+zFmM9e2rADqU0BfsgPIYRdBqqeQy7S9kFf9EC7cfh8kKMw55tM2DbMnBmJHLcsXjSLuImpF3G6rW8wwK/C5hcLccYyXdTckzmYyuy3Thvci1wlFRIqJ/JkpwxgVxFeiiDruT0uiRctMUGs6ay0ROqk7OWq83xWh05pmU2MRAREQAREQARHIhIAEi0woqY0IiIAIiECrJ1BLBIacdq1+9jTAOhxSzk5+Ojn5M9/9MKY8y3e5zKjHZW7GDvxt8eWAuGV0Ze0W/I8OedY1mAxj7RY6QSlgOLUUElFHOLfd1pyiaREV3KnONE+7wSgSULA4ADYb9hasD4xpn16GVVVX+DqDFZgqhlbbPCUag7UyWCeDIglrjLAujlNb52fHoiC66XabPkTH9MB8uaFHVKFGRTeXx42pNKP4LsflRtov26iIxu1gLBYvgqARCPg9rhgUi1A0GqiKeCIYnMc2YzbKYbghWDjpwvTsy2Bim7NJUnjk/DB9IYuyO4JFZ/zs3NcU2Xl/8z2IY8K4P9uLqNicuNvNuSg44PnC55yxYVPQtWjZBgPCtBmNxxOfBaugXP4kYjvRX+3m2nUhIiACIiACIiACHZOABIuOOe+6ahEQAREQAREQgbZDINVZTgcVd2QzmoI/d0P6oB4x2+hi2dYwiBdD4OhmVEE5RAsKGnSEsj1fq2B0hDIFEiMuEvUsYG2q5kE1dSr64hqOgh0DY+QIBRleE8WC72GP83ohVFCwqdcri2gFOqJ3hNER/SGMqahmVnc8RaIbnpuFjE8GMj6ZyAnlKkXGulLLsHPcLJoet3uiNkVFLBr3bI6E+ni8nkqXyxVCDQtoGrblhns7FreLKoOxnpVVsWJEZMT83QqilVUROy8HJS/0alUEkmIFRQlGPHFt8t50HMwUL7on1w3XTE8YhS7ewzGKinjvsDvok4Juel5ICq2tao6bYjCOUIG+XetLK90VwbAHUVfQNF0+d9TlhWgR8vs8iMoyrapQlM+9hMDd1kTopmCnPkVABERABERABNouAQkWbXfuNHIREAEREAEREIH2TcCJpnBqKNDZyX+70ejgZDRBHwgTg+HJZGHp8XB+01cFgcLukhQsGFFBJ3p/2I+wNTAWhKYjdDGsTRWjTxMreF3jYUz91AO2CLYt7DXYAzCmfloIq8hCcGjoiqITenCSN4WU52AUiLZ6/eTAxi7pqIFwCjseCHhQn8IMRSPxGGqRVCHIIsfjcm8wPa5OKJlu+jxuBFhYnqpwzA2XZOc8vw8lLqwwHJbDUMtiMxyW4Ug0zpoZ0TzGm+jV2gg4kUAUI5imjEKik8aMIiPFRM4f720nXRnXOAWMSs5re3dCVxNpllo/JrVmDFNltbb5bfTxJMWKxHMf9zbDrnxut7uwZ5c8o6winOdyx808l2fTJsTXoVZR3Od1sx05RcCSz3alFGv0WVGHIiACIiACIiACzUFAgkVzUNY5REAEREAEREAERCA7Ak70Ax2WTkFevnPXNR1RdGAOgnWFRtHHZZr9IFDQ0enGO4+h85NOT37GHd2p0RTF+J0589lfrTu3sxty07ZOESvo+KWDd1fY72EULFhIexrsU9iLMF5js6VHSY6NPEfBmIaLP4+Bcaw17Yx3of6EiagJZIKyraqqWG9EVPRA7RGXFbPzLCgWPo/VFSJFARJ8BYJVkUQaMHwfiUVtb9xnM4ojjMIXm4OhSAmEjIoAdlr37l7A666tIHjTTpR634oAnMdcB17sjM/H/FFc7IUJCiCVYQxzz/u52J7TOQAAIABJREFUADnceC/z/uY9yyLtnG/ep/ye0VFM39auHdCOCFFTRAUYtOvrT104ybo5iTRhkUgsjzVrkAYqEI3EukfjVp7H60KUlWn4vZ7cSNyKhMLmZjwXyvj8wDPDiUbhM0LRVnomiYAIiIAIiIAItDkCEiza3JRpwCIgAiIgAiIgAh2AgONworOSTium+qAQwaK8jkOaQkQhLBciRSGcn3E4Peng5P56/Gr68TmP5TF0hLJtEYzHMcqiF4wOLRb3jbfmPPkpYgX/7ToatjeMgsCgpDGagjUqWOB6fZJRcy8Tsj8Rdkjy/M/gnQXOa3olcs4HfO7NUCw2QZTY7DbNDS6EVUQjlg9RFj6U2HbB3eiybbMKvxv4LgoAq3FgeVU4ikxSBnyXNkWMGKJr4rlIBYWf24wI1dwT1BLnSxUrcP7O0KEgQCVSuuXgJi902aYvbtseG6ncMJ+lmL0g7lvep4yO4hrh/cvnQUL8ojO/vUdaJIWLOuvGtMR8NuM5E6Ij0jwhKxxWiGV3QQq4vFAk1jUaszwFef4KPN1tRFQUhqriBsSLeEGhL1xaFo9DsOCaoWDtST7b+TdDLxEQAREQAREQARFoMwQkWLSZqdJARUAEREAEREAEOiABOikpVNBxSXGBvztOTDqhKGjws0I4OZkXn2IFHX1OrvxEUVa86PzicUxTxO+cCAs6tbh7u9q0Ra2ItxMhcgTGdAqMKa4WwBhJcQeMYgWjLHg9P9tRjHRQzXEZZDoRdjiM0R+sEcJoD6beqvZFpzOciRQcQiiavglyxA9oCM8khCc4tqFP+BF9sdZ02T2siI3d+WYEkxkz3C6oUXBexuwgduzHc/2uAGpWdM0JeIrzUXUbNSxCvxzTQ7uqm2PWMzhH1065LqTrycE8d0ayrz6IoumJ3F7bYoLcKGASQAWTmMsyQ4ZpY2KNqG0ZVbhRea8X455m2jfUpUmIF2uTp2tTadwyQKQmaQSS0RUmxAkfBInciqpwZ5fL3Q9rJGAaZh7Wibe8ItI3ZsWDEC5sP54BkahdBHGjAoJX2OvxFPt9rjUVwQif62Z7j8zRAhIBERABERABEWh/BCRYtL851RWJgAiIgAiIgAi0DwLOv9PorKcQwSgJfkYBgz/TqUlvPOtY5CKiwhEhKEwwNRSd6HRY8Rj+zJz5LOzLlEVMS8Pc+Kxjkeivmvzx3MndoiSTkRUUXfrA9oedCWO9Cl4PnblPwF6Bsdg2r3vLq5mECud8rF0xDPYxbDhsCuzb9DFVA9MKR2Ihl9+zCU7tkphp9vZ43BE4JisN21wVQponziuc251dtuFHzQoTykW+1+cKmYY7jNoX5cgptQK79itQiTdYmO+vgkmsaNFV+/8nZ50SE1l7TNOVj7rq+VCihiEEZiyczrxvPabbLIW8BqHR9mDeKxAh1SduWLkQLVbB8cx7lKnfKChy/bO+xWaY0n21kvltwmEkUoihMEV+OBzrV1UVH2CY8d5I/9a1KhL1Qpgocpmu7rjRTY87uhGLLOjzmp3yc3wb8DzYgBRSFlTNyoJ8XxjCBvti4fYOk06rCedFXYuACIiACIiACDQTAQkWzQRapxEBERABERABERCBLAjQ6exET3DHPf/N5kRJ0FnPz7h7n8IFUyD1YoQFc+Inv2NbJw0I+6Iz30kvxXQhzJNPJ7sjcrS4OJHKJq1eBYWJI2ETYEz99AlsPoyCwPew8mYsqv2zKUyOk6yZYot1B96E7QV7FEZnc10vzksEWZwqMEkbkPZlJVNB4bMeLGsRj5sbMXXIBOVyeXxweVt2mLurbctcj9/nG5bFQtzrUQhhZSgSLVtTXG6jhoUEi7qoN8P3FCuKCgKecDieh7CZAr/X1TUSi/fDXBb6/J61cET3RJF1fpfnMWy/22PmoJpFrm2a3RF74UFqrxJE2RRjcS3G+uD9yggqihZK79MM89dSp0hGVxgQJYyNZVWuaCTu2xyMQoC2ciF0dQ6F493iMdtnmfFOcdu0PB481hFVgfH68TDp5vW6w3gmePBgQGoxowKFuFGRO+5E5rXUZem8IiACIiACIiACIpAVAQkWWeFSYxEQAREQAREQARFoNgJOaicn9RMjKmh0kNN5SbGCDnwad16zSC8/53Fxbu2GiMG2NIocPJb1K/rBmLKIefTpHG9VNQ/S6lXsgPFNhnGHOXelM0JkOexd2BoYRZsWcdCnjJN8OTbOB3fFfwNjuqo6x8W6IXBsx3xeD3ZIG2viECvglISf0e7Enz0uOxaN2WVRw1phxGx/HCshirT2XstY6fNhg77HVeb1uKqQ2z5UEawKTxjZO9pS4g2uV680Aj6vy1UZi0FqMvLhRB6KyIm+McPuGQ9H+8YtowCCRMg0rU5YKQFUIVmDe9YDdcrvtiFAuowlMWypZyopfM+1xHvVSfEm1u2cwJqScjNYFfUh8sqPmhVFhmUPtQyrK57pAYhbITwLCiw73iUcsWM5Xg8Ltq9FQe6QyzS75Pi9xYbPU4XaF3F31NyAdVWCSC6lEmvna0aXJwIiIAIiIALtiYAEi/Y0m7oWERABERABERCB9kTAibKgo8mpW8Hrc+pZMKc9d/YzSoJOcxRehkIBp2fSsZlatDbVWUWnJ1NF0RKFn2GJYr7pr+ZOCZUiAjAKhHUqWA+C42VaHA6QUQuMrFjJMbeSyaYjOQhjEXDOxdOwLbUrMkhNZZdXhsOFef5SiBVeOLYNl5tphIyuEDK6oZZ6LhO8oCB30HQbEaR8iQSwaxpyVDHKHvyYG/CWAsTmyqAtsaKVLIjkMMzi0qDX7XLleDyuroim6AHhIhd3qoV5LnK77E6Yw/XRuM37NRfqItL8mBsRWYH0b3YXrO7euK19OK7ctrGn3k7cryziXmNdlNZ1+RpNfQhQcHzv27VmLGa5QxEkCOPzwGX6UPvEE4nYAayPSkRb5KD4TT7WiN+KcWHECrCm8JG1Eanhyn0+92a3y12EtVaC3+M+b9yEYFGf4egYERABERABERABEWgRAhIsWgS7TioCIiACIiACIiACtRJw0jjxPfXfa4yicFJBcUc/UgYlHJkJ0QGG7DHULEw6+WlOP/yZURYUKFKFEKYS4Wcmi0C35JykiBV0+m8HYwQIxzY3OfaZeGckCSNFtow1A0Gg0S8rZaxM1cOiyIysKIK9CFvkjC+TsSWjLOzNleHy/Dx/zGO4InBwmx7TLvV53CysjXT1RiAv4CtHapeNFcFQBRyRSxA7s87ldQVzAr7NBXm+yt/sPEipghp9puvXIdNB4chE6jXMXlfMVy9k9crHYrYgSmxC5EUMBbhzET3hxUqOIoDCA2HC7XYbYeyY72xC2fB73UVIFxVEmrAcOKmXxG2Lhbd5D7NvvdoxgQ2bggbudW8oHIVOaRYZcbsL1pE3jkWAmJtCPOK9+Hwd1gbTP/lR38aNmhUh23JZVUgw54cKhlRQhTgmkOP3xINhxOv89PdAz4h2vG50aSIgAiIgAiLQnghIsGhPs6lrEQEREAEREAERaI8E6KTkLn4n/REdlhQpuKufBbSXwOjcd5ykFC2wQ9+kcsHi23RU8d98Tn0L9uNEWPC9RYUKTlhazQqmfzoCVgyjk5bX9RWsDEaxorW8OCdMV8U0W5wLRn7MSnLOaowUi1gUF37qsNfv2eh2mz7ssN7kcpsbI+HYEjtqxKJu5H2KRKuwUTri89klyG1fkRfwUtyw8nJ88RSGW507E+EkqwGrcSYEXBCbEC1jVrmQ5gue5whuSGgQdiek8IrjpiuHYJHH8iTYMR/CZz7cr7lYA9gU7/L5fK4CpAMrj1jxLn6fe2YoYgchXGibfCbk236bRBQdRKwcrIuuEC+6uky7i9fjznNDvYwbibVSZhsQKSCM4QEZwFNyOJ89KL5djDopBqMt8F3vssr4imjUinTvglIpEiza/srQFYiACIiACIhAByEgwaKDTLQuUwREQAREQAREoM0RcGpLUGBwak3QYcl/v/E7RhswLRTrJbCANl9sRwc6s0NhM/eWHbV09DMig07/pTBGAbAWBD9jn9WKFjc+N9OEs8wBV22bRkwbxR3prMFB8YVFtZ0i4wvx89ewn4kVLeWETym03QNjYk2NebDVMIo/2aSCcrgm3pMRLtGHpswvD1ZFInBmBzoVBgK5OT5jdfHmWLQ85PX7PWanApS5sIzNubm+eO9uBRYKOzspw37Wn35pHQSwK56VZHw2Jg3BMnHk7QkyzQ/EBzfuuhhCK1CL28QcWn607MzwKNyOXqT/6QGnM9O8lcAx3R03c9AyUAVDERatY2KbcBSLlm0wOhUEXHgGWFg/eGbbEQhbVRaewFhOfGb3MFn3xLDXsOA2FkVnLJr8qGVDH3O5I5GIDynEgjm5XttCJA9TjWGdtbgw3YTI1LUIiIAIiIAIiEA7IyDBop1NqC5HBERABERABESg3RGgk5KOcDrwnbQefGc6J0ZYLIVRqKCywM97wvhvvO5wWvFzOrTp5KLDnwW6mUZqI/yiK7CDN+L1ePx+v8t724uzsZnXiGGHtxmzLBccZTGIFY5owjE05YtRJL+ADYINhB0G+xR2D2wxxInWlreffJmei4IR6wpwHrYwaoiYctp+o+KItuB8hboU5brzcr2e3l3zzfUbK61unXO9PbrkG9hxH0FUhZPey8L5mnp+mnLu22PfiagmiA35iJawEF3BkAoTARcUEr0IgYpAvCjH/ceaFhTqIFDhJ5cZNeNm1I5bOfgU5UpQt8RwhxCgkWsbLtRftngPK61Pe1wxP78msyocS9QkwmPfxFsZ9IYSZPrrhEgLLgxkhrJ7QNrC3wST6wxtoIExAgeVtvEw6IK1Fs/1e2K5Rf7ObtNYjboWEiza/7rRFYqACIiACIhAuyEgwaLdTKUuRAREQAREQAREoK0SqCNKIZEuKO3a6LR0UkNxdz9fbLMGxnoKNL5YY4GFqilUVMAYBbCW+c+5s9vrdfngQh0QDEUhVCBljW1Xxm3mQjficHtt2bnfFPUtUlIY0fG/H+xUjg1GQYVFtW+BLU1eV6uY2pQx0/lHrj/AShsqGFSTzsmZb75zHjjXPCcd1k7kiUSKVrEqqh1EIqUPHMibYrF4vuF2b8Rm+W6m11iN+8wP9zJqDkCkQHoobJnPRzH1ErfhCsIX7TFdcDqbriBqWCxj0WQUW96Ayt3FFZXhaDgci7DmSeu9bI2skQjYKJKNoAqTz/k4hIkyBE4Uokh737hl9rAhKEPhDeAZ3gviVzz20xMihnYR6F6W120WoA5KFGnlgtForHJzOBpbv6FS6cQaaXLUjQiIgAiIgAiIQNMTkGDR9Ix1BhEQAREQAREQARFoEAFHMEgKF47D2om2oCNqFR1bMNZ9oNN/HYzpn5geaj2MtSD4774InFp0mq7HjtxcOFQLEVYRhFARQGwGjjexdRe5alwmnaKJHfxNLFbk4Bzbwg6Esdg2x8sUVzfBlibH0CB2jXVwiqjgFD0mU0Z+NLiuRh0RGU6UCy9Fu+vrOaHJQtg/O7op1nbyBE40FHzLdp7tssvgXP4BtQU6mx5IFAy+sKzBiJjwQJAIuj2uVSigXIHIpn7MCIXq26xNYEfgtM7J8VZ5PO5yv88T6t2d+qNeHYQAloNdgggdiqJMIZYPUSIMK0NNFFZo38i6FtGojeo21hqkgsrH2oliHZWgLfQu9yqklltfXhnZhOd5dPjAriafYXjWKNKigywgXaYIiIAIiIAItGUCEiza8uxp7CIgAiIgAiIgAh2CAJytznU6OezpdHJ2WlOwYPTEChiLP3PnP0UKpiqih7MURgdqIm0RhApoFFYxdu8irsLczIT5MDecXKgJbIQRWVEVjyf6tprCoZvi+Ge6KkZW7ACjWEGhZRnsPRhrWLTmneTkz2iV1jzGDnFv8CJT7o/qrtkRmCjw8eXMmQvHpYpB/K4x67TwfLw3Gd20ye9358ai1rhcny8f2XuKwiFEEplGJRzL3VBg243bz4b8xTRAKKJsRlF4vSLH9K70ezxrC3O9lTk+N1NCydncMVY155lrB89iazPELjMes1wogrIOq4QCaW4kFgtDoKDA3BurFsvIhTR/Rl48FkdEhiuMDsI5AR+EDdNXkOf3dS3KZZo5CZ4dY/3oKkVABERABESgzRNw/gHf5i9EFyACIiACIiACIiACHZVAcvc4N6JQBKDznzUhOtGxBWMUAJ20jLhwCnbzZyflkxNNkcAHkaLJnFopYgXz9u8CuyE5zu/w/gaM77NgW6IWGlIPoqOuB113QsTgPcAX1zfFg1RnP3/mfwc50Ups56Td2koUqE9heZyf9xrHwLVehJoVhsdjDvB7PQPhXC5CWqiBEDCGuF3uPJfLDrvc7oUoxt0NoyhkkeSAz7sc2+SXmi7ju0DAuwI/Vx44qW9rq+WipdZEBLB+EnVQYAUQJgZiTQzCWpiE92GMoMAiDaHeUA6E5y74LOTzeTZDvChE7aEljNbJCXgXYt3MxHcrkPavsme3/BDWT5M925sIg7oVAREQAREQARHooAQUYdFBJ16XLQIiIAIiIAIi0H4IMBICDi4KEHS20inl1Figs5Qv/u44OxN50ZOfN0kURXVk01IqbY82p8DyYcthL8CmwliDo1GKV7ef2dWVZEogKdw5QoQjzvHw6tY57xk6hZ30TYl2/L9GiixyoqF4D/aAMxllj93YIW8xoKl3AIUpoi4rF/ViEHFhxFGPe7PX6w6jZnI4N+Bdjl316wyXXer1eio65ftDnQpzVIMg04XQPto5z/IqRN1UIAyuBLFwi7CoUOoEwjSqsCNVWHeIGKWWZbhQ3wQRX/Ymr8e9Fgtls8/rqkD9isQzv3NhTry8kkEXeomACIiACIiACIhA2yDghEa3jdFqlCIgAiIgAiIgAiIgAtUSoJMVRqdmGMYIBaYsYp0FpotiOhB+5tRcoAM33kiO2WxmhM7hHrCDYJOT4/oA7x/CWDxcYkU2NNU2nQDXF6MaaE5anRrXebKAtRNtQYGD/23EVFGNFYXO9cz7j+nOkN0nUdR+WSgcXVlZFVvgNs0vEHUx2+NxlWOnfDcMJOJxu5ehXsU8yCjzAn7vcp/XXYqIDEeE1Ix3EALJZ7MjWpQjqqIUwsVCy7J+wM8/YH2sgnSxgSmj4vE40/5VYp2sh8AVK8jzrUfkzgoIXz5EWiRSk/12tyFKX9dB1o4uUwREQAREQATaAwFFWLSHWdQ1iIAIiIAIiIAIdGgCaTn80/Py0/naEuLEljlJRldwHJ1hg2H8N6hTd4ORFczzrx3AHXoVN+zikyKDI1Q4Dv4611QyOolinnPfOBu6GpQ+h2IIx0RhEO8UDtfCuWyiEHIAu+BRY8bOjbiNCogWeaGY5TFtuzNS/6wuzAtsqKyKrDYNexUiLpDNx46iBkEiuiIlSulnsJQ2rWFrp6WPrqUGC0UGisxM4ReBUBGCsLUQtSp6wEwIYBaiLgogepUh5VgFvo/iowpUsdgQiVrrPTFzE+qelAd8HokVLT3JOr8IiIAIiIAIiEBWBCRYZIVLjUVABERABERABESg9RGoI8d+nU7bZroi/rvzYNjEpBPufby/Sj8sHK5Kd9NMk9COT+OkgnKEh2zXPQUKR/Bww4ncKOnSkkIKo57odKbjuADVs8OWZW6Mxe1obq53vQ8Fk6vC0ZGIplgKR/S6SCTO4tuVeZYdi8Fwf8jh3I4Xbl3Pb6whpw4RAixsG8JWFeS1mBW3Q7Zh98UntuWyKiFObMLaWorIiqjb49pcGYxU+Lye+KJlG7K9F9oxbV2aCIiACIiACIhAWyAgwaItzJLGKAIiIAIiIAIiIAJtmwAdwRQq9oTRsTwjafPxLrGibc9ti48+KQo4hbXp3K+Pg9YROlhzgv+NxAiJBkUmOSnX2A/6YxQHx8b1no/d8aviVtwbDNplqEWwEcWS3ZbbXo/a3NgdH/dDsKCTWql8Wnx1tYoBcP04ayeEtVEGsctEtAUid8zVtmF5Y3H+apQi0qIYayvqto0o6p5E1xSXN4rw1iooaBAiIAIiIAIiIAIdhoAEiw4z1bpQERABERABERABEWheAimpoPrgzENhX8O6wpASJ1Fgm3U29BKBxiDgCA4NiUagY5j/feREa/C9PuJH+vWwDwoWFO42wfwwnisUjVleGMWJEjiig+s2VCA7lBGDaGFrZ3xjLIu234dTzwLCF9cR1zcjdjyItmCh7bWm25XDq8SX0VAkFkQSqURKtBaoUdT2YesKREAEREAEREAEWgUBFd1uFdOgQYiACIiACIiACIhA+yKQIlbk4cpodATTMRuEfQFjIeLGcAa3L3C6mvoScJy59T3eOY4REE4NDLORCnA7Y2PfrN1C0YIvOp4pZPDFegOV4Ug8CrGCQl5iDLXUN2joder4NkaAAgRroySLxXPdhGiojYIIHWsT8oeV4zunHksbuzoNVwREQAREQAREQAT+n4AiLLQaREAEREAEREAEREAEGpVASnFg7ijvBfPB+sO6wd6AraYztlFPqs46OoH0YvP15cEd7BQLGF3RmK/U8Tk/U7BwzpM+ft0fjUm/DfdVg2jF9UEBLHX9GMm2ibXjHFdHjYw2TEZDFwEREAEREAERaK8EJFi015nVdYmACIiACIiACIhAyxKgI20CbA/YchiLDk+HfQ6jQzjxQkHhlh2lzt7mCTRy6pt0YaGx+VAQSU1blS6MSKhobOJtvL+6inK38cvT8EVABERABERABERgKwISLLQoREAEREAEREAEREAEGo1ASnRFd3R6EIyRFaNgS2HfwLirPPGSWNFo2NVR4xLgzvVGS50rh3PjTo56EwEREAEREAEREAERaN8EGu0f4u0bk65OBERABERABERABEQgCwLcFMNC2/Ng5TCGUTwHc3L3S6zIAqaaNjsBRjk0dkqoZr8InVAEREAEREAEREAEREAE2iIBCRZtcdY0ZhEQAREQAREQARFohQRSCm3nYHhdYYyuYAHhj2ArYUp30wrnTUPaikBjFfAWWhEQAREQAREQAREQAREQgSwJKCVUlsDUXAREQAREQAREQAREoFYCXny7E2x7WB6sGPY2TKmgtHDaEgGJa21ptjRWERABERABERABERCBdkNAERbtZip1ISIgAiIgAiIgAiLQcgTSalf8EiNhwe0FsE9gK5yRqW5Fy82RzpwVgUTx7UYu6J3VANRYBERABERABERABERABDoiAUVYdMRZ1zWLgAiIgAiIgAiIQNMQ4GaYIhijKcpgm2HzIVJYTXM69SoCDSdQQ1FsRVg0HK16EAEREAEREAEREAEREIGsCUiwyBqZDhABERABERABERABEUglkBJd0Q+fHwyLwWbBvoSFREsEWjOBq5/kMt3qlSi6rQiL1jxzGpsIiIAIiIAIiIAIiEB7JKCUUO1xVnVNIiACIiACIiACItD8BNw45XiYL3nq+XgvgSm6ovnnQmdsGIGEWKGXCIiACIiACIiACIiACIhA8xNQhEXzM9cZRUAEREAEREAERKA9EijERfWArYUxwmIpbEuh7fZ4wbqmdkuA6aBMRVe02/nVhYmACIiACIiACIiACLRiAhIsWvHkaGgiIAIiIAIiIAIi0EYIMGp3LGwQLB+2BkbhQi8RaPUEVMOi1U+RBigCIiACIiACIiACItCBCEiw6ECTrUsVAREQAREQAREQgSYi4Ee/w2ELYEynsxim6Iomgq1uRUAEREAEREAEREAEREAERKC9ElANi/Y6s7ouERABERABERABEWg+Al1wqqGwKthK2I+wRO2KbfszU5ReIiACIiACIiACIiACIiACIiACIlA3AUVY1M1ILURABERABERABERABKohMGvFZn7KiArWrugM2wM2AzZNwERABERABERABERABERABERABEQgWwISLLIlpvYiIAIiIAIiIAIiIAKpBNz4JQDbBCuDvQ+Ls4GiK7RQREAEREAEREAEREAEREAEREAEsiEgwSIbWmorAiIgAiIgAiIgAiKQTsCHD5bBlsLehW0QIhEQAREQAREQAREQAREQAREQARGoDwHVsKgPNR0jAiIgAiIgAiIgAiLgEPDihyiM0RUUL2yhEQEREAEREAEREAEREAEREAEREIH6EJBgUR9qOkYEREAEREAEREAEOjiBZP0KUuC/J0fBusNijmChdFAdfIHo8kVABERABERABERABERABESgHgQkWNQDmg4RAREQAREQAREQARFIEGDBbQoV+TA/bJ0jWIiPCIiACIiACIiACIiACIiACIiACGRLQIJFtsTUXgREQAREQAREQAREwCHAemi5MEZWsI5FWGhEQAREQAREQAREQAREQAREQAREoL4EVHS7vuR0nAiIgAiIgAiIgAiIQAEQ8N+TrF9Bs4REBERABERABERABERABERABERABOpLQBEW9SWn40RABERABERABERABHoCQQ6MURbljmCh+hVaGCIgAiIgAiIgAiIgAiIgAiIgAvUhIMGiPtR0jAiIgAiIgAiIgAiIAAkwumIirBusUkhEQAREQAREQAREQAREQAREQAREoCEEJFg0hJ6OFQEREAEREAEREIGOTWAhLr8EFoBVdGwUunoREAEREAEREAEREAEREAEREIGGElANi4YS1PEiIAIiIAIiIAIi0HEJsMj2i7B8GGtY6CUCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiAC9SbgrveROlAEREAEREAEREAEmpFAXn5B4aAj3J9uAAAgAElEQVShI0YWdercpXxz2SbbsqxmPL1O1UYI9B80ZNjE7XbcZeTYbSb27N2nn9vj8ZRt2lja2obftVuPngOHDBvh9wdyuJ5b2/hSx9OlW/ceVcFgZWseo8YmAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAk1OADpF0dV3PPjElz9uiMxasdmmTZu3quyPF152tcfj9Tb5AHSCNkHgkKOOO+nlj76e76yR1PcP5/xY/OdLr76JIkFLX8zgYSNHP/LSO9NSx/fmZ3N/POiI357Q0mOr7vxjJ0zafubyMmv8ttvt2BrHpzGJgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIQLMQMPG6/5nX3ps2b/Xm404767zho8aOHz9p+53+ctk1N3+9dGPs5gee/G+zDEQnabUEuEauuPmehxwh6+Krb76bzv9JO+yy2y577L3fYceceNqt/3n65S9+KAlTuNhxtz33aamLYaTCezMXrXlt6uxF+xx02JFDho8aw/Hc/vBzr3H8x576h3Nbamw1nZf3Hce2w6577NXaxqbxiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiECzEdj7gEOPoLP0V4cccXT6SQ8/9qTf87sDDz/6+GYbkE7U6ggcecKpZ3Id/POWex/Oy88vqGmAFAdeeO/zbz9buK6SUQ4tcSEX/eumO2csXl/Vq2+/Aennv+bO/zxJUaVv/4GDW2JsNZ3zylv//Qj5durStVtrGpfGIgIiIAIiIAIiIAIiIAIi0D4JmO3zsnRVIiACIiACIiAC7YHALQ8+9RJrERyy6zZDbbzSr+nhl6ZMDQRyc487cLfJ7eF62+I1FKKoyOSdfrEH60Vghuy1q1cs/+zjD96JRMLh9Ovx+fz+idvvtCvrTODHQGlJyfovPv3o/Y0bSorre+2vT5uzeGPphpKTD9tnF5Q1qbWuCc/7/DufzXn6oXvvuOuGK/9R33PW5zhGgjDC4+P33n79ir+cdUp6H6zR8t7MxWteePKh+2791z/+Wp9zNMUxz7w9dWZhp86dD9p5XKsSUupzrdmsVc4Xnz0jx4yfmFdQUFhZXr55ztczpi9dsmhBfc6tY0RABERABERABERABERABERABERABERABERABNo4gf99MW/F7Q8/+2pNl8EUOl/9WBpF3eKcNn6pbW74rB/C1FwzlhSH0utG/PXy625Nv6BDjzr+5PdnLVmX3pYO8fpefE5ubh77O/VPf/17pn2MHj9hUm5eXn6m7RurXb+Bg4dyrCec/sc/19QnBTrWt2iscza0H5fb7WZEyI3/fuz5hvbVksdnu1aZdu75dz/7Jn2tfr1sUxwldTq15LXo3CIgAiIgAiIgAiIgAiLQ3gl42vsF6vpEQAREQAREQATaLoHOSEMTx6umK3j5mcf+89Vn0z4Kh6qq2u5Vtr2Ru/Bi/ZA99j3gkCUL53336nNPPrJm1Ypl0AEKOnft1v3dN15+IfWqTvrDeX87/5KrbmQkxYN33nj1kvnz5np8Xl8nTPCC776dXV8C4VCoKhaLRl2my5VpH/O+nVNvgSTTc1TXjmuZn9e2nm+47G/ncGd/Q87TmMcOHjpilM8fCHw3Z+aXjdlvc/aV7VqdtOOuu//7qZenYEm5Xnr60QdnffnZNCyxaFGnLl2CwYqK8s1lm5pz/DqXCIiACIiACIiACIiACIiACIiACIiACIiACIhAKyHw7tcLVz/+6vuftZLhaBhJAr8/52+XcPf5ZTfc+QAdwrWBYfHrmcvLrCde/3BGEbz2jQ3x8dc++PyOR55/vTH67dm7bz+KMI3RV3ofA4cMG0Fm5178z+uaov+m6POAw446jmPebufdftkU/TdHn9msVWQ36/LerMVrP5j9w3pG4jTH+HQOERABERABERABERABERABERABERABERABERCBNkLgvqdffXf6grUVdTnF28jltIth9urTrz/TQN3/7Ovv1xUNwHljoWumgmLkRVMAYPH1r5dujI2dMGn7hvZ/wRXX3/bx3OWlDe2nuuO9Xp+PBb/veeKlt5ui/6bo8y+XX3sL0yDVVsy8Kc7bWH1ms1Z5zr9fc8s9FNe232X3PRtrDOpHBERABERABERABERABERABERABERABERABESgnRBgbQLu8OYu/XZySW3+Mi6++ua7v/xxQ6TfgEFD6rqYfQ467EjO30G/OeZ3dbWt7/cURR575b3pjMYZPmrs+Pr2w+NOP++iyzjeTsn0TQ3pq7pj733qlSkU4JhmqbH7bor+Hnrx7Y9f+uDL75ui7+boM5u12h1V47/4oSR8xc33PNQcY9M5REAEREAEREAEREAEREAEREAEREAEREAEREAE2hiBYSPHjKMDmTvf29jQ2+VwWeR62rzVm6+46e7/ZHKBjMJ45eOZC1i8OZP29W3D6A1Gcny+aF2Qa2X/Xx957Mix20zMtr/DjjnxNK63vv0HDs722EzaH3PyGX9i/7/81UG/zqR9tm3cHo9nz/0OPoyRBdkem96eQhDn+l+33vdoQ/tqieOzXasUq776sTTaVHPfEgx0ThEQAREQAREQAREQAREQAREQAREQAREQAREQgUYmQEf0W599t7SRu2233XXr0at3l27dezTFBR54+NHH0+E+evzEyXX1z3oQTK/zuzPO+WtdbRvyPcWQg4747QmvfjJrIceWapdef8f92fR93Glnncfjuds+m+Mybdu1W4+eTF911W33P5bpMU674aPHbVPXMVff8eATHP9N9z3+s6LndR1X3feOWHjU735/Vn2Oz+SYQE5O7oDBQ4dn0jbbNtmsVfb92tTZixqrFkq2Y1V7ERABERABERABERABERCB/ydQa5FEgRIBERABERABERCBlibw1svPP9W7X/+Bbbnwb3MxZE2Jh//7v0+4k78pzsnd+0sXL5w/79vZX9fVvxNFwPmrq219v2ckwZMo5v0vCACL5s395u9/OvW4s4779a8euefW67+c/smH69euWZVN3/sedPhRvLbidWtWZ3Ncpm03lKxf9/m0j97bc/9DDs+mLgQFmWf/N22Wx+P11nYuR6j6ccnC+ZmOqaZ24ydtvxO/mzv7yxkN7aum4y/61013NlUKpmzW6tARo8f2HzRk2FsvPfdkU12r+hUBERABERABERABERABERABERABERABERABEWgHBLgrnTUTbvz3Y8+3g8tp0kvYZvIOO3OH/d4HHHpEY5+IkQxTv1+56a+XX3drJn1zt/ozb0+dmUnb+rQZPX7CpPdmLV7LlFP8uT59OMfw2v72zxtuZ/RDUwtje0Gs4BwdfeLpZ2c6Zta+eP7dz76pqz3TIA0aOnxkXe0y+f7yG+96kCm2mGYqk/bZtvH5/P5p81aVUbTI9ti62me7VhkFxLkvLOrUua6+9b0IiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiEAHJ3D9vY88S9GC6Y46OIpaL/+M8y++nM5w1nRobE7jt91uR/a9x74HHFJX33Ryfzp/TflfLr/2lrra1ud7RhK8N3PRGhaEbsi10mm+36FHHvPi+zPmsn7BoUcdf3J9xpPNMWQz5cv5K5nqLJPjGFUxY0lx6O/X3HJPJu0bqw2ZPPLSO9Maq7/0fibtuOvuXE/7Hnz4UY19jmzWKs99zxMvvf30W1PrjBpq7HGqPxEQAREQAREQAREQAREQga0JKCWUVoUIiIAIiIAIiECrJ/DC4w/9m47bw4896fetfrAYYF2pe7gTnkWNM72WTl26dmP0RK++/QbUdsywkaPHrV65fOnGDSXFmfadabvtdtl9T7ad9+2cOqMmxmyz7Xa5eXn587+dXWfbTM+f2o7RELl5BQXnnnL0IfW5Vo7vkutuv48RGtff8/Az4VCo6qTD9tnltReeerQ+48nmmHgsFnvp6cceZI2ISTvssltdx7LGA4WVubO//qK2thRxBg0bMaqu/pzvff5AoKa2+QWFRUOGjxrz7eyvsk4H5UdhinETJ+/ANEu1r9Ux4/j93Nlf1XpdmV5Parts1ioFpInb7/yL+XObZq3WZ/w6RgREQAREQAREQAREQAQ6MgGzI1+8rl0EREAEREAERKDtEHj5o6/nB+AMPWiXcYMtvLIZ+e777H/wb44/9UyKBHded8XFi+Z/t9XudtZ/+Net9z363GMP3FObc5i1ByorKsqrOz/T/fzhr/+4cvioseN/WDT/+z/+7ogD1q5auTy97euffrPk3TdefoFj4Xes9/Dbk8/4IzLSdPng7ddf/s9dN13jHHPKH/9y8R8vuPQqJzXP+2+/9tKl553+u1BVVZBjvuCK629jGqBIJBzeFo7XOF6zvpg+lcfH4B1fMPebWY/ce9sN1Y13l1/us/8Rx518+sAhw0agvMKaf99yzRXffP3FZ2w7cfuddj3oiGN+hyF15XnGTpi8fc8+fft/gPOn9kXB4PH777r5qBNPOws1JQaQcZ/+AwexMPdXn039qGxj6QanPcf84J03Xr3sh8ULs5m/1LYsPv38O9Pn3H7NZRc+dt8dN2XTD/leeeu/H9lj3wMP5XFffPrxBw/dfcu1X0z76P1s+mloWxYkf+uzuUv/99p/n73k3N+fkN4fIwTO/PPfr+BcMk0R58JhaeMVDFZWPH7fnTcvWTjvO+fY2x9+7rUJELX2mTy8N0WR6sbINXTKWX++6JhTzvhT1+49e82fO2fWWccf9qtNpRtKUtvvssfe+93z5Mv/u+bv5/9h1LgJkxgFwXm+9h9/PovMarr+nXff61fX3fPIM+TMNrzPLjjjhN8s/3HJIv5+2G9/d+q+hxxxdDQSiXDN0Zz1xHu6dEPxet4TwcrKivRzUEA5/vdnn0+xKRqNRl584qH7HIEpm7V6+7WXX3TsKX84Z+jI0WO9Xq8vB8oa7wOyZH0W57xk//qLTz827YN33mrofOt4ERABERABERABERABERCBzAlkvLMv8y7VUgREQAREQAREQAQan8BLTz/6ICMMdt1z3wMy7Z2RDlfcdPd/WE+BosUv9vrVgaefd+Fl1R3PXeEHH3nsibX1ffUdDz7xwHNvVuuwPfms8y+85cGnXqqCs/XZR+6/q9/AwUPpdE7vj87cfgMGDXE+P/fif15320PPvDJi9LgJvfv2H3jy2edf6ERosDbDORddcS18qd/ce/M1l9PBzPoUx5129nk8HvpN7uhtJk6mE5uiQhHEBTqze/cbMJA78wcPHTGKjun0MTDH/2U33PkAU+FMRmqe0uL168ZOmLT9vU++MsVJu7X7Pgccsg0KL/fq238APyP7ivLNZaPGT5w0Dg51FmUes82k7br36tOXv+/4i1/u03fAoME834DBw0bApxyhY95py3eOqa7ok7rm9hDMEQWjF5986L662qZ+T1HnCRTo5nVSEFq/dvWqcRO32wHZs3pm009jtF23ZtXKaR+++/Y+B/36SM5Zep8jx24zMQ9hDmSIEi69YrFolJELXFMDcR2DhgwfiaX9swLcLBTOSBzoaYXVjZFRGnc99uKbZ//t0qsQODGd9xPEiG1PRP2G9PaM5uFnZ0Mow5oc8Mqzjz/ENXA57iWus+r651q86vb7H6NYcv9t11354ZQ3XqFwd/HVt9zttGe/0Ey8UYhr3Xv27rN508ZSri8WvGZ0SL8Bg7fcF6nnYGTVc+98Opv3ZyUWYdfuPXpSeOI9zXbZrFXeG3sdcMjhFEt4TRAuEpEe5EtRjuuaRkEjF+pkY8y3+hABERABERABERABERABERABERABERABERABEWhnBOiMZZ0BigKZXBod49x1zjz59z/z2nvcmX/RVTff9cHsH9b/8cLLrk7v47RzLvjHR98sLakpVRN3mbMvFiNOP5YREvzuqtvuf8w5/uYHnvwvIwHS2+6538GHsS13o//u9D/9hT9fffsDjyfSREFISC38e+GVN97B7+ncZT9sc8O9jz7nOGpT+2Z0BdtW9136GP586dU3OddCRzO/Z0QEPzvxzHMvSG9P4YHfnYXokUzYvz5tzuKHXnz740zaZtvmrc++W3r7w8++ms1xrHPx9uffL6NAQyGAxyLrUSeui6+XbYpnUpcjm/Nl0tZZB8ee+odza2vPMT791idf1dUni1czxVVN7ejgn7m8zNr/10ce67T5zwtvfTRj8fqq9PRQ9z396ruc72NOPuNPTluue35WnQDGNk4x8QMOO+o455izL7jkX6efd9FWAiEjPXjev1x2zc11XRfXM8/7+GsffO6kRON9wGu989EX3mjoWqWgyfo4CLbw1TUWfS8CIiACIiACIiACIiACIiACIiACIiACIiACItDOCXBnMx2bmeTfv/epV6awADGdzXVhufT6O+6no5O1ChwRgUIFP3v+3c++ST+efd/9+H+rTf9CIYEpqXgsIzFSj+VY3p+1ZN2z/5s2K9XpWVMh34uvvvluOmu5i5sCzCXX3vbvmq6Fggvb1HWt/P640846rzaHstMH0/3Qcc30V+n9slD2tXc99FT65zvsusde7HvvA3/9m7rGQqHo66UbYxSH6mqb7ffky7GzuHimxzIi4MHn3/zwyTc++oJRBqnHMb0XBZC3Z3y/vLEc1siKNYiCUG01IjgGjmXavFVljPqo7Vo+nru8lGu4rut99OV3P2UkUXXtGJXD+WM0T+r3jHj4XVqEBcWE6QvWVpBZattr7vzPk+yDwmF153DENwpndY11xJjxE9gXC57X1pZC3Ydzfizm/cq5Sm3La33nqwWrGrJWeexD//3fJ5kWQK/ruvS9CIiACIiACIiACIiACIhAwwkoJVTDGaoHERABERABERCBehKg0/bOR557nSmOXGbdRahZ94HHMLVTbac8+sTTz/7N8aec8eZ/n32CefeZH5+O2AMOOzqx+3v6R+/9L/V4ChpMfzSvhsK7B2BXOlMKLfz+2znp9S1O+sN5f2PBY+b7Zwof9stzDRs1Zvyi+XO3EkYm7/SLPZiSh9ET3876asb1l//tnJquhSlz2JcTYVHbNTO90ZqVK5ZtKF5X4y57igmXYac8C3Nfe8mfz07vL1hZXu7UH0j9jqmc+PuieVtfT3of/QYOGkKBJ5O22S4bZJvqQwEiveZCbf0wooDMr7ro3DNY5yO1LVNLvYDUUqi90X/yTrvuke140tsjo9fgh1+aMpVpy+w66qxwLB+/+/brFMBqml9yZ8TNtzO//Ly2sXFemT6suna8Xy745/W3Mw3VA3fccFVqP6xX8sQDd92S+tnIMeMnMoLhuccevMf5nH2wQDhrj9TEvgxrle3rKgzPNo7o9+3ML2q9rr9ece2tvP5Lzvn98el1Y5D5rMFrlWNBlq3hi5ByraFzr+NFQAREQAREQAREQAREQAQah4AEi8bhqF5EQAREQAREQATqQeCKm+95aNy22+945jGH7MMi1XV18dnH709hmx1+8cu9a2rLXeMXXnlDQgz45wV/PI31HdiWqWroUObP6UWWWdCXqYKqc1xSMHB29L/9ygtPp56X0SFHn3T62VPfn/Imz+d8d+hRx5/cA7Ud3njxmcdT26O+b/7QEaPH0hE9cuz4iVf+7Y+n1VQgmcfNmPbhe3zfbe/9DqqLzaQdd9l9ztczptfW7sDDjz6ezvm7b7jyEhbATm+bk5ufHw6HQumfD0C+/wg+X7nsxyV1jYO1AdgmtSB0Xcdk+r0TKePz+34WKVHb8UeecOqZs778bNqC776ZXV27T1FLgp+P3mbbyZmOo7p2dPLfjZRTrLFw2pEH7OGIV7X1Of3j95LreY9q1/Mk1Bfh8XXN66hx22zLiI5vZv5UMD31ddgxJ57GOb/npqsurW7O09tjHe1moeD0Z8mx8fvTz7/wMgoRLJhe0/WgGPf7vNd223v/DNbqrruXrF+7hsJZTf2xXse+Bx525Muon8Hi3Vuv1Tys1XCD1iqjNpjiqinWakPWko4VAREQAREQAREQAREQgY5MQIJFR559XbsIiIAIiIAItCAB1oSgA/1fF55z+ndzZn6ZyVDWrl65glEEqE89qbr2FBeYCioUClX940+nHsdixWzHHf9nJHPp06maKi7w+zHbbLsd3yFYbOUY/fXRJ5ziRBhQmEg97577HXQYU0I9+8h9W9If7fLLffZn2qfXX3j6sS+nf/KztDrDUISYEQJ0ILPo8dIlixbUdt3vv/3aS6hzvYlO99raMQ1Ros7EF59Nq63dSWed9zfye+eNl59Pb0fnLa1sY+mG9O8GILwEWsUiRqrUNU9syzZLFy+cX1fbbL/H0Ep4TCEKl2dyLAUOpt6qbX2x+Db7KsBEZtJnTW3Ov+SqGzmv553y20OrY1jdcbNmTJ/Kz0ePm1jtemZUQ2lJ8XpGNtQ2Nop0FBnmzv7qi/R2rEPB8Ux59b/PZnJ9E5HS6cclC+c7EQ1MNfb7c/52yXOPPXAPI5Zq6oP35udTP3x3r/0PPpw1Q2o7F6+rrrV64pnn/BVBV67H77+z2joXFAQbvFaTkUNNsVYzYa02IiACIiACIiACIiACIiACWxOQYKFVIQIiIAIiIAIi0CIEzvzzxVdwZ/OU117MyJHqDJKRGAMGD0s4xdNfx55y5jnDIQrcdMWF52Hz9g/O97857pQz+g8aMow7zFetWPYjRYDUY4eOHD2WO+KXQ0FI/Zypduis5Wc8Jj0KZOc99v7VhpL16z6f9tF7FC7+cvm1t9z12ItvfvnpJx9QiEkfH8fGzxhV8ei9t99QF3iO99lH77+bBbF33G3PfWpqP3H7nXbld7O++MkBXt2LfTCS5L9PP/IAndvpbSim8LMfFm4d6cKoiR8XLZhX13j5PaMx6GR3UgRlckymbRi9UBUMVg4c/FMUR10vZDIKsDaFaZhmTW0ZOcLvYpiUuvqr6XumdDriuJNPf+2FJx/NJArF6YcRBpxjRxBL75/zyuiQusZFwWIh0nUFKysrUtuO33a7HQcPHzn6tReeejQ9HVZNfbIGxeIF389lNBALUl9wxfW33X/bdVdef+kFWwpw13Tso/++/UZGHVHkqKkNhYbe/foPnFnLWqXwyPoWM3BfLYdQlt4X55Qp2qCrbBWVldVaHTw8sY5+yHBt1zUP+l4EREAEREAEREAEREAERKDhBCRYNJyhehABERABERABEciSwLCRY8YxNdKrzz7xcJaHGiWo0cD0OxQTUo9lapc//OWSK+d9O2cmHbTOd8j0VHTWX/9xJWsqrF65bOniatLLcCwrl/64JD0906FHH39yl27dejB9DWtXOOmlnL6ZsmfurK+/OP3cCy9F4eZlFEzuv+36K8895ehDnOiO1DHyuvn7R++8+Sp3pGdy7U/cf9ctdNSfevafL66p/fhJO+yEJmV0NNfU5hd77Zeo+/H+W6/+t7o2O+221778PD0agdEprEuxDF7dTMZLh/HSDNtm0l96G6ZHYtqiTI6lGMCaC6x5wuuo7pg+uDh+vnbVyuWZ9Fldm70POOQIrsdXkL4o2z4oeLFOQ/pxRZ27dKXINufLzz+tq89ttt1hJ9RF2ardnvsfcjiPfef1l7aKqKmuT84d67EEArm5L7w341tGC519/GH73Xfrdf+sawz8nqnWZs749JPfnnTGHyl4VHcMI174+Zyvar6uCZN22JlMalqrFGj4DGiMtUrxLhuRKRMOaiMCIiACIiACIiACIiACIlB/AhIs6s9OR4qACIiACIiACNSTgFN097tvZn2VbRfYwJ3L1EQWPI2px570h3MvYEqjO667/KJUYeGsv15yJVPU/PuWa68YNHTEqOoiBVjbIj26gru4GV3x4pOP3E/ncXqBYAokyMQ0ZI99Dzjk9HP/dulH77z12uF7TB71wO3X/6u6CAaOlYW4+Z4qqNR1/YzseP6xB+9l3Y7ho8dtU117FgxnAeV0QSW17QQ4eYvXrVldUxoqFopmVMSctDoIZENnfF1piZxz0em9vI4URnVdc23fo1bCB9169OrtOL7r6uudN156nrvxmTarurY77b5nQqj56rOpH9XVV03fs+A5BSroRXOy7YPrubp6F5xT9jW7Fsc+vycLRizMrkbY2BFrhuvn+wzvs22Rqol9ck1v3FBSfMSe249hmqdsrumhu26+ltFGv/7t706taa0ySqY2VhQkeCznuro+uFb5+dT3//dG6vf1WauMcsmk3kg2DNRWBERABERABERABERABESg/gQkWNSfnY4UAREQAREQARGoJ4HO2MXNQ0uxuzzbLlAjYRgd76n1FLib+zfHn3omnfYzpv5UqJovRkAcg6gH7jAv3VC8njUNmBIq/ZzdkaZmTdoO+9+ccMqZFCqmfjDlTYoX38z88vPU45AFqB9/Z17/g3+xzdBLzzv9d6lpqKq7rhFjxk+gA3n6Rz8VD8/09fTD991JEeSwapzALLY8Ysy4CdXVL0jtf9CwEaPmz/1mVnXnZIQJ0wd9OOWNV9KjTJx0RXXV22C/dL4zPVImbTO99vR25E1x4Pjfn31+Jn3cetWlFxx/0B7bV7eLnlEXXDcUK6pLPZRJ/2zD9cx6CjUJVTX1w0LvnRHSgOW8Mr0NBRk60hd89221xcKd9hO223EX/pwesUCRietiJupkZFJ7JHG/JAULinqMcGBkT6YMnHbTP35/ClOnVbdW2YbXNe/bWV/XxoprlemtViz9YXH6+Zku6pAjjz2R99r8uXN+tp6zWavsl+2bcq1my07tRUAEREAEREAEREAEREAEUINSEERABERABERABESguQmEsMWa5+zS9SfhItMX09WMQMVtChOpx+x1wKFHULR48amH73c+5y7vf91236PrVq9acfXF553p1I9YvWLZ0tRjmXOfkRkb1q9b63xORzKLdD/98L139Ordtz8/T3eeou5zV37+9qsvPJNJOiHu8KcTmIW7q0sXVRsDpqTiThSpyqkAACAASURBVPfd99n/4PR2Q1CjgM7p77+Z/XVtfXTv0bM3+6mujVPU+8UnHrov/XtGTDByYykKBtQ1T6wtwqLi6bU+6joum+9ZJPutl59/at+DDj+K9RbqOjaMvFA1RRic8Ps//plO69uvuezCuvqp7XuuZ4pbFMSy6Wcn1CXhMenrmX1gnW+zZMG87+qqPcHIGaYXS08x1qf/gEFcF1jvWwl0NY2R4gfP9+CdN17NdFSZRrGk9/fGi888TnGOheDTv+N9WPda7dV7A1K/VRcx9Mt9DzyUUSUNXascF9d2U67VbNaC2oqACIiACIiACIiACIiACPxEIKv/qBI0ERABERABERABEWgMAk5aJie1S6Z9HnPyGX/iDus3X3ruydRjdttrv4O4i/xjpGVK/AMHO+dv+Pdjz1FsuPhPpxzLqAZn9zX83T+rHeHk2g8GK7YULD7j/Isus2zLQmHsG4eMGDWGfabvgi+EYsHPsQk+nMn4R42bsC3bffrhO29n0j69DVP+9Bs4eCgFltTvIFgkxleb45UighcVqJmKJ73fXn369T/smBNPm/PVjOnpNQHYdvCwkaPXIfyksqKivK5xsy3bZFqgu67+avr+ruuv/MdmpK/61+33PwYNKDEP2b5223u/g869+J/X/QfO+equO5v+eL0UB5CCqcbC6NX1x+LUjKJg2qr071kgHaVAtioqnd5uwuQdd2Fdj/TPmQaNnxXXIFKlt+/UpWs33iOs1fLOGy8/z0gkplPLhoPT1klP5aRAcz5nwW3WlKlLJEDQUE4VQizSz837+vTzLryM0RcvP/PYf9K/z2atMqUbRc2mXqv14adjREAEREAEREAEREAERKAjE5Bg0ZFnX9cuAiIgAiIgAi1E4Ivpn3xAJ/gxp/zhHKZ/yWQYI8duM/Gks86/kEW103PXj5kwaTum9IEusZHO+b9fdfPdO+++169uueoff3V2r2O3dyJSgsWpU8/nh3eUv4dDoSq+U1g4/rSzz78bTnGmxGFefNZ24E791OOC+JK/07ma2fjHT2S7L6dP/bCu9nSmcvd3ajsTO/GTpTv+r727jqsie/8A/t01dlfdtGtNFJBGUEHE7u5c1+7EDmzFFjtR7AQDFYsQRGmQFgQVCwNbsXZ/80HH3zjey70XLi7qh9fLl3LnzJlz3jPXP84z53k+qt0hFo3GG+lie8wBRYnF3/GmOmoSYIeK/Nqjp85ZjFROy+dNU1jUGzs41K1JUV6nkh4W4FEXQNUcs3IcO0WmjxncG/dm/R43Dyy2q9sfdjT06Dd09NKNuw4eP7hvp7oFpTPqHzs+cG9GTZm9EJbqjKV9jz4DkbJs39ZNa1AYXH4O6lJI7yl2/WDXgrQdUpXpGhqbKdqhge8B2v6kYDyo6YFnTNqXWDMj+IKvN9KCOc61H4/vkLj7RtoWaciwAwOf5RUCYWJNGrENnlX8W+jmtfQ87PrA79J5YeeRfCeGkL0tRdGz2l5I34X/B7asWbYA33W5mWbP6rvgmrq1WdS5p2xDAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKfKECVrb1GgVfefDmdGjCbQurWnUymkYVYzOLM6GXU/zibj/FgqW8rW/MjUebXU76YpF26vzl60OTH/87ee7SNdJ2SzftOojPkf5J+jne0Mfn7br16o9/HzobemnnsbNB4oLvul2HT+896fdJMWUs+uK8XkNGf7TQj0X0cTMWOMp3jyzZuNP1dEi8wpRM8vks3rDDxTM86UOAASlw3ANikp1cTvjI2w4YNXEaxiEuQDdr26l7yLVH/9Ss27CptO2qbS7HPcIS70gX1Ft17N4L505xcPyQSkveP9xhqs5jNn/1lj3wU6etNto0F2oZ4Bk6ERh7vV7TVu0y6hP3E8/c1kNnzsNnxKSZ8zVN4ZRR/4PHTpkFS/SPYuwZtYU7xu3iERiNQIS8LcaF45PnLUtP0YU2eCa3u3kFSNuaWFS3xjUVpW7C84BjG/cd85KegyDJhfiU572H2k2Ufj7IbtIMtK8mpKkSP5+zfOP2oKTU141atu8sbYtn7lzsrfSAXZfeA4fD09Lati5+RwBj5dYDx/Bdlc/NvHpNW1xD7A/pobwjr6WOnDxrgbT/XoNHjUc7fSPTquLnaItr7j11/iKuochXk2e1Q4++g3AN1FzRxrPIPihAAQpQgAIUoAAFKEABClCAAhSgAAUoQIEvXACL+liYx8Ih3pTv1LP/ECMhJz9SHyEggEX36YtXO2HxFouVimo4gMDVMygGC6tHfMMT0BeCA0gf89EiqBBYwLEVzvuPShc8sZDtFXH1/p4T58Kw2I6FVhShFs/FuBQFCnB85zGfYK+LV+41ad2ha51GzVtjrAGJ916iP/nb8G5+EYmL1m8/oM4ta9Gha0+MFQvamMvZqOQH5y+lPFO0MN24VfsuaDtvpdPOMdMclsJq+ZZ9bmLARbxe/Wat26MdFpPhiAX24KsP327af9xbnmZKPAcpcxQFZZTNAYartru6qzNHbbXBM3T8QvRVjNPVKzh26Dj7ObgfWEBH2icEBxC8Ep8NtBFqRzTQ1vWl/fQdNnZyYNL9V3gGHFY57ULwCLtdsIsAC+5N23TshgAYxnrk3MXLGQU2DnqHxCGY12fYmEm73X1D0ae8Zgd2P6AvfG8QtJGnx8K9wPEJsxetRLAGfSFYgX4RBJOOfZnTnsN4dsQUaTiGHRx4ltAHglF1G7do06xd5x6+MTcf7zruE4I22GmB7x6+xwvWOO/Fc472SHclN0ZwAMGNrYc9LvQfOcEeAbRj56OuiOmrxPYYGxwP+4TFN2zRtmObLj374nuGgB/+b1B07zR9VsdOn7/MP+HOC/n3JDueC/ZJAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKfCECWGgcOHridCxcYqFT/gcLrFgIxc4FZVPCQirersYC6PCJMxxQT0DeFjsLsMsAi5TydDM4B9f1ib7+EAu70nPFt8wV7ezA2+oIcIhjxkLu+FmLVsjT7WBXBxZqEVxQ57ZgEXX8zIXLcQ4WbrHILRYNl5+PuW5xPXUOY0B7LJQrSkuEPmc7btgmjhXBCvsFKzYoC1bgOoamVauhPYIdqsaN/hFUweK4qrbaPo75YscA3r5X9AxhIR6BJ/jLA1naHgvqQGBHCp4lRWPBMyqk4VokDQwoGgN2jPhfvpuGPk4FX7qpqN6LVe36jXEcAYPR9nMXy/tBWjEEMqTjwA4QsZ6LtD0COTuOegfK+0DQArtR8L0R+8F3VaxXgvbY6SJ+D7AbKaPnBXMX+0HAT1kAAimzcN/EtpsOuJ9Fmixl90uTZxV94P+C/Wf8I7V9/9kfBShAAQpQgAIUoAAFKEABClCAAhSgAAUo8JUIICiBt+LxFneD5m064I1yVQu7mk4dRbvl5yAFDwISitLzYAzY5VCwUJGiiq716+9/FMTCsZmllY20boS0LYIKbbv+3U/Tt7kR6FB3/gjCyNNdKRovAh8wzmjxVzxPfINfWbBE2r+YIqtzrwHDNL0n2mxfrGSpP5FiDMEJ7GjAv1HoWZvXUKcvBEZ09AyMEEzDjpnaDZu1QoojTQImqBWB4FdGqauq1rCpnVFaIzyTuDa+U3pCvQtlY0c/GdWTwXfDsmbtenjWFQW5ENjAd0EdG9wPdeqOoLYFnlX5biVF19DkWcX52K2h7o4ndebENhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKJCNAqihgJ0YWDhXdRnUJcDb8CjUrKotj1NA2wKaPKtifY9h46fN1fY42B8FKEABClCAAhSgAAUokDWB77N2Os+mAAUoQAEKUIACFPhaBfQMTcySryQmvHqZlqZqjuLb+/Gx0RGq2vI4BbQtkLlnNYrPqrZvBPujAAUoQAEKUIACFKBAFgUYsMgiIE+nAAUoQAEKUIACX6MAsvboGRibXYqOCFdnfpbWtes9uH/v7r07t2+p055tKKAtAY2fVSG1Fa59KTpSrWdbW+NkPxSgAAUoQAEKUIACFKCAagEGLFQbsQUFKEABClCAAhT45gSq2dSpj3oLoYHnfVVN/veChQrrGhiZqtNWVV88TgFNBTR5VtG3lW29Ro8epN5PSoiL0fRabE8BClCAAhSgAAUoQAEKZK8AAxbZ68veKUABClCAAhSgwBcpUKte4+YYeICv9xlVE7Cp26gZCoqr01ZVXzxOAU0FNHlWS5YuU65CJb0qgX5nPf8VfjS9FttTgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKDAZxTAjgn/hDsvDnqHxKlz2Z3HfIJRnLtIsRIl1WnPNhTQloCmz+po+7mLURy+cav2XbQ1BvZDAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIAC2STQf+QEeyzq/j1o5DhVlzCrZl0LbVduPXBMVVsep4C2BTR5VvMXKPCzb8yNR14RV+/n/eHHH7U9FvZHAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACWhQoWLhoMe/Ia6lno5IfCHW3f8+o6++Fny2up84hYFG1hk1tLQ6DXVFApYAmzyo6Gz5h+jw8qwNHT5yusnM2oAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAgf9OIHfuPHnW7Tp8Gou63fsNGaVqJIPsJs1A22VOuw+pasvjFNCmgKbPanWbOg2CklJfuwfEJGOnhTbHwr4oQAEKUIACFKAABShAAQpQgAIUoAAFKEABClBADQEEFZxcTviUrVhJN6PmWMTddsQzAAGI3e6+odg9oaw9CmyLqXhOBsXdKFSkWHE1hsImFMhQQJNnde37wNphn7B4Ic6WJ6OOa9Vv3Pxc7K0nCFhYWtvW5W2gAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKECB/0AAxYWDrzx443/5btqISTPnl62gU1k6DBTK7vx3/6EnAmOvI1gRKCzq4u+Fa7fuMzK3rIE32cX2CGrUb9a6/XY3r/TAxpnQyyk6egZG/8G0eMmvUEDTZ9Uv7tZTPIco+m7boGlL6c6JXLlz5zavXtPWYfXm3SHXHv2DYEXTNh27fYVsnBIFKEABClCAAhSgAAW+KoHvvqrZcDIUoAAFKEABClCAAp8IGJiYW462n7vY1KJGTRx89TIt7cmTx4/y5StQ4Kd8+fLjs7QXL57v3LTa8cDOLesH202e2aR1h67f58qV682b16+fPHr0EG+x/ywUtUDbf4Ufj+OHXRymjh12787tWySngLYENHlWN69eOr9b3yEje/QfZodgxT/Cz1PhuX775s2bX3//o6C4SygmIjxk7qSRgyLDggO0NU72QwEKUIACFKAABShAAQpkjwADFtnjyl4pQAEKUIACFKBAjhPQMzQ2q1mnUdMKunoGP//y229pL54/F+INNyLDggLOnjp+RFjrfSgOuliJUqVrN2rWWt/Q1PyPQoWLCGvAbx6k3rsbFxke6nPmxNEbyVeTctwEOaCvRkCTZzV/gZ9/sW3QpIWJRXXrosVLlUagQniUHyTGx0YH+HqdiQgN8v9qYDgRClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClAgJwigRktOGIeiMSCdoDbG9sOPP/1UtmIlXW30ldk+fv3t9z909AyMylbQqfyd8JPZfngeBShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUOCrE6hibGYRmvz4X9sGTVvmtMmZVbOuhbFZWNWqk9WxOaxy2rXpgPvZrPaj6fnf58qVq02Xnn13HfcJCbn26B/MB392HPUORBBF0/4+Z/ttRzz9B4+dMutzXpPXogAFKEABCmSHwPfZ0Sn7pAAFKEABClCAAhSgAAUoQAEKUEC7AoamVauhx9evXr7Ubs9Z7612w3dBFAQustKbgYm5ZaOW7TunPX/+LCv9aHpusZKl/tx66Mz5qfOXr0+5dSN51vjh/Uf37drmWtLleH0j06q6Bkammvb5udr/ImwHgRt3gnwucV6HAhSgAAWyUyB3dnbOvilAAQpQgAIUoAAFKEABClCAAhTQjgBSFKGnqPCQQO30qL1eTC2tbNCbkblljaz0OnSc/Ryc//TJ48dZ6UeTc0v9WbY8dnT8K/z0atuwZniQv594fjmdynpDxk6dfePa1SRN+vycbStXMTLB9S7HxUR9zuvyWhSgAAUoQIHsEOAOi+xQZZ8UoAAFKEABClCAAhSgAAUokOME8hco8HPnXgOG5cqd+8PLewULFSlapnzFSjlusAoGVEnf0PhG8tWkRw8fpOak8QrZkvKJOxCy8qZ/1Ro2tavZ1KmPuT1/9vTJ55gjnonlW/a5/fP2n7d/t25gJQ1W4PomVatbe55wO3jvzu1bn2M8mblG5SqG7wIWl2IZsMgMIM+hAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKPC5BRo0b9MBNQn6j5xgj2ujZsEBj4CoGUvWbP7cY9H0ehjrhfiU5/NXb9mj6bnZ3d7S2rYuXN38IhLxd7mKlfUyc03ng6f9xLoRdvbzlmSmD03PsV+wYoN/wp0X4i4F6fl6hibmMC9dtnxFTfv9nO1nLV3nHJSU+jpPnrx5P+d1eS0KUIACFKBAdghwh0V2qLJPClCAAhSgAAUoQAEKUIACFMhxAl4njh66fjXpcu8hoyYUKVaiZOtOPXpjcX335rUrctxgZQMqL4wThZ+jL4YG5bSxmlWzSq9bcWC70zr8bWRmUV3TMVrVrt8Y6aRiI8NDce6zp9mfEgrXQ5HttUsdZsRFXQyTjjlv3h9+mL5o1aZ1wrHkK4kJms7nc7bXMzIxv5IYH/f69atXn/O6vBYFKEABClAgOwQYsMgOVfZJAQpQgAIUoAAFKEABClCAAjlOAAu66x3nz8LC/7gZ8x1RL+Hwvh1briUlJqCOQY4bsGRAuobGZvg1JwYsTC1q1Ex78eL54b07tmCMmaljMXD0pOn/CD97nDesQh/PnmZ/SqiRk2ctuJqYcGnruuWL5Pd+ssOytQ9T799zXuu4MCc/F0jHVa5CJd1L0ZHhOXmcHBsFKEABClBAXQEW3VZXiu0oQAEKUIACFKAABShAAQpQ4IsWQFqlRw9S77969fJlvaat2mEyzdt27tGqY/deWCxvbKlX+m7KrZs5cZL6hqbmKAotBCyCc9L4cufOk8fIvFqN6IjQ4Pv37qRgBwvqWGgyRus6DZoYmlatdsrNdV/KzevJ7wIWT7K16LZZNetaCLRMGNK7y9s3b95Ix9tv+Lgp1WrWrt+1aS1zPBeazOVzt0UqKzzX4s6Uz319Xo8CFKAABSigbQEGLLQtyv4oQAEKUIACFKAABShAAQpQIMcJ1KhVt+HY6fOXldOprPfqZVoaBoiFarxdf/vmjeSI0ED/nBqswFhRTwG7AbJ7IV/TG6cn7PzAW/4RIYEXcO5F4e9GLdp2wi6Wl8K2C3X6w+4KBGM2OC6YJdaLyO4dFt36Dh6J4MopN5e90jG27957QJ9hdpN6t2tcK/Xe3TvqjP+/bFPF2MwC1xcCFiH/5Th4bQpQgAIUoIC2BJgSSluS7IcCFKAABShAAQpQgAIUoAAFcqQA6hEsd97ndk2oRfBXy7rVrwv/eP7s2dNcuXPnxhv0e7duWB0TEab1nQvm1Wva6huZVs0qCt6g1zUwNo0KDwnMal/aPh87FdDnxeCA8/gbgR+4IpChzrVq1m3YFDsyPNyPuMbHRkX8lC9ffpyX9uLZM3XOz0ybosVLlqrdoGnLPc7rV0l3UDRt07HbuJkLlo8f3KtzTky9pWiuOXXnTWbuC8+hAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKPBNCIgL4Uj3E5h0/1UlfUPjHUe9A0OuPfqnZYduf2sboXXnv/qEJj/+1zM86W5W+65YWd8AfXXuNWBYZvoqVKRY8T8KFS6SmXNVnbPMac9hjA3XQFsEH/A7djCoOhfHtx3x9Mc90NGtYojf23Xr1R/nW1rb1lXn/My0GTBq4rSAxHsvf/n1t9/F85EWDM+FNp+F7HQXx33AIyDqoHdIXGYc/utzsDPnz3IVdP7rcfD6FKAABShAAQpQgAIUoAAFKEABClCAAhSgAAU+u8DPwgq1f8KdFyi2jIsXK1Gq9KngSzeDrzx4I6Yi0tageg+1m4iFdyeXEz5Z7ROL6ejL0MyiuqZ9fSf8HPYJix88ZvJMTc9V1R59e0deS3Xzi0gU26KmBYznrXTaqep87K7AvBascf6QlgmBjvS5CjUtVJ2fmePfCz/HzkddWbR++wHx/P4jJ9gHJaW+bta2U/fM9KnonOx0F6+HBf/gqw/fzlm+cbu2xv05+5m2cOXGTQfcz37Oa/JaFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAVyhAAWqxs0b9MhT568ecUBoWjxxDmLV+XLn7+ANgeJBesKlfSqSK+V2f4nzV2yGgvqeX/48UdN+zAyt6yBAEC9Ji3banquqvbYFYG+Zztu2CZtu8X11DkESVSdj90VWHAvr6OrL7btM2zMJPSJXSWqzs/M8Wo2deqj/zqNmrcuWKhI0WVOuw/5xtx4ZFW7fuPM9KfsnOx0F6+JAFZWdt5oc76a9oU0bXAfP3Phck3PZXsKUIACFPi6BVjD4uu+v5wdBShAAQpQgAIUoAAFKEABCrwXQL2CU26u+16/fvVKRImLuhg2b7LdENS00CYUikhfvhQTJb1WZvuvYmxuIXR1USwWrkk/1W3qNkD7kAC/LO/0kF/XvLq1LT4LC7pwTnrsYkjAeexYETIu/aFsrNZ1GjRB+ij3Q/t3JcbHRovtfvjhh/SgzAvhhmgyT3XbtmjX5a9HDx+kIqB0wDMw2laoZXH/7p2U0mXKV9BGcEkcR3a6i9fQrWJsin9Hhgb5qzv/nNLOQNhBk7/Az79kx3OZU+bIcVCAAhSgQOYEGLDInBvPogAFKEABClCAAhSgAAUoQAEKKBTAwrcm6Zsy2jmBN9Er6RsYR4UFBWSGu2JlPYObQpXxB/fvZbmWhvz6ppZWNvgsPPDjgEX4+wLcVYzNLJSNGXUk3r5582btkrnTpW1+EPIc4fe0Fy+eZ2a+GZ0D59rCzorTRw/uR7AkKT4uxtfj5LGHqffvTZi9aKXzoTPnf/ujYKGM+sBx7J4oVrLUnxm1y0538bq6Bkamr169fBkXFRGmiZW6c9CkT3lbBIRQfF1ZH+IOmkg1nmsENjI7FqQoy+y5PI8CFKAABShAAQpQgAIUoAAFKEABClCAAhSgQI4Q+D5XrlzjZy1aUat+4+bSASG1EuofdOk9cLiygfboN3Q0UvUg3ZSyNljM7Tts7OTTIfG30HbXcZ8QRYvlqOWA49Ji0EhlNHD0xOmoAWBTr1Ez6TWwUDx2+vxlq7a5HF+6addBr4tX7p0JvZyyaN22/fjjsHrz7l6DR43XBjLqf5yNSn6Aa0r7K1y0eAmMGQXOFV0Huytw3H7Big3y4wgc4JgmKbpwjxw37z2ywnn/UbF4t6Lr2jZo0gJ9K0r/hD6Qnmrxhh0uymx6DRk9Aam50Af+4DlAHQm015b77wULFUaNlU37j3sPsps0I6P7hKLxSKuFNgULFy2G1GGomTJ0nP0cZbtFMpqDsms1bdOx29bDHhd8Y24+Rv0PfC9Qf0RRe+yqwX09F3vrif/lu2l4xsV2rTv16L1qu6s7CrW7egXHoti6+Fyijgnuvfy+oyg3+sEzg37wvfxrwPAxW4XgEuaKHTLycaAN5nkyKO4G7umSjTtd5R4WVrXqTJ63bG1GvhiL/NnWxveGfVCAAhSgQMYCSqPdhKMABShAAQpQgAIUoAAFKEABCnyrAggUdP67/9BiJUqWPnva3Q0OHf/qNxj1LvBvBC7u3Um5hRRTcqM7Kbdv4rNSf5Ytj5RT8uPYNbFs857D1W3qNPBwP+L66EHq/bZd/+73V/9hdssdpk+Utq8i7ATA7xHv0/6YWFS3Xrpx10EEN5B2qqVQkHtA5xb1gs77eKEdFtD1jEzMnz99+gSLrb/+/kdBYYNFYvFSf5bJI6za4px7KSm3snpfS5UpV6FQkWLFsUMBfUr7u5ty6+btG9eviWOXX2uQ3eQZ2Bmwftn8TwqBCxmh0lNCqbPDAm/PT563dE3rzn/1Ea+BVFLjBvXsqGh+WNx+9vTJ48BzZz3kx3GPj7ns2d68fZe/EGiS3zc9Q2OzYeOnzY2NvBjqecLtYN3GzdvgGYi+GBrktHLxPG24495iAR/BB4zPrJp1rROHXfZIU2aJ48aiPHZxuOzaurFsxUq6G/a4eeBeI7WZqUWNmsImn7xLZ08ZK52nqjnITXCNWUvXOSNggfu8Qng2K1TWrYLvhRBvy4PPpOcUEb4sG/cd88JzcWT/Dmc9AxOzQUKx96Ouu7ffup58FTtTcN7zp0+eIKj1WEjNVaxk6T/xXH4n1JfJl7/AJ3VkEIDC9wXPGIwRmLK0tq2LZ7pI0WIlOvToM9D71LHD4jjwTCxav21/rfpNWuC7+e///v23UYt2nRq2bNvp6IHdH2qt/D1o5Dj5cyudi66BsSnmMnFo764+Z04czer3hedTgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFMi0QPd+Q0bhLfoeQhABnSC9Ed6ux9vaTVp36Iq3w+cs37hd0QWwkI1zsZCs6PiMJWs24/zGrdp3EY9jcdQ/4c4LeXqoeSuddvpEX3+I4AMWb/Hm+m5331AUqq6kb2iM68xfvWWPoutg4RrH5btEMo0iORE7PtA33mRX1J/DKqdd2NkhPybaYBeIovPmrti0IzDp/ocaI8rGioVpvKmPMazbdfi0jp6B05xc/wAAHZBJREFUEd789whLvDNk3NTZis7DG/cYl7I+sVsF/Q2fMH2evM24GQsccQwL7Tj2U758+eGuyDYz7liEP38p5RnuLwICCHbhecNzgbnJx1NOiFZgPO269eqP3QoHvUPicA7GBYML8SnPEXCQnqfJHHAe2uM5RaBO7KdqDZvauK702cUx3A/s9sAuDCz24zOxKHvdxi3aSMeB3UV41kdPnbNI1bOI5yQg8d5LIZbxMwqkB1958KZb38Ej8X3AXMUUYmI/Y6Y5LMX42nTp2RefoR12GWEuYhuM1S/u9lNlu6SE2Mn3e0+dv4jdGcVKlCqtaow8TgEKUIACFKAABShAAQpQgAIUoAAFKEABClAgWwVmO27YhoVP7CTAwi+CBDuP+QSLqWWOno9MWi+81a5oEEjJ4xtz45GidDLigr18URxvn4vBEWmfbn4RiWt2HjqJt8sPnQ295OoZFPOLkHdHbINFbqTrUTSOrn0GjcAcxDf2tQk2bdGqTegbuwIU9YvFYBwvWbpMOfE4FoIPeAREYVH+j0KFiyg6DymZcFzVWKc4OK5D/0jrg37RHoEKfIbFZvn5WPTHMbxtr6xvjAltkLZI3gbBEQQQVI0LxzV1R2ALz4tneNJdMY0YAldYnMd48MzIr1u/Wev2OLZw7dZ93pHXUksI0QqxzcqtB47hGHY6SM/TZA4IoCBYIQ/+4NnGuISyEr9K++491G4irtmgeZsO4udiOjOk4pK2FQNtjVq276zKc/8Z/8gNe496durZf4g8yCc/17hqNSu0EXdBiccRvBltP3ex+Du+axgr6pgouj52lOA4HFWNj8cpQAEKUED7Aiy6rX1T9kgBClCAAhSgAAUoQAEKUIACX7gAChpfTUy4dP1q0uW2wtvaKBI8bfTAv1+/fpX+9j9S2yibIgpuR4YGBchTziC1zZjpDstSbt24vt5x/izp+ReFQtXb1q/4sKiKY1hAx4J/RGig/9Bx0+YIL/eXsuvfvd3jRw8fiOcinY6Q5eiRorEYmFS1RCqe+3dTbmv7dphUrW796mVaWlRYSKCivjEffC4tPt6sXece2Bmy02m1Y+q9u3cUnYeUUOg3o/HijX/sLECKn7mTRg36R/jBW/tNWnfsivP8vE5/EnCwsq3X6J+3b9/6eZ8+oaxvsTC58OL+J6mJkL4I1xB3WGQ0Pk3chXX/35Zt2n0IewEGdm3VQExF1VTYxYNAGQqT+/t6nZFfDzss8Jltw6YtZ08YMQCF1cU2T58+fox/P33y6KPnQt05YOcCAlIJcdGR65d+nLbLqnaDxjGR4SHSZw51K3oPsZt4zvPUcWmKtMrvd1rEx0RFSMcvBgoiQgIUBtrEtkh7VqGSXhWkxBo2YdrcLWuWLXA/tF/pDpmRk2YtwD10nGv/oUYLgkHYhREfE/khiGVsXs0Kz8KlmKhPAlsw7zdi/FSM4cCOzeu1/b1hfxSgAAUooFqAAQvVRmxBAQpQgAIUoAAFKEABClCAAt+QAN5uL1ehkm6g31lPBBn6DBszefeW9SvjY98tvGKXRSGhzgBqT8hZsOCJBeuLIe8W7KU/qLWAFDOrFs6aok6NBryhjvNRjwJpglYtmDVFWs8AfWER/VpSQryi22NWzapWeLC/n7ZvHRaSy1bQqYy6GmIAR36NuKiIMAQehMXhGjiGRePBY6bMQrDFeY3jQmVjErh/fJlBwAJvx4+bMd8R154+ZkgfMSiENF3ibo4ABQv81Wzq1I8KDwkUYjsPlV0bfb15gxm9fClv4+/reRqfyYucZ9UdacXKlK9YacqIfj3EYAWeIexYQN+okaEoIFVe513AItDPx1NeR6VAgV9+wRzkz5i6c0A9FezYmDV+eH/p/UWxdwTyQgPO+0rn3a577wFI2bR60Wx78XPcb9RkCfE/d1YaTMFx1Oa4d+f2LfnncksxsIF6FPfv3klZu3juNGX3Ds8Fdvs4r3VciDoeYjsUfkfdEq8TR4Wg0LsfY6EtgpGKAmPN2nbqjmcb5qxdoe3/OdgfBShAAfUEGLBQz4mtKEABClCAAhSgAAUoQAEKUOAbEUAxYywaI+jQsmO3v/MX+Pnn9cscPhSIFtNEJV9JTJCTYCdGvvz5C4QFfRooQNABQY4Thw7sVofSQAhYYBEdxaIvC6+D73Ba8yEPP87X0auSXtvgUnRkuLw/LDgXLV6ylHxxWZ3rqmqDN9TRBovRytpi4V94ET8QaXrQBjVBEGDBgrKyHSFo926HxUuFOywQnEEqqLS0tBeThGLIuAbOwb3q//6teHiJBcrFsSHAhLoSF3w8TmU0N/SP+gaKxnfm+GEXBDvaC4vzGfWhiXvDFm07IgCyd+uG1V4n/39BHYvmpcuWr4jrXAwJVLgLoVzFSukBi7VL5k6XjwcBpRtXryTKP1dnDkhjlp5+KcDPJ0J2bas69RvjeFjgxwEL1DNBWwRXcE2kLxOLhztMGTNUPg4zSysbdZ5LpI7CuXhuVsyfMUlRIEnsG2NAAMJ1l/NG8bMBoyZOQ3qnhdPGj5QGqvSNzKqKwUfp2HDvB46elO554azHKfH5UvV94HEKUIACFNCuAAMW2vVkbxSgAAUoQAEKUIACFKAABSjwhQuIdQRiLoYFd+s7ZBRS0UjTMFWorFcFU0xMiIuRTxVvemPRXEyJJB7Hbolywlvxh/ft2JLRwqu0P0OTdwELLPrPnzp2GNLYSI+LxZgvRUd8ErAQa0uECgvP2r4deEMdfYb4Z9w3FrEr6xuaIMDTa/DoCUgDtctpzfKMxpPRDosuvQYMQyHnhdPGjRAyIH1YkG/XtVd/LPBjR8GN5KtJ8l0UeFMfi+gXznpmGLAQa4Pg7X/5GNH37i3rVuoZmphjt4ayOajrjqCWnf3cJVcux8ctnjk5vbA7frC7Z9DoyTPE3RExkWEh8mshaFCmvE6lpPi4GHlQAW3/LFdB51Ls/6dAEs9XZw416zZsCsudG1d/UhTduk6DJuhLGowrXqp0GewQOeqyJ70APWpf7DnhF2ZhZVPHrl/XtvLAQJFiJUriHAREVD2XuNdoA6Mzxw4dyKh9Ddt6Dc+ednfDvcf4V21zOT5w9MTpqxfOnnpo7/bN4rlwL1ay1J/CVzdS3l+rTt17ibVAsmNnkqr58jgFKEABCrwTYMCCTwIFKEABClCAAhSgAAUoQAEKUEAiUEko0Ix8OlhoR37+3ZvXrpACoQ4Dfle0s8HI1KI6dkPI39Kv07hFG5xz8ojLXnWwsShdxcTcAgWlTx89uF/RAq+Q3t8I9RtQa0Dep6GZZXWMQdExda6fURsEUFBbQdWiLhbTsfthycadrkgZ5LRq8bwXz58/y6hv7LBATiZ5GxQOHygs5MdEhIcg6CMeR/HnQXaTZqBGwc3rV68kvE/bJT3fvHpNW6QJCleQpkvaDvcbvyNdkKIxblu3YjHSC/UePGqCsjmo695/5AR7LN4vmzN1nDQ1UY/+Q0djQd/71NHDuEZCbPRH9R/wWdESJUsjAON/zvuT2haYA+piKHo2ca6qOTRu1aHLw9T79zwlOz5wHnYf1KhVryECQtKaKEjvhOMvBOBNB9zPrtt95Ay+O92a1ba4IGSr+vS5tKiOz8KDLpxT9RwKgUEDtNkjBIrk9WCk52IHBgINuG+zlq5zPugVHKtvZFp1dN+ubTYsXzBb2hbfXXy3ribGx0k/x/yQhgs1a/C5sp0tqsbM4xSgAAUokHUBBiyybsgeKEABClCAAhSgAAUoQAEKUOArEqikb2AsrGdGI4XTtg0rl0hz4mOaQnmLKsjtjzfc5dPGYn5Y4KeLsdVq1q6Ht7/FtDmquMoKF8FiPAIDSIejqH0lPUPja0mX4xXVwzASCn9jl0dGC72qxqDoONImIaUOCi+rCj6Evy+8jTfl79y+eWPfNqe1qq6Z98cffxQyPaWnepL+9Bw4fAyCHo7z7MdL5zTIbvKM3wsWKrxGqG8AM0X3xKy6dS2k94JlRtcX3+hH/Q1F7XD/9jpvWG0p3Etxd4u8nTruGC+erVAhtZL3qWPpgQn8YOEdxavxuVCX/Rrmid0F8mv8Wa6iDj5TNFcLq1p1cEwo+u6v6RywkG9du37js2fc3eS7eayFdFDYgRIuS3WG4uu4zowlazYjADNt9KBenZvYmCFop+j68MFzI8TYPtkVJG2PAIKQ9koX37PjB/ftzOi+Gb8fg1BrZlLtRs1abVq5aG5za6MKnifcDsrPK1m6bDl8hu+N9Fjrzj16/ybcmHNep9xxzVghMKbqWeVxClCAAhTIHgEGLLLHlb1SgAIUoAAFKEABClCAAhSgwBcqUFFYYBfWS/PqGZma73Vev0o+DaSEuhwXEyUvOI3aAUjHEyZ7exyLrwiCIIUSdkSow2Jgam6Jdkdd92xXVCsDxcCRiidWCBzI+0NaIVwvMiwoQJ1radIGi/p4u1+dVFNIrXT75vVk9L9x+aI5ioocfzJ2YWKv39emEI8hjU+7br0HIADj7/Ou+DV+8HZ/ZyFNFHatpApVmbEbBTsApH1ih4eRmWUNRUEk+bVRWwHBH0VplsS2O53WLsdifutOPXpn1r3jX/0Goyj1hmXzZ4l9IFgwfdEqpzx58+RF+i9dA2NT7GTAbgX5dcS0RYpSV6EmBs5RVENF1Rzw7P76+x8Fg4U4ivyaDVu065ReHyQk4KOaGqiTgh0ZY/p3b9fKxkQHu1/kwQ5pX4ZCwCImIjQ4ozZoX76Srj6+N/4+XqeFOu2pGT2jRYuXKIXjS2ZNHtPIonKp1Yvm2GMnjKJzihQrXhKf37qRfE08ju9LvxHjpmInFYJG6QXjFRRe1+R7wrYUoAAFKJB5AQYsMm/HMylAAQpQgAIUoAAFKEABClDgKxPAW+J4kxwL8/u3bVr77OnTJ9IpYhFVWaAAb4+jbbhsh0WJ0n+WxXk3ZYvpGdGh5gWOYwyK2lWorFsFi/ExEZ/WOCgv1MrA9aKFGhzavj2oB4E+gy8oL7gtvaYQKPDF2+wHd2/dpM5YUCBbvhOibpOWbRG02L/DaZ3YB9IezVy6dkvKzRvJsyeMGCDujhCMr0ivg/Re2JkhDyLJx4IAEN7ORyqmjBarESRAqqNa9Rs3l/ehrnvz9l3+QmBFmjIJgRfUxnCcaz8+LupimJC5yPBm8rWP5iJeT4gpFMK/ESiQjgEBM9Sg8PU4eSyj4JCyOSBQh/7iZfUvsIivZ2BshqCKPFWSkDGtIOqJoKC3OsE43Cd1nkvdKkamGIuH+xFXVc8NxoA2e7duXC3fDSU/94/CRYri+Xr0IPW+eAwF4fMX+PnnretXLK6sb2SiKECoagw8TgEKUIAC2hNgwEJ7luyJAhSgAAUoQAEKUIACFKAABb5wgYrCQjGm8EZ4y3/X5nUf1a7A53gLHcEARbUhjM2rWd2/dydFWhAa5yAFEP6+q6CYszIuA5OqllhYjgwLVrhLQkfXwAjnonaDvA9h4Ty9xkZifGy0tm9HFWMzC7xpHyakLVKnb4epY4b1bF3fSr4bRdm5SDklbGD4KHWTTd1GzbAY7n3yXfokBGrmr3HeI7wsX3rC0F5dkKoJ9wXHhMxT6Ts6xB9Tyxo2eJtfvjNAfv2mbTt1Fxatf9m9Zf1KVfPCbg3UisAuCWlbddzLVaysJ5RbKO914ughMbUV0jjZTZ272OfMiaM7hGLXCM6gZoe4O0U+HmFDQPp1X7x49lE9kPbCLhQEfKQ1PpTNRdEchNIYZdA+5dbN69Lzhk2YPu+m8FAjCCKvjfGLEC1QdzcCgoFIc6bOc4kdJhiDn9dpd1X3A2NAm9dq7IqArZCR6qnYZyFhywXScG1cvjB9BxAKcqcI+bhUXZPHKUABClAg+wQYsMg+W/ZMAQpQgAIUoAAFKEABClCAAl+YQMXK+umFfj3d3Q4qSrmDdFA4nnjp02AA0t0gbZF8yngzHZ/9JKRSkh8rW0GnMhanpZ/jbX8doaA20uEoq0Eh1lBIiIv5pOB2iVJlyqI/aXFkLAD/lC9f/qzeDgQsUJ9AVZoe8Tp4k12+EyCjMeQSIhbyGhb6xmZVsUtDiEs8gOXEWYtW1qhVt+HiWZPsRG8hNVFp9Csvdm5qUaPmJSGog1RHYlFt+fWxkD566pxFXkKhaXnqKNwb7KiRnvOdkHoKARR5WiN13PWNTauir4j3NSYqCJXTF67btl9IUXR16sj+f+FYUaHqtqK5iGMQ5ygNmKA4fI8Bw+yuJFyKxQ4L6XjVnUM+YZcBzpP6G5lb1kB6MRTVxs4IBPLQBkEj/C2s/T8R4icfBW6U3V/sNJI/l0hvhbRS8nMqVzE0wT1XJ3iAMeB8MZCT0fOF9E/SNFsTZi9amSoEGREoEutbqHPNrH6PeD4FKEABCigXYMCCTwcFKEABClCAAhSgAAUoQAEKUOC9gBiQcN3lvFERCgpu43Nh88MN6XG82W5oalFNXIiWHku+knQZv6PmgvRz/L7b3Te0VafuvaSfY4EYuziCzvt4KbsxaIOF17vC6/DyNtilgM9+ylegAP5uJuwe2HnsbLB59Zq2WbnRWOwtL+QqCvFXLx1UZq6FgISwweKjHRZIgYSgB45NcXBc175Hn4FIlbVLqCchXkOI8fyAfz9/9uSjFF7CDouaUeEhgev3HPVYsWWfG4JB0nFhMX+Z0+5DwqL309njRwyQj3nS3CWrt7ieOvdHocJFcAxv5Lft2rNfeLC/n3zXiDruH9I5Pbh/r3IVI5ON+455YV7D/u7QXAwCiXN59n4hXj6mq4kJl/CZmMIJtTumLVq1CanMls2dOk6emkndOTx6mJpeK6JE6XcBr8JCcQiHlZt3LZ09ZSwCF5gzAj8Y84I1znvRBmPB7hapK8aDZw5jko4dwSjpc4n0ULvcfUO69B44XD5HzA21LtR5huQe4jkIVs1aus4ZuybEz9KE7RXiv1H4vJ6QbmzxzEl2uJdIM4Zjd2Q7TNQZA9tQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFNC6wNbDHhcOnQ29JO6KkF9g4dqt+0KTH/9bsFCRotJj2CmBz4dPnOGw85hPsLzGwartru44jje6rWzrNeozbMykC/Epz0+HJtzGIri0LxRlRlssaCuboEdY4h2vi1c+qmEgtm3cqn0XnD9vpdPOMdMclgZfefBmubBYr2xO6iLqG5lWRb+NWrbvrO45mrbzi7v9dPGGHS7S81w9g2KCklJfH/ENT8D1l2zc6Sq+4S+26zVk9AQcW+G8/6i4eI639/FZ++69B6AP/HvtzkOnmrTu0BV/xs1Y4Ogbc+PRkXMXL5etWElX0VhbdOjaE+e5eARG47pno5IfnL+U8gy7aeTt1XFvJBSvRn/Hzkddwf1HX1hYl/aFoubekddSfaKvP1RUKwPBMc/wpLsnAmOvY9F99Y6DJ9CnPEAg9qnuHBBACLn26J9NB9zPdu0zaMTxC9FXYYQaFugfzyy+G7gP4rNp26BJCxybvWz9VjzXCD7AStF4EABB//iO9R85wR7PMBzElGnieBFgwPmo66HO84MgSkDivZc7jnoHouh4s3ade6zZeegk+thz4lwYapiI/WB8+HzR+u0HMJaZS9ZuEY8hgIhjljVr11PnumxDAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUCBbBbDoadugaUtlF9nsctL3ZFDcR7sr0Ba5+f0v303DgieCE+Lb2mI/SCuEBWYcF/9sPXTmvFh7QXq98TMXLsdiKhZ4FY0DgQcsWLt6BccqOo7dGdgVgOugH4dVTruwCJ5VOCwEBybdfyUPsGS1X+n5Z0Ivp2C80s/qNm7RBp9jgRsBIcxPfk3Mb9U2l+P+CXdeiLshxAACAi1w3nXcJ0TqL/Ynv1fSvmEt3g/Mfd2uw6fFAt/yMajjjl0qGCcCFc4HT/uJxdXlfdVu2KwVgil29vOWKPJFwAVBHPEe2y9YsUHc4SFvr8kc+g0fNwXPTHoQwnHDNgSGMBb8jsCXw+rNu1HrQ7wG+sYOFanrdjevgHpNW7VTNG6k3hLbIrCnKE0Xgg6Ym3RnhKpnrEf/YXbSMRz3j77Wc+CIsfIdNfhOeUVcvY+2CIxJ02qVLlu+YnowQ0jRpep6PE4BClCAAhSgAAUoQAEKUIACFKAABShAAQpQ4D8XwNvcinLuY2CoKyHWwFA0UNSQwOIvFv71DI3NlE0GNRWQeimjyQr1kcspC2iI52HhXvp2eVbxUCfBuGo1q6z2k9H52G0A48xeQ7poj90BCDJIF61xf8wsrWwQQNJkxwkcUbBZnXFpyx3BgozGKJS6KIPFfWW1OeRjVXcOeK7EGilIM4UgTfDVh2+xU0XZ/PUMTcwxFiz6qzJCcO83Ic2XsnbYGYO+VPUjPw4H7EhBvRb5DhxpW1wbtUMU9Y/AT0bz1HRMbE8BClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIU+B92MCAlECkyJ2BgYm559HxkkpgSK3O98CwKUIACFKCAZgIsuq2ZF1tTgAIUoAAFKEABClCAAhSgAAUokMMF8IZ95SqGJjGR4SE5fKg5cnio9eDkcsInNOC8L4paR0eEqVUAO0dOhoOiAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABCvxXAkj9lF64WShK/V+N4Uu8LtJGobA86lV07zdkFNJpIa0WinB/ifPhmClAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIAC/6lAs7aduiNgYWRuWeM/HcgXdHEUJnf1DIpBQXcLq1p1MHTUpoCjiUV16y9oKhwqBShAAQp8wQK5v+Cxc+gUoAAFKEABClCAAhSgAAUoQAEKUOATgUr6hsb/vH37VshlFE4e1QLlKlbW27DXzePFixfPe7SsW/361aTLOAtF1uEYGxkeqroXtqAABShAAQpkXYABi6wbsgcKUIACFKAABShAAQpQgAIUoAAFcpCAjp6B0ZXE+Lg0YQE+Bw0rRw7lp3z58jtu3nP4f999993Azi3q30i+miQO1MzSyuZSTORFOubIW8dBUYACFPgqBVh0+6u8rZwUBShAAQpQgAIUoAAFKEABClDg2xXQ0dU3jIuKCPt2BdSfec+BI8aWLlu+4qxxw/tLgxUoXF7Npk798GB/P/V7Y0sKUIACFKBA1gQYsMiaH8+mAAUoQAEKUIACFKAABShAAQpQIAcJ/PLrb78XKlKsONNBqXdTmrXr0uNKwqVY71PHDkvPqFq9pi0sz3ufOaFeT2xFAQpQgAIUyLoAAxZZN2QPFKAABShAAQpQgAIUoAAFKEABCuQQgYq6VQwxFKQyyiFDyrHDyJ07T56SpcuUi4+NipAPsk2Xnn1fPH/+7IKP1+kcOwEOjAIUoAAFvjoBBiy+ulvKCVGAAhSgAAUoQAEKUIACFKAABb5dAZ33AYv4mCgGLFQ8Bm/fvnnz6mVaGnZSSJvqGRqbNWzepuNRl93bXwoFLL7dp4kzpwAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpkUmCKg+M6z/Cku5k8/Zs7bdG6bfsDEu+9NKtmXevHn37KZ2Vbr9HJoLgbF+JTnpcqU67CNwfCCVOAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFtCGw3c0rYP0eNw9t9PUt9FG0eMlSbn4RiaHJj/8V/wRfffi2ZYduf38L8+ccKUABClAgZwnkzlnD4WgoQAEKUIACFKAABShAAQpQgAIUoEDmBL7PlSuXjq6+octO5w2Z6+HbOyvl1o3rnRtZm6JmhZ6hidmjB6n3D+/bviUmIjzk29PgjClAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACWhD4vWChwtgtUEnf0FgL3bELClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQAEKUIACFKAABShAAQpQgAIUoAAFKEABClCAAhSgAAUoQIFvTeD/AMRAp16fSAweAAAAAElFTkSuQmCC"},{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO3deXhcZ33o8e97zuz7aDTaV8tabEne5C12bCdO0pAVAoFcErZCA5fL0qe3D225lEKhpfTe2xZKe7ml6QOFtPQGkpIFkpA9xI7jfV+1SyNptMxo9n3O/UOOiBPHlmzJI1vv53nOY2vOOe95z2jmp/e8q9DpdIc0TWtEkiTpXQghOoWqqvFcLmcudGYkSVq4VFVNKIXOhCRJVwcZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhEZLCRJmhFdoTMgzY7FakOv16OhkUokSKVShc6StEjIYLGAGUxW1m/ZzobNW2lpW4HT6SCTThGLRlF0Omw2O4oi6O88yY4Xn+XZp35BPCGDhzQ/5FIAC5DN7eWjn/kDbrzpBva+9gKvv/ISx44cZDIQJK9p5xyr0xtZuqydm+78ADfcsIVvfekzHDh0rEA5l65VqqomUFU1DmhyWxhb24bt2v977nXtvzzwgGY06GZ1bnXjCu1nL+zSSjyOgt+H3K6tTVXVuKooylc0TdMjFVzd8rX8xV9/iz/61IfY8dpOcrn8rM4PB/wYi6pZUmYjmNLzvR//DGMuzLFjJ+Ypx9JioShKVtZZLCCf+/Jf8Hd/+gX6BoZmdZ5QVBxOJwLIZtJ4ior5zJfu58l/e4j7PvYgz/76pXeck04licfjc5RzaTGQwWKh0Dtprrbz+p7Dsz61pLqRP/nanyPE1M+KzsDKlSuw67OU1i/n63/7/Xecc+bAa/zj33/vcnMtLSayzmJhbMLg0p58Zacm5iAtT12b9oMf/lADvfb4yzsLfm9yu/o3VVXjslPWAqGlJznSOc773nv7ZadVUlKB3z+EuaicWMA/B7mTJJAVnAvIvl2/4b999X/Rvnwpw4P9BIPBS0qntnUVtUVm/FGNKq+FF59/cY5zKi02soJzgZkcHeSzH3wPN939Ib7wZ39DWWkx/T1nGOjpZtQ/zMTYOBNjfiYDY4yNjhIJh8+bjkGvks3kWdmxnoO7dwGgM1r54pe/xsPf+0tGJ0JX8raka4QMFgtMLpvm1489zK8fexiD0UxNQyM1dUsoLa9g6fJ21hfdiKekFHeRB6vVymDPaX716L/x/K+fm04jm82jqgqbtm7l25/7LgC33/8Z1m+6noEjW/jZo0+d58qCxtYVjA/1Egz+NphYbXZi0cj5MysULBYz8VjsvLtNVhd33nMPv/zZwyRSmQvet9FkwWa3MjE2duE3SCocWcF59W6KqtMa2zu0v/3xk9qnP/3J6deb192sPfTIk9o///gn06998NNf0p7de0b71c5D2hO/2a+1L1t6Tlqf+crfat//8SPaI8++ojksBg3QbMVV2s+fe1XTCTRHeYP2jW9/65xzbrnvM9off/mPNUC78+Nf1G7Zvumc/X/6vZ9q//bUq9qdd9ysIRTt81//jvbLnYe0NSuXn3PcB37vv2uPvrBL+8EjT2v/+NBDc1LJK7e53WQF51Uun8ty5sg+/vxP/oCb737/9OtDfV0sX7ORx37y0PRrP/vB/2Lf4RN8/XMf5tEnnqGhccn0PqO9hNtuWsfnP/4hBoMpyoqdAPzOPffzyhP/TlaD0vJqbGbrW64uuPfDH+Gxf/9XAOqXNCFQp/dWLVtHU4mOp556DqPZxG0f/ixV9izf/ft/ZOPGzdPHbbr9fm7evJKP3L6Fzz7wPr79zW+ind134613zOG7JV0uGSyuAR5vGeHAxPTPkdE+znR2c+jgwenXmtfeSLUjx/7DJ6ioqGLY55ve9/6P/1eio8O0bXoPxbo4XYNjqAYL93304+zbtQOA4tJyIvHJ6XOa1t5AnUels29kan/Zufvvuf8TPPnIT7AXuxCKjU98/D6+/fWvYjbZiCSiwNl6lD/6Mg995y9JpDLc9bEv8J5btgLQsu4mHvjIffPwbkmXSgaLhUjR8b77P4GnyHXRQyvqW/jTb/4lP/z+WztY5Xniscf4yCcfBMBodfHHX/sm3/nmV8jmNKxWK8lYAoD6tvW89/Ybsdet5AtfeJAvf/5Bcnn4+O//GeUeB1ouDwhuvv1uqqsbptKzOPijr/452fRUPYTNU86GDeuoObt/+brtrGut5vHHn8LjKeXO+z/Jf/7L3zEZSaDTG9G0HACf/MM/p7qsiHg0gs5o4e73f5B8NoeiM/Lfv/JnfP9//9UcvaHSXJCjThcioXDvJ7/IBz50HxPDvRzat4e+nm7Gx0bRNA2z1UFVbT2rN26hotTN97/9NXa9seecJHRGK3/zo58TGjxFdfNqXvnPf+FHP/wxALfd/znuvmUjO3bt5+57P8g3fv8T1Ky+hffftZ1fPv44reu2UWrL87PHn+fBBz/BwEiQfGgAR+1qxroPsaRtHb/68Xdp3vZBzJkA1c0rePaxn3LvR36X115+iY716/jKZz9CT/8Q3/7hk7TWOrj3d24klc3T1LGNb3zjq3T2jmAhzNMv7uZTv/dx0jkVTcvywr//ExlPM41e+MbXvlGAN186H1VVEzJYLGBCKNQ2LqNt5Wpq6huw2WwIAZlUksHeLo7s383JEyfQ3jZs/U2q3siaDZuJjPs4efLUW1Pm+t+5m8oyDy8/8wT+0XEAlndsZtWqlYz0d/LKC8+Ry2ssXb4Kp83I/j1vYDQ76Nh4Hb7uk/T29qHqjXRcdz3+vtP09Q1QWddEfX0NB3fvIHq25FLd0ILIROnvH5y+elN7Bw6Lnv273yCvaZRUVJNPJ7j53gdprq9k+YoWfu8DdxCJy7k5Fgo5RF1uC2q7/7N/qr12tFtrX95Y8LzI7dxNtoZIC4aiM7Jx2zYe/odvc+T4mUJnRzoPGSykBeHeB/+QtuZ6ghMTFz9YKggZLKSCs3kq+dAH7uCnDz+MIuRHcqGSvxmp4N730U/z9E//iXAsiUAUOjvSu5DBQiosoeOOO+/g8Z//HJ1qIJO/8BgSqXBksJAKqrqlg8jAEcZDcUwOB/G39AKVFhYZLKSCWrZyDYf37wagtLSMsWE5Wc9CJYOFVFDeMi+jvgFA0NjUQFdnd6GzJL0LGSykgpoMTFJaWc2qrXeS9p9gIpIsdJakdyG7e0sFZXWV8K1/eAiLmuVbf/wFevp9Fz9JuuLk2BBJkmZEVdWEfAyRJGlGZLCQJGlGZLCQJGlGZLCQJGlGZLCQJGlGZLCQJGlGZLCQJGlGFE3TZMCQJOmCNE1TFU3T5AQCkiRdkKZpcloiSZJmRgYLSZJmRAYLSZJmRAYLSZJmRAYLaVESQtbrz5YMFu+ivrGZTTfcTGNLa6GzMudUnY41GzbPWXor1qybs7Tmk6rT8cGPfort77mL67ffittT/I5j7A4nLW0rC5C7hU9X6AwsVHUNTbz0zJNUVNfO63UURSWfz83rNd5u3XVbyOXzc5KWEILi0rI5SWu2VFUll5v5e1dU7OXAntfpPHn8XY+pW9rE8ODAXGTvmrMoShaKouByF83qnFw2i8FoZGigb55yNaV2SQMABqNxXq/zJiEELe2rGPFNfSEsVutlpef2FDMZCEz/vPnGWzBbrHRsnLuSy1sZjEaEEAghcBd7Z3Xu0qZlDPReeI5Pb0kZgfHRGaXnnOVn6mq3KIKF3mDA7nTN6pyDe3exsmPD9M/lVTUAmMwWDEYjJrMFRVEwGE04XG4ADAYjZRVVM76GEAKnuwghBCVlFbPK36VqX7OOU0cPExgfw+5wcte99+Mq8mCx2tDpdFRU12Kx2nCevSeX++w+vZ6mZW3A1F/osooqdDo9dQ2N9HSewmqzA/D6Ky9gtdnY/8ZOrDY7FpsNh8uNyWSek3u0O1wgBEaTGYdjdr9Tb2k5K9asp2PjZoRQ0On0VNXWs2LNehRVpWPj9bg9xeTzeZavWI2nuOSC6bmL3vkYcy1bFI8her0Bj7cEg8GI0WQiHJoklUySSafJ5rIAZ39OYXc4EYpCeDKIxzv1Ydl6823k8zksVhtNy9rI5bIoikLnqRMsX7Gaqto6/u/f/BU33X43mqbxzOM/n1G+zBYL2WwWs8XCsvZV3H7PfdgdTuKxKPF4FJvNQSQcwj/sIxoOE5oMEo9HiYbDJOIxhFAoKi6e+uI4XSTicUAjFo0QCYem0onFpq9nMBqxWu2EJgMoioKiqmSzU/eyYcuNGI1G6hubObD7dZwuN0cP7qOhaRkWq5V4LMrE+BiqqnLfJz7Nob1vsKSxBYPRyPrN2zCZzDz+yMNs3LqdVWs38thP/5X2VR0oqsre119j07abyOfz/PrJxzAaTdTUNxCLRcnncqg6Hfl8Hp1Oh9lixWQ2Y7XasNjsJBNxVFUlnU6TTMQpLa/k9VdfxGZ38LH/+kUmAxOkUklURcVgNBGNhEinUgz7BvEP++jrPkNwYhyAYd8Ae3a+Ov1+1DcuZ8P1N/DIjx/i5tvuZu+u12huXcHSluVomkZTazu7Xn0Ru8OJoqroDQYMBiP5fB6b3UGxt4TertNz9Cld+BZFsNA0bTpQFBV7Ka2oJJNOExgfI5VMEgoFScbjAKzdtJWXnnkSgFg0itVmI5/L4RvoRVEUKqprePz/PUzbqg7KKqrwD/uIRSNU1dZjszs4cmAvAFabHVeRB7vDibe0DJ1Oj6vIg9FkQq83kMvlKK+spqfzFKlkks6Tx3j+l79AVVU0TQNA1emx2R04nC5sdgduj4cljc2YLBYUIQBBJBIiFAwQmBgnGg5PfVnSaVLJxDnP8zX1S7ntfR+kv6eL+sYmPN4SDu/fw8mjhwiMj+EtKePw/t2YLVZ6zpyiorqGZW0ref5Xj3PLnfdw8uhhKqqnSlfRcIijB/dRU7eE7bfdzT9/939y3babqK5bQjwWpbi0jFBwgqUtrfzgu3/NksYWLBYrRw7uAyCVStJ1+gRlldXUL23CbLVhs9tJJZJkshli0QiJRJx0Oo2m5VFUHYqi4PYUU1Vbj9VqY2LUzxu/eWk6MGuAePPfs48pRqNp+v71BgOZdPqcz0VL20qe/+Uv0PJ58pqG3eHk6IE9rOzYQGBinN+88AyaNhV8HS43DocLvcGAqqo4XG7KK6sRioI2R/U/C92iCRYmi4XdO1656LHGt9QdmM1myqtqGRrso7l1Ja8+//TZJjeN8TE/a9Zv4tF/+yFrN22huKSUF55+gsD4GACxaIRYNALAyaOHznut67bdxOjwEEazmUw6haZpZLPZ6f25XI5AKjnjZ+gL8XhLeOrRn+Lr78XucNK4rJWauiX0n32Gd7rdjI4MUVpeSeuqNbz2wq/ZuPVGKmvqGPMPMz7mp3XlGkrKKzlyYC/L2ldx/NB+Ok8eI51OkU4laWlbSTwWpevUcZKJBH3dZ8hls9TWN/D8rx4nHPrtamP5fJ6hgb5Z1wnp9QZGhgZRVRWnu2g6sMJUoICp37cGJOK/LVXVL22iv6frnLQS8RgjQ4O43B78Qz7u/uAD/Oj738Ht8bLj5efIZqaWUszlcgQnxqdLKDAVkG65855FEygAVCHEVwG10BmZT3qDntr6pfR0nrrosdlslrbVa6mpX4pvoJf+nm7Wb95G56njpJMJ+nu6sFitjPgGScTjDPb34HC6GPH1s3LtRjLp9Dlfigtpbl1B16nj5LLZ6Uej+dCx8XrGR0cY7OuZvkenq4hEIk776rX0dZ1Bp9OjAZ0nj2G2WPEN9FJVU0+Rx8vuHa+w7ZbbCU6MU1xSSmlFFWMjw0TDIUKTwak0MxkcThf+4SHC4UlCweB06S2TydC+ei3xWGw6gF6qomIvvoE+8vk8Y/6RGadXWl5Jc9sKauoaplu4QsHA1GNMOsWaDZsZGuyn6/QJLFYbjS3LL1gZqigKZouV0ZGhy7qfq4UQIo8QIsVUUL5mN51Op7mKPAXPx9s3RVEKnofZbptuuPnC96TqNEATiqKJebg/i9VW8Pfgt/eqFjwPV2oTQqQXRWtINptlMjBR6Gy8Q/4qLMIqyoU/Mqo6VUidr+J5PBadl3QvRX4WfTyuBYsiWEhzQ1GUiwbdTDo1/f/F9Dy/GAghRErTNEOhMyLNhTfbAyRpbgkhMrJkcQ1R1KurnloIgcFovuryvVjJYHENyeeyFz9oAXEXl7LxpvdS17xKjgK9CiyKfhbSwqOoKuu23UHHtrvw9Z7CP9BFLDKzJmepMGTJYpExmm0YjOaLHDX1V37e/9oLlXRqqtt97gqPvJVmT1ZwLiJ2t5eb7n4Ak8nIMz//EZMT/vMeJ4Q4p2fkfHEVl7Fk2RpGBroY6r14hzmpcIQQGfkYchFCQHMVbG5Xqaksgswk4ViGA2dg53FIpi+exhzmhstp7dCpKhs2baKssppRXw8vPvXIeY97t0Ch6gyYbXYUoRIJjV920+jk+Aj7f/M0sgXn6iCDxbuwm+HWtbBxObS3tVK56rN4qjeSSYYZ6NzFh3VJ/N2v8stnXuX5/XlOD85fXoRQaGxdjdPt4eSRvUQmAxc/6TwioQl8PScpLy9FYXaVoYqqo3nlJlZv/h1isTCvP/tz/IOdl5SPc8lAcbVYFGNDZkMA21bA1x8s5q47tlOz8uPUb/4GOkcL6Bx4K5pxlq3EXtpBRfMdXH/99ayvOkqRcYxjfZCehwYJs9XKvb/7+6y+/j0YzA76zhwhl83MOp18Po+vv4e+zlMc3vvGOQOtLkZvMNK24SZWbrwZh8vDcH8no74LTyRztRBCmR4gKJ2fECIvSxZvoQi4dxt85I4aqq77NmbPCsrLq1BVleHhYWBqBGImk8HhcBAKaUxqy2i69d+52/xlqrzP8Nf/oTEentt8pZIJzhw/iKOoHEWnx2A0k0q8+xfdYDCSzWbPO12fr78XX3/vrPOQSScZ7D7BYM8pctkMQ30Xr2MQioLLUwoaBMeHZ33N+aLqDFjtXix2D86iCiyOYoQmCE0MEJoYJBQcIpOOFzqbC46s4HyLj94CH3tvE7aW/4G9bC2aplFXV4eqqvh8PlKpFPF4nO7ubm655RbMZjPRaJRUKkU0HGBoz59xYt/jfPVHELy8wZXvYDCZqaxvIRGLMurredc+FWarjVXrt6JpGof2/IbEHI6l0BtMVNS3kIiGGfX1cLG/xDZHEfd++k8wma08+i9/zdhQ/5zl5VKoOgPe8gbW3NqIyeYhMlaPojOh6nSAIB2PMDncTXRyFF/vfiKTIwXN70IihMjIx5Cztq2A//H77yVf+UUa2rbj8XjQ6/Xo9Xq6urowGo1UVlaSy+Ww2Wxks1lcLhcGgwGTyYTRZMFdfSNq/Bjllm5eOwL5OSzV5rJZJif8REMBNO3dKxbtDie33/dplndcTzwcxNc3F/UKU/K5LKGJEWKR4IyOV1SVtdvuorhiCdFQgP7OozM6z2Ays2z1JlyeEiKTE7OalPfdmK1ulq29m6Z1W2i9eRJ3tZ/wmEo25SSbTaOqOvJinKKaCUwWByZ9FaGgj2xmfqYNuNoIIfIyWABuG3zr8w24Wr9Evz9Le3s7RqMRs9lMPp8nGAzidrux2Wzkcjk8Hg8mkwnD2VmTYrEYfX19VFXX4qq6AV3gUfxjEboKMNWBpml4SitwF5cx0H2SwZ5zp31TVBVPaQUWi5VkIj6vTaTZbIZEPI7BZKb7xH7Gh2dWsqhZ0sL7f/cPWNq2lnh4jGHf5ZVILDYP7dfdi7u8nrymZ+i0jqHTCjq1CfI6BAKDdYTi+iG0vInmrT4S0TykqgiOD6DJPiAyWLzpgZvg9nsexF79HtatW08qlcJgMCCEIBgMUlZWRiqVIhAIEIlEsNlsqKrK4OAgdrsdg8GAzWZDr9cjVBNjY0HqLTt5Zg9krvDnLJfN0nvmGKeP7KHr5OF3VISWVNZz9wOfY9nKdfgHu2c8Uc+lGh/uo/v4PkZ93TNuajUaDTQtX4XN4aD31GGG+i+9IlUIhdYNd1GxbCmlzZ3k8yPkUtUISiCvmy45ZJIQmUijaV0UVWk4yhLEAhqqVsXkeD+LvfJTBgvAaoI/+VgRlWu/QlVdK/39/ezcuZOWlhYA9Ho9+XyeaDSKwWAgm81isVgwm82kUimMZ6em1zSNdDqNxWIhoxQT7vkZ48EknQUoXeSyWaLhSXLZd9Zr6PQGWlZtxO4sZtTXi/8y/2pfnEYmnZxVn4x4NIqv9xRnju7l1NED09PbXQq7q4zr7qmhtqMXuzeEw2vD4oDImBtFUVH1BgxmjUTqV3jrxzA7U0QnbMQnVXLaBLm4l0Q0TjIxx7XWVxkZLIAP3wh33Xk71rr7MJstTE5OUlNTg8ViQQiBqqp0dnZSU1NDJpPBarUyMTE1p4PX652eebqnpwer1Tq1PIDJRjgSo878Or/eC5kFNL4rlYgx3N9FcGKUnlNHSCXmr9bfaLbiKiohmYjBrB53NMKhIBOjI+fMSXopapasZflNOXTmGGG/Bd/h9eRzJjJJM0IooGnEYwNk0kliY2sY6c5gtTeQTVqxuS2kU2Okwk4mJxb3wkOy6RS4eQ04StvR6Qwkk0mSySTWswvvvDk2oqGhgUAggMvlQgiByWSanhFKCIHZbKa5uRmYmilqZGSEtGkl2zpcOK2TxApQRyaEoL6pDU3T6Os8cU4zqn+wB/9gz7znYe22O1i2ejM7nn2EE/t3nPcYRZl6H+djVTad3oTd7SY6OYar3Etf11oyKQOZMR2app0tEebQ6c2ULnWTjkdIRVagsR9XVZCJwQTZXBa7sxGhqIu+7mLRDyRzWMHsbCQSiZDL5XA4HHi9XnQ6HYlEgnA4jBCC0dFR0uk0Op0OvV6Poijkcjk0TSMajRKJRKannDMYDKRzBiyuOsxXZqGxd/CWVfHeBz7DXR/+FBU1SwqSh1Q8ht5gpq5pBeI80/EZjCZuuPN+tt55PyaLbc6vbzI7MLsgFW5n+JSbdDKJ2TWCoh9BKHnQNITOT/XKYzSsH6VpcxclTa8wcMSOwWglG1tLKrwORdUjkEPoF33JQlUgl4kxHhnHZDJRVVU1NXP02BjJZJLS0lJCoRCJRGJ6qn7dWxbFebPiU6fTYbdPrcrldDop8hQjUhpKgT5jpVX12JzFGE1G9IbZdaMRQmC2WEmnUmQvoafomw7tep5kMk4oMHreOgujyUJNUzs2hxtfzynOHNl9ydc6n2w2RSKs4KoYIJsqRWcwkgiBTm8nlwOhAHknGlEiE3nsxSZKGwzUrhnnyPOVCEwUV1bj7zyItsgrOEGWLMjmIBrsorq6mlgsNl1Z6XQ6qampQVEUotEo9fX1mM1mwuEw2WwWIQS5XI7k2en7nU4nqqpy8uRJjEYjdpuVfGqcXIGmoezvOsnxg7s49MbLjPhmtzZHRU09n/jCV3jfRz6N2XLpa6Fm0imO7n6Jgc5j590fDU+y75Wn6D5xgODY3NcEJ+NhUrE0/fs3Mt5TTf3G18hoLxILRRFianEggY2+PRvwHVvCSGccvVGleRMggri89WTTSdKJiJxPFFmyIBiB6NgRrI2/fSv6+vo4duwYt912G8lkcroUARCLxab6Mng8+P1+XC4Xbrcbi8WCpmnYbDaEEGQiXYSCI1d4VOpvhQJjPPnTf0Kn6mbdi9NsseOtrKO8Zgn7X3+Z7lPn/7JfLk3Lc3TvbzhxcBfZzHy8URpjw6fx1iwnnQmgN2aoW5VncvgwwYFa9PpaEAKDyUts3InZOUJgKEYuK7A5rpuq/AyOEg4Os9ibTkEOJEMIaC0fIu24jboljeh0OqxWKxaLZbrnYFlZGXq9HoBAIIBer8dqtTI0NERJSck5q5i5XC7C4TD7n/4SR0708fjOqdJLIeSyWTKX8CUMTQaIx8KMjQxx/OCec2bsng/zUbn5pmwmhaekHouzlkx6kOXb7NStEAT9E6RCteSyGRRVh6rLUtY8gs6YIjyaZ9JXjJZTiYwOMtC9Z9H35JRNp0DPCNyyOkMqq1Lf+h7S6fR05WUwGJxuHs1ms0xOTlJWVobRaERVVdxuN36/n1AohMs1taJ3PB7njR3Pku/7Hj98RpuXXpyKokxFuXnqfanl8/h6O+k8cZhMeoZfEiFQVN0Fu6IXQi6Xxmi0YXOWYnHaKGkIMuFL0bO7BVVxkc0kyaaT5HOCTNyJrdgHuSJyuQgTvRmG+w4THOst9G0UnAwWQC4POhXayvvwND1APPHbjlZGoxGLxcLY2NhUPYTdTjgcnh4boijKdG9Pk8nEyMgIBw4cYOL494lMdPODXzLndRbFZdWs33ILJpOJSCh43o5Xl2uqOXNmQ7ZNZgtNy9vJpNMkE4kZnXOlxWMB7DYvBluY4toEr/3EidnSihAKOr0BRdEhFIVMwoSjZJzuN1xMDir0ndjLyODMxrNc62SwOKvXD9taE1TUthJKuXG5XAwPD2OxWLDZbCSTSTKZDCaTCb/fj8lkIpFIAGAymbDb7YyOjhIIBBjqfBXr5L/y/Sfy9J5/1rpLpjeY6Nh6B9ffdh9llbV0Hz8wy7VDBbWN7SxtW08sHCCVPH+HrDf7IMzki9++Zj2f+G9/SN3SJg7tff2yWk/mSy6bJhYeQ69V0bsfDMYmFFVHLpsiFQuhqDrQIDTci+9omsBggNOHX5MlireQnbLOiiXh/zwBreufpXTNOrLZLKqqTgcEq9XK+Pg4RUVF1NbWkk5P1QOYzVMT38bjcWKxGLHJfkyjf89rh7PsPD73+cxm0owNDxCcGCeX10gkE7M6X1VV1m69laWtayku8fL8L37yriWTmT5OTAYnSGeylJRX43QXkZzHHqGXIxoe5fj+Z3AVVWF3hTFbXSiqfqqvhaKSSSeIhvwEx/uIx4KLvgPW+chgcdb+TviLv3+Gv/3fN5BSrsdkcpLP54nFYuj1epxOJ6FQCLvdzsDAABaLBafTCVm01zIAAAr9SURBVEwFi1HfMQL7/ohjp8b4P0/MT3WCpuU5uf83hCb8aFqOSGhmQ8XflMtl8fWcpKquEb1ORVV1l/0YM9DTyRP/8SMcThfRSOiy0ppv2UyScX8n4/6zw/bP9tAViAVX17IQyclv3ua2TU7+4qufx129DX/IhLe0ApfLhclkYnx8HLvdjqqq060j42N+dj//PXKD/8qR0wG+8xgF6d79bkorKkklk4SCATRNQ1V1FJdVkIhFCV/iXJ5vp6o6FFUhky5QO7E07+TkN+fROZBi166dVFlPU1s0SiwSANWOorPgcrsJh8Po9XpCwTHOHHkR/+4/INb3GE/sSPDPv7rSs31fXCwSQafT07ayA73BwGRgglgkRGqWjzAXomn5Rbei+GIjhMjLksW70KuwvgU2t0FHixlvzUaKKlbjLG4AoRDwn2Lfjl/wq1d62XEMxhboYloebwlbtt/KqH8YRVHY8dJz071Ur8TaINK1QQiRkcFiBsqKBGuWapS6QVUhEoejvXC8b966OpxD1emwWB3EY5EZzuotaF/dQf3SZlRVZe+u1xga7Gf7rXfy8nNPs3LDNiwWCwdef5lIeIFGOWlBkYsMzdBIQOPpPVdmla63E0JQXF7Hpls/ROfRPRzb/eIFezxW1tSxccuNnD5+hKce/Sn5s2Mampa3Mdjfi9nqYMPN92K2WIhFwux7/aXLjngGoxlncRmR4DjJ+BzPVMxUsNTrjaSS8zsNoHRhMljMUKE+pDq9kbLqpbSs2UbV0hUM9Z5iYuT8s1tt2HIjdruDX/zHT8i9bfbvpc2tPPfUf6KoOob6uymvXkI2l7/sQCGEwqrNt9LQuo4jb7zIsT0vzWnLghCCto7NVC9t5+ieV+g9fWTO0pZmRwaLBS6bSePrOYHf14Neb0RVdVMjJt/yhRRCsPa6LfR2ncE/9M6l0SxWKztefm5qnEgmzQuPPYTT7cXvu/wJcPQGIxV1TZRVLSE45uP4vpfR5rKuUwhKqhqpbekgl9cY6DrxjkAoXRmyNWTB04hHQ5w+uIMT+18hHBx7x5flxlvvZPACiwdlMplzWj9SyTjh4PicfOnymkYyFkWvV+k6upvxkTlex1HTyOay2Bxu/AOd+HpPsxC7lF/rZGvINaCiqgar3c6ZE/MzjPx83r7KuqrTozcYSSXi89O5SQjMFjvpVOKSlm2ULp8QIrPoJ7+5mun0euoamq5ooIB31t/kshmS8ej89YLUNBKxsAwUBSaDxVWsrqGJY4f2FTob0iIhg8VVLJ/LEpqc3fgQSbpUMlhctQSx6NwteixJFyODRQHo9QbcHu9lpqLhH/a941WhKFRW12IyW857lre0fHo9lLczGAu0boF0VZDBogCWr1iNzW5Hr7/0Riir3U77mnV4vCUsa191TtqxWJSSsvJ3nFNZU4feYKCssvq8aba0rbzgNT3eEppb2ymtqKRxWesl5126OslgUQBCCAb7emY1ma7Vdu4iPHVLGjmyfw/lldWcOHJw+vV8PkdldR39PV3U1Decc14iFkNRFIYH+7HZHRiMJhxO9/T+t68parXZz/m5oqqGU8eOUOwtveItMFLhyU5ZV5gQglg0QmVNLcHABGuvu55IOITV5sDucGJzOKiqrcdqs1FZU09peSWqqrJx600M9veysmMDqqrStmotmUyapS2t9HadJp/LYbZYsVhsnDp+mGXtq/CWltNz5tT0dRPxGA3Ny0gmEly37SbCoUnCkwFWr99EMh6nY+Nmuk6dZPX668jncmzYcgNDg/2s2bAJvd5AQ1MLqqJS29BI15mTV2YUnbQgyDk4rzCLzUZVTR3+4SHqlzbjKvJQU9dANpNGCEH7mnUUebwEJ8ZoX72Ona88T0VlNb1dZ8jlcxSXlOIfGsRkNjM67CMYmMA/5CMcmho5WuwtJR6LYTSZpr7IQjDmHwagdeUaxvzDeEvLSSXiDPb34Sn24vYU03nqOFW19aTTaXz9PXhLyhgdGWIyGKCyupZgcAKj0cSpY0fQGwwcObDnslY2l64+Qoi8fAy5gsxm69nh5jayuSx1DU2oOh25XI6yiip8A32EQ0GGfYP093YjEBiMRsqrqslm0qiKQkV1LalkkomxUbyl5UyMj06n7x/20dDUQiIWQygK4bc0q1rtDlRVh8lsweMtJZNOIRQFq82G3mDA4XITi4QpKi45e80a0qkUiqJS5PGiaVMrm+sNRlLJBTQVmHTFyO7eV1hJWQU2h4OeM6fwlpYTDk2iKAoGo5F8LofD5WZ8dGpa8GQiTmV1Lf5hH0XFJaRTSTSgsrqW44cP0Laqg6MHz+2UpTcYqGtoJDA2dk4gsVhtVNbU4hvoQyDODvs2kM1mMBqNxGJRDHojiqpgMBgJBsaxWGwIRSGVTLCksZnD+/fQuqqDYwdlR7DFRgiRQQiRYmpkjtwW+KYoigZo123drglF0dZu2jrv1xSKoqmqqq29boum1+u1tddtKfj7ILcrvwkh0rJkcRVpWtaG3emaHsh17ND+eZ96v331WowmM3ktDxoc3vcG2XlY2Eha2GTJQm4LZvN4SzQhxHn3KYqqNS5rPe++DVtu1Kw2uwZo6zZv1Wx2xzn7a+qXattuuU3TGwznPb92yVJNp9cX/P4X+iaESMsKTqngLFYrn/rClzBbrNOv2Z2u6f+7ioqIhKbWJBHKuR9ZRVEor6xGKAotrStJv2URZ1XV4XIX0X3m1PQyBW8/3+kqumDLztuPX8xk06lUcJlMhkN73yCbzeAuKkan02GxWMmk01TXN2B3uNA0jWw2y/Xbb2Wgt3t6btGSsgoQAk9xCbFYlMG+HixWG06Xm8qaWkrLK+k6fYL6xma0fI6NW2+kr+sMFVU1pFJJquqWkMtmsTuc6A0GTCYzTnfR1L8uN9dt3Y6vv5eKyhoQUFVTTzKRIJvJYDSZ5mWt2YVI9rOQFox0OkVNfQMVVTXY7E4MJiNllVUM9HTRtnotOr2BaCREPp9ndGRqaXqnuwhV1WG2WDAaTaSTSQLjY6zo2EDT8jaCE+Mc3LuLxpY2zBYrE2OjRCNhLBYrKzrWo9PpKC2vRK83YDZbGBrop25pEw6Xi4qqWtKp1PRask3L20glk1RU12A0mfCWlaMoKpHwwl6Fba7IfhbSglJRWUNfTyeJeIxMOo2qqMRjMeLRCNFwCLPZes7guaqaOgZ6u0gmElPzeghoaV9JPp9jxDeIpmm4izyMjvhIJhOUVVbiH/JRVbcEi9XGsG+Awb4e0qkUwcA4LW0rSMRj6PUG0pk0E+OjBCbG8JaV8/qrL1JWUTndbNy0rI0R30Ch3qqCkCULacGIx6Ikk0mSiQQCpor5uSyB8TGymQyR8CQebynBiXEA8vk80XCI8VE/2Wx2egav4cF+DAYjldW1xGJRQsEADqeLwPg4DqcTk9nMkQN7SCbilJZXcfLoQWqXNNLX3cnGrdvpOXMSvd5AYGJ8qjfr8BCR8CT5fB6z1YYiBL6BXiYDEwV8t64sOQendM1qWt5O16nj5GaxrGLz8nYcLjd7dr46jzm7Osk5OKVrlqZpswoUAAaTiWgkPE85uvoJRVGS+XxeznoiXVuEQI6KnTuKoqQUIcQ8TcksSQUkA8Wckq0hkiTNmAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiAwWkiTNiE4I0amq6tJCZ0SSpIVLCNH1/wGOFRf0P85NKgAAAABJRU5ErkJggg=="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydCcBNVdfH9Zb0Nr/NyZh5zEyGIg0KDUoTpUGSoURJEUJUpEgZQwgpkjQqQxSZ5zkkDSqNGtDwrd91t++6zrnD4xnuvc//ZHfvc88+++z9O+fss/dae62VI4c2ERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABEchiAkdk8fl1ehEQAREQAREQAREQAREQAREQAREQARHINgSOsO2EE086mXTcCSeeeOxxxx2f65j//jdnzpxHH3VUzpz/sY08+/bt3bvru293rlu9Yuk/f//9d7YBpIaKgAiIgAhkawJSWGTry6/Gi4AIiEDiEch/buGiufPkK3DkUUcdtfPrr3Z8tnHdGk3QEu86qUYiIAKZR6DtQ91679796y+jnu//ROadVWdKbwJ58hcstPOrL79AAJneZas8ERCBxCNQsVrNCx/q8dTAd954bcKeP//4o0iJ0mXzFSxUJPc5+fKfduaZZ6OYiLXWg5/u3W3Ys0/0iDV/RuRDidJ/xISpfN57W+MGGXEOlSkCIiACIiACEJDCQveBCIiACIhAQhCofmHdyzp069P/3CLFS4ZW6Kcfdn0/cfSwQQjq9u7dsychKqtKiIAIiEAmEahS48KLhk5880P6v1ol8568d8+ff2bSqXWadCRQvvL5NUdOeW/u0oWfzL3z2noXpGPRKkoERCABCRyd65hjBox6ZVq1WnUuiVQ902P8/vtvu3db1/4H/fxff+3b949t/1pyx7Gv18PtWm5cu2pFVja1RJlyFce//dHiX37+6ccLS+c7JSvronOLgAiIgAikNoGjUrt5ap0IiIAIiEAyEKjf6IamvQYMH0tdv/lqxxdrli9ZyGStcLGSpQsWKVaiZfuHu9eqe1n9Vk2uvoxJUjK0SXUUAREQgfQgUNP6PsrZvH7tKikr0oNo1pRRvc7F9TjzGWflPidraqCzioAIZCaBJ18YNdEpK77/9puvF8+fN3v96hXLPt+yeaONdbd/t/Obr3/+8YddKCgys16Hc64KVavX4vivd2z//HDK0bEiIAIiIAIiEI2AFBbRCGm/CIiACIhAhhI465w8+bo+9dxwTvJMry4Pjhs+qD/KCndSzOl7PTtsTKnzKlR+fOCIcW2bXRcQ3mkTAREQgexAAOsz2rl4/tzZ2aG9qdrGIsVLlaFtG0xgmaptVLtEQAT+nwDxKPjrX9uuq1u1tK23+SHZ+ZQpX6kqbdi8Yd3qZG+L6i8CIiACIpDYBP6T2NVT7URABERABFKdwF33duyC2fyrY0cMHjN0YL9QZQVtX7Jg3pzbr7201q7vv91Z86JLr7ioXsNrUp2J2icCIiACECCmT6GiJUrxfdWyxZ+KSvISwHc9tV+zYumi5G2Fai4CIhArgcnjRg4l74Y1K5engrKCtpQ6r2JlPrPaNVWs10D5REAEREAEkpeAFBbJe+1UcxEQARFIegJHH50r16UNG13P6rORg/r38WvQN1/u2P70Yw+3Z3+zlvc9mPQNVwNEQAREIAYC9a+98RaXDTciMRyiLAlI4PgTTjwpd558BaiaFBYJeIFUJRHIAAJlKlSuRrFLP/3kowwoPtOLPOnk/52SJ3/BQpx43arlSzK9AjqhCIiACIhAtiIghUW2utxqrAiIgAgkFoFipcqUQ5AT9Of7RaTavT/99UkE4C5bscr55+TNXzCxWqLaiIAIiED6EjjCtvqNbmzqSv1y+9Yt6XsGlZZZBIqVKluOc6GcN4XF4sw6r84jAiKQdQQYr3L2pQs/mZt1tUi/MxcvU66C68dMYbE0/UpWSSIgAiIgAiJwKAEpLHRXiIAIiIAIZBmBc4sUL8nJd1nkwWiV+Puvv/6a/9HM9//5+++/Tzjp5JOj5dd+ERABEUhmAtVrX1zPrcr/bfevv/z+22+7k7k92bnuxUuXLU/7t2/9bBPXMjuzUNtFIDsQOPKoo44qWaZcRdq6fNGCj1Ohza499GPWjf2cCm1SG0RABERABBKXgBQWiXttVDMREAERSHkCJ5p9OY10gQmjNfiJLh3aXFu3Sqn1CloaDZX2i4AIJDmBJs1bt3NN+OarHREt0JK8qSlf/RKl969MXrtymawrUv5qq4EikCNH0RKlz2Ns+9WO7dtiWZSTDMyKlz4v0I+tXr5kYTLUV3UUAREQARFIbgJHJXf1VXsREAEREIFkJvCXmU1Qf/MKFZPFxC8WtZCUzG1W3UVABEQgGgGsz86/4KJLXb6vd3zxebRjtD9xCRQvs1/Qt27lMvl9T9zLpJr5EFj2xQGjoJyW5W9L/5C1fN4TxcyHQNkKVQLxK1YtXbggVSCVLFs+YDGyetmiT1OlTWqHCIiACIhA4hKQwiJxr41qJgIiIAIpT+CrL7Zvo5G58+YrcNRROXP+9de+fSnfaDUwSwiYwOUcOzHClm9NyPJ7llRCJxWBGAk0u+e+B8m6588//mCV7tdfbpfCIkZ2iZbNLt+xBQsVLU691ipQbaJdHtUndgK8P4ta+q+lZZZQXGjzIeACbqeKNQIW0S7g9qpli6Ww0J0vAiIgAiKQ4QTkEirDEesEIiAC2ZEAq9EsHWPp6OzY/ljbbEH7AqtNc+Y8+uiCRYqViPU45ROBWAkEn8UjLX8ZS2UtlbTffMc/wfw8v/8J+R7r6ZRPBA6bQN4C5xZu0OjGW4h1sGDurBkU6JS7h124Csh0AuZGpfx/jjzySAJur1+tQLWZfgF0wvQicIQVRCpt6dT0KjRVyylboXLAwiJVFBZmXVGJ9uzdu2fPxrWrV6TqdVO7REAEREAEEoeAFBaJcy1UExEQgRQhEDSdp389y1J5+/uEFGlaujfj22+++pLgfRRcsVqNC9P9BCpQBPYTQHHIc4iQhVWi0bbjLQPxVXJFy6j9IpDeBO66t2MXBNwTRg15zhbnH0f5+EFP7/OovMwhUCIYeHfb5o3rf9u9+9f0OutJ/zvl1NPPPDt3tPKOsC1aHu3PXgRsXJorDQtqUPxzLzG+PTZ7EYuvtTybKJ7N6+lf61atWBrf0YmZu0zQxRXKin379u5NzFpmTK2Ci1eOCF3EEuImLWNOqlJFQAREQAQCAw5tIiACIiAC6U+ASd0plgpZCgictHkTmDfz/bfZU6P2JfXESAQyiEBBKxdlxbeW1phLqID/7fAtZAKKYIY8/2ZQfVSsCHgSyFewUJH6jW5oinXFuGGD+p+ZO09eMn71xefbhCw5CZQqWyGwMnnV8vRzo3LhJVdcOWPJxq+mf7JyS7VadS7xInPaGWedPeyV6TMXbvl+z7VNbm+RnPRU6/QmELQwPMnKjXdsyrgWN1DrLO1O73qlUnnOuuKzjevW4NYvFdpWvsr5NWlHqliMxHlNuPfPtuRci8Z5uLKLgAiIgAikhYAUFmmhpmNEQAREIDqBYywLgiZWdseyojt6iSma48N3pk2haVVqXlj3eIu+naLNVLOygECItRORQX+wtNZStPgVzu0F1hUaJ2XBdcvOp2z94KO9nHXFzz/9+ANCZ3h8/eWO7dmZSzK3vdR5FSpT//T0+97ukR5P4krx6KNz5brPvnvx6T/85SmVq19Qh/hQlavXqpPMDFX3dCXAew1lxfGR3CN6nJH3KHHGTrckq50IlyTV4lf8xzanhFmzYsmidL0bk6Mw4r6WtHSeJazntYmACIiACGQCAU3EMwGyTiECIpAtCbBCe7Ml/LxmK9PpeK/28kXz5+EaCsHLxVdcdW28xyu/CEQhgOIBoW8eS0Us8WxG2nB1gWCG51bPrm6vTCOA66BLGlzTGLdBWFcQbPu4448/AZ/hP3z/7c60VAQl8Jlnn8O9ry0LCHD98p1bmEDFOVanY6Da3HnzFXDN2fn1l1+EN417xwlN2bd4/rzZWdB8nTIxCSB8ZXEIbhLjUTzwbsRVIkG34zkuMSlkYK3KlK9cleLXrFiaEsL9wsVLlTnOXia0ae2KZYszEF2iFo3FrbO6lavQRL1KqpcIiEDKEZDCIuUuqRokAiKQIAQwAWdFN5un+5kEqWeWV+Mf295+fdLLVKTh9U1uy/IKqQKpRoBJNooKVsWxMhSXFpE2F7uCfIFn11xIpRoTtScBCbBqnngDL48Y9AzWFaecdtoZVNN0FV8TsDneKrMC/+W35iwaPumtWfEeq/zpQ6B46XIVWJ1sXmF+37R+zar0KdWUH0FB6OYNa1f37HjvIe6e9u75889N61av5Hyfzp31wesTx7yYXudWOUlPAKU97zeUDvH0Kz9b/m8s/eTejUlPIgMaQB/urKpSxX3SeRWrVgfVH7///tu2zzauzwBsiV4kzwqW87iEksIi0a+W6icCIpAyBKSwSJlLqYaIgAgkGAFWotW1dJElAvhqi0Bg2qSXR7O7QpXqtQoXK1lasEQgnQgwyeT5w9JptaUvLXkqLILuo1x+3GUwOdUmAplCoHrti+tVqVm77i7TTrw0ZEBfTnry/049jc9d36XNuqL2ZfWvIibG99/tRMioLQsIOMHl2lXLlhCAN72q0OPBNs2f7Prgvc2uqns+90x4uSi4brmybrWbr7igUqtbGtVLz3OnVxtUTpYRwHIQ14i4LI3VUgIlRylL9S3lt4RrKG0eBPIXKlLMDNtORriPQjEVIJWrXK0G7diwZuVyFhmlQpvS0IZf7RgWEZyZhmN1iAiIgAiIQBoISGGRBmg6RAREQARiIIDCglU4WFr8FkP+bJ1l6+YN65aZaygg3NDsrtbZGoYany4EQhQQxazACyyhqNhg1hKRVpQilMF9FMdoUpouV0KFRCPACnysK8g35One3X7/7bdAQNsTTjr5ZD5/+P47gsXHvRGYmYNWLlk4P+6DdUC6EDiw0jod3UFRsc+3bN44cdTQ59y94lVZgv2uW7V8yT9//x3Nqixd2qpCkobAKVbTfHHWFplBNUu4l+N+kgzBB2DZ8pXhlGPtyqWLU+XZO6/SfguLDWtXLo/zvkmV7Cj2UDgzRsSlmjYREAEREIFMIKDBRiZA1ilEQASyJQEUFqxAYwWb+toYboHXxr44hGxXNLqxKX6/YzhEWUQgGgGeP5QPBSyxqvT7KAfg1zuvJZQW0YJzRzu39otATAQaXndzsyIlSpfdumnDuikTXhrhDjrBlunyffcvP+OCJe7NCZmksIgbXbodUKpcxUDA7ZVLFy1It0JVkAgcHgHGVyyo2WEK/HiUWSy+mW1pjaV0sxY6vKYk3tFlylcKxK9YsfjTTxKvdvHX6LQzzjr7nLz5C3Lk5vVr082tXfw1ydIjsLjFQnetJY0Ns/RS6OQiIALZiYA0xNnpaqutIiACmUmAoIS482CQi9BJLjmi0J8xfeqrHbr26X/Kaaef0eDam2995aVhz2fmBdO5UpIAz+FGS7kt4Roqmr9u4ld8ZgnTf5I2EchQAhYb+dhWD3bpyUkG9On6UOiK3P8ed1zAneDu3b/8Em8ljrVjnZBp7cpsGSQ1XmTpnv/kU049zV2DNcuXLEz3E6hAEYiTgFkeOhdQWHEdzd9RrA7dGXh3/mkJl53bLWXHOAYx0S5VrlIVMjqXfOYZavfePXv2mEe4ff+aO6XQeETEuzjCLOyOPPI/Rx51VM6ciz75aNY7U18dH9OJLFOFqjUuKF66bPnxLw4eEH4Mbqns3/++/mrH9ngsPXgnHWnbb7t3B8ZATvHN943BuDix1O/U0888q2K1GhdQB9qFVVgsxyVoHsaSuET7wpKUdQl6kVQtERCB1CMghUXqXVO1SAREIDEIMLljFRsD9DS580iMZmReLfbt27v3dVtdfGfbBx65vlnzVumhsLAZ4FFM2n6xALap6nf33CLFS5Y8r3wl5r0fffDu9J9//GFX5l21hD/TqVbDwpZwf/GDpUgKCwQ5+CdmYkpw0T0J3zpVMOkJ3Hr3fQ+ccVbucxbPnzt7zox33gxtEEGz+Xvv3r1x34sFChUtTp+AO6lvvtqBkCXmLW+Bcwtf1/SOu0cOeroPwb/DD6TcwsVLlTF5VO4tm9av/ebLHQgwD9nIV7ZilfNPPe2MMxd+PGfm7l9/4bmKe8tlErRcuXIdY4YmP8Z6cI06l1xe57IGV5/8v1NO/earL7+YPnnCmPWrVyyLdvxd9z306GVXNrrh4dZ33BQeJPusc/Lkoy07TQL4/bfffB2trNLlKgYEl+SN9xpEK9tv/3+PPfa4v//+52+Cbsdaxtl58ua/6vqmt48dNqj/b3aRQo87Otcxx7DA2sKgfIWLqWhlcq2q1LjgojPPPifPFrMYWvrpxx9FO0b7M5UA7zksgHF5iED6qzjOzvuURTgcg8WitjAC3P9FS5Qqy8+MzUjxQDrF+pdYFRaMbweOnvTmccefcOLMd96c4voYnueHevQdWKtuvQa4G7TH9vcX+vXqOnbYc0/71SX/uYWLNr2rTfuL6jW8hkVD5Ftlbuw639u8ablK++NXMIbevH5NVAsLlOX3d+7V95qbmjWnjhxrupp9He5q0ogxajw8EigvrqCKWGIsKReLCXRhVBUREIHUJiCFRWpfX7VOBEQgawgwIcRk2FlVxCw4yJrqJs5ZX3t55NDbW93/EJO8ytUvqMOqrHhrh5CswXU33dq46Z0tzR1HFSZsCLomjBw8cNizT/aIpLhgRdjQidM++OmHXd+3ufXaK5joufOz+q1l+4e7X33jLXfYSrm/Rr/wzJMTRw8bFKl+1OWZFydMRXjIZO2zjetwpXBgu+Ka65u0aNepKxPE96ZNfuWprh3vRXETS5tZudv1qeeGE6jX5d9lUqWmDetU9RMgxlJuiuVhgonPbVxBESgyWoBRJqNFLSHgDayIttWnKYZEzUkUAqefeXbu2+5p15E+6ekej7QPrxd9Dr/FEjC5SfNW7Vo/2LUXgqE/LLABfQ/HIrCfvXLbAVdoFs7gb5SaA/p06zRnxtvTvFg8+uTAYfS/5q58yXvTXpsYmqfuFVdd265zz6fy5CtwLr+zcrdv94fahfeFl1/d+Gb6tgIWgJZ89EnNrr64umlPcKsRdUPwfkuLezs0tL48T/6ChThgx/ZtW559/NGOH779xmS/Amh3t37Pv4gAPjTPzXfecx999sAnuj8c6eQt7+/UzZY7H1mtVp1LnMKCPvb+zj37Fi99Xnl37Kz3pk9FmEdgXb/ynMJitYd1BfFFbrz97jYFCxctARsTKD6KUicqGJ8MrLRu3fHRXk64+OrYEYOf6PJAm1jK69z72cEoeL74fOtnb02eOJZjELy2fahb72ub3N6CFdesCn97yivjejx0bwsvZQjcb7itRZvWDz7a0+SnAVdmbCi9nnvysUdiqYfyZAoBXJSeYwnXh1GVbiE1QtmPsoJjGaMEgm4TK0rvyP+nVKLMeRUQ0tPPDR/wVE/7mpO/6cvtX04+jzyKX/b/zf94tswIYzf9W3h/G+mOwFETygry0OfzWbRkmfOGTpj2AdZd7lie35btH+nup7Cwfqjt/V169T366Fy5UFhuMisKFBi4tnrupdfecmVv+2zj+kgxczifGVOcMsTOT1/Je2uVucI7x94VjHHv7/J4v7kfvvdWqIVJptzx6XMS5nE8L8R/ya5Bx9OHpEoRAREQAREQAREQARHIOgKY2FuqaekBSzdaOjB5z7paJc+ZB45+dbox+7ffsHG+Qim/1jBZGj7prVkc79LS7T//476jcIhEAqGWyxtqBo8A69mRE98ILZfvocoCr3KZPLpjsBwJzdOs5X0PhpfnXMNEu1pMiues3v4Dx89b9+XPo6a8P2/Bpp2/8zfCxmjHp/p+hCiW/mOpsqWnLfW2dF2IO4xDENi+Iy01sNTBUiVLOYOBu1Mdl9qXRQR69B8yOtIze0OzFq3Z3/7Rx/tFq+LQiW9+SN7FW3/YR5/w6eZv/wjvX9zfi7bu2nvZldfd6Fcmx5O3+oV1LwvNc+/Djz3hVSblYZVBXtx/uD6cvvedBWs/d33wI737vxCtHewvVqpsubfnr9nm1Ycv+fynv6vUuPAiv3JQVLjjxr4569Nezw4b896i9Tvcbyhc/I5FSO/yVa99cT3y3dKibQdXf849Y8nGr1weFDeR2oOwj7yhfT+CSuoUzpHrla9gIRSscW0oClo90LlH6HvOlV24WEnc90TduEYcU/fyKxuRGavEcdNnL/S61iXKlKsYXiCLAh7rP3iUyz9pxvyVU+cs3eDuR1Z8R62EMmQKAbsm3OPXWrrV0gEFXLST8+601NgSfcDDlk7j/ah35MHkmt7V+n7uexaTRGN6uPvrX3vjLZyLZ42yChYuVgLlNL9N/2TVFqwlUDrc3rp9J7+xKm5Yyb9wy/d7UFw4JTnK9Glzl28K7QN4xiPVmWNHvz7jY46h/y5iVnjkR1nhxqdO+Xy4bc/s461Nx1liPHm+pQK69zP7Cuh8IiAC2ZWALCyy65VXu0VABDKawOl2AlaWsiINP+RpcoWR0ZVMxPJxC1Wr7mX161xa/yrcSuz8+ssdsdQTZcWLk9/9qJDZ42MZMezZJ3pMGT96OH54mUTe90iPJ5u1bPcgq8ycb97wcnFfwm9YObDKzO2/p8Mjj7EiltXLmMmzihVB0ZWNm9y2cN7sD/3q58pj/9oVSxe7fOdfcNGl1Ie/WX3LRJNA45T3Qt9ej0ZqL25JBr/8xvsIBhfMnTWjU+vbb2LF9IWXXN7w2ZGvTGOlbCy8skEeVqfjyoC4FKwIXR7FVzduMliVSBBSXPCwiu4om5gyVsIdAEFK+c7vuEbBjzF/88mqVVa0c05WorL6lHLYz+/OpQ9/k9flcSv1yMNvviv3tIo1te5YVt9jCYabpEFP9ejs1TpnDeZcQ0Ui0PbW665AMMTKXo5DgYFgv5O5NsItDxYLCJT+tmWvuCjy6wPpc92q3R/Nn5Q7JwpWrN/4+7VxI4diEVDqvAqVEcpT7qUNG10/bdLLowePn/o+ffDHs2a8g+UFfssRdNG34UYq2lWEi63QnSHjOH0AACAASURBVEEdzPX6NiwqcCPCkuTHnn5hJAqHltYf+1kjoHTmHG+/PullLCD4Tl/5wstT36O+Bc3aza8ORUuWPo999P+LPv5oJtYFTlk0/6OZ7/d+uN09rIJGicHvWJFQP6/yeD+UqVC5GvuchQWK737Dxr7Gu4Rz8H7avvWzTax+Rklwi7lkefyR+++Jxsjtp7zH+r0wkvuI33hXTps0blTNi+rVR6ldrsr5NfnNbjHfoO1n5c6Tl3cKxxMYnNXY8C9ZtnwlrEde6NfTLD8+mnlexarV/zFzmnWrli8Jrx+KLK4vlhdd77/ntvfenPwKSowx02YugHnVmnUunjpxzIuxtCsoAGfcRH94wBWa+r9Y6MWUB66MT3nXEMfCcwtTRPDO4v3HKn6UarzfsHrinfmL5cV1He87xrq4QqVsrFNdYr97X/KOpQ7s4/ryN67eOJby2HiP8s7dZoljuR+oK7/zDuU79zTndHmpE+d171fO4VxA/ptZ94+zqjoca6kgg6gf59e66BIyfTL7g3dxw9R/+MtTTjKLOiyTH2jR9FrnQo8xq1dhWOUxNsZKrt0dN15FOS7fd+b3Diu8fkPHvuZ+ixZEvM1DXR9noc+Pu77/rnnjy2vTf3Msbgm/+mL7toJFipU4wxQhO8ySK2rjEi8Dz8wVlnC5+lbiVU81EgEREIHUJCCFRWpeV7VKBEQg6wkwAWNyV8BSwK2HttgIYDKOAJ6J12VXXnvjmKEDo64uxsAeiwwEZUy07rn56ktD3S+9NGRAXyZmuHyqUqN2Xdx5eNWmVNkKlfgdYZUzfUfpcEfrDg8jYGrbrHH9T+fO+qDLEwOGIswqVqpMuUitKmVCH/YjlFw8f95sviOY6vHMkNEItAY/3bsbipV6V113U59BI8cjLKTdfnEoEAI99cJLr5Bn+aIFH9/brHED50LKTUpPN4fjsZFO+VzHWQtZ2bvVEj72Pf3sh1DAbzN+vXGVgdsa/Hs3sARPhCoIanDzRj5c7DCBrWBpgSX8viOQ4e91lrjW2yxdaamyJVyBrbDEuAt3U5wHYc1OS5stYYVFPlwOEPOGfdQBRQbKkT0mFEIgw++4JnCKjQMxOTJLIGPn1naYBHj2O5qP8f19wOPdEPB4FYmAmN9d8O1Ip7UwF3ucD3PKNUFxoO9ZsWTBJ/SJsVbZ5PkEFg1sP+7aFagXfeC9nbr34fvwAU/2fKHf4135jrsPl9e8+JV5ftyUd+mDUcDgCsi5/nAuraK5tqL/w5INZcWSBfPmtG9+8zVO6GY3/h/PmzIXhQXCcxTU4fE1ENoVKVE64D/+rSkTx7m6Ucb9d950NdYXUyaM9l35XLzUfpdPn21Yt+bcosVLPtSz73P8Pf21CWO6dbjndqdAsrLHorAg9giKZi/lD9YS1BEGFnB7EeVgkYGygvq0bXZd/ZVLFgZ8oTvXYBUsQG2s14lrjIVO/UY3BJQy+L1//OH7WlIXXDuxr3PvZwajBLnqgvK4ufPccH3FDhT03Ce9Bgwfi7ICN1X33ta4gXOLtXHtKvqvQ7aaF116Bcos2HS8p9n1Lg4Lf69duXQxCgvaF2u7LB99JO9V+m6E2ixY2GL9H/1xqBD6oCLV/8VMGL70B7yreNdt8jmSdw/v0AKWePdxHMo+rHZOtoRrqJqWeD+hPHDjDq4ZcaDcuwtFFWNg3qHh1k1D7TfuXxQVXu4aGUOjsODd97ollBoFLSE05v3IvYGyjXcx7kNx41grWM9P7JN3K4sVsNbiveqUGryrUWKku2uf0uUrV7WycyxZ8PEcPjNyq2yxYih/3sz33m7/aO+nCxQuWnzpwk/mMk6NFm8GizjXpw8z11WhygpX57mmKOY5ZtzJb4w5/dqDNTF9DftRFDtlhcvv3mEEIM9IJhlYNvc/9xr3oOZ0GQhaRYuACIhAKAEpLHQ/iIAIiED6E2DihVCRCRoDW1zTsDqNxEQJIRQTbz6ZMDmho5uweQYGTsYJOS5NChYpWuLJRx9sG6vfWqwYZrw19TWCvrJqNxaFxR2t2neqdH6t2igZwpUVXF7ObTKcTSgsEKh5KSxQJDhzdbcfn77d+z7/IhO2/j27PoSygvLWrFi6CIUF/uEj3T7OfcbHs95/xykWOnTr0/80UyrMfv+tN1BWuPJcOZTpp7C4/tbmrVi1i6DugbtvuS403oUtoGYilcOMS3x9qqf/rZ7QJSJIIeg9PPwEIqENINYFyginnODZRFCDlQYrr/3GTAHXMSEbQp1rwn5DiHpT8Le59olQJXTbZn8U8KCJYgThEArQkZZWWyJwML8jJMJ6hDr/an0Mygz8WdP3oAgJCGUsudgdAeFMFCsTjyqkz08+rkPo81xyfKkzq2uddQp/I3RilS2/IXQK7Ue5tgjWXOwXngOEZvS3lIOgk3shvF8lP4IY1wc7YWiG978IznHVgVL1lZeGP+9H2HSkgTaZTDyuQCrEzEHov+v7b3fGG8+G/pFzIvD61gTYWE/gZo7V/B++M22KU1aQ50TrrFzdL2147Q0I0bE4QEEc2ibnLsoMOyLGrzALilH00QjJ77v9+obhioDPt27eSF9Of8xq3XABGopcF7vjz7DYEgjjRzzX9/FId3PJsvvdHW1ct3oFdcGyBSu2bg+0uiM09hEKJlYlw+S/xx5/vJfCwllXfP7Zpg0orLF8Q6CHFQLxkUKVPaw+5rzxCPaJL+GUFbwjn+nV5UHXtv+ZqY377mdJ4/ZXDrrXmjfz/bdRnFMm902LGxvU/WLbFgS+vhvWGMS/IMOo5/s/ER40/lhjw74/ft8dj5CS5xHhMiv1uR4kFMUIpOn3UO7yyTNN3tAxVKTqHta+KP2XK9v1Hc7iDmE7fRD9Ff0W/RfCfMZ+7CMf+0jOeoDvtM0JRTmOfCT6A8qjv3P5XH8JB5fXMTkQtylEOM87A+UC5UUav7CfPhdlE/m5hhxL4v4KBGYOtoc2uc1ZSbh9keKo3B1ynNdX2skGiyZR8qJ4m2GJY6pbusESixQYA0yxhHIV5lh58X7AVehs++Reoq2wO6Tvj2fcTdwIYothhRWPkjhKuzx306eiMMWamD6x0c233YV1HZYV0ZQVFIgrqKNzHXMM74dRFtvH6yQowYlpwdiYMenWzRtYjOG5te/Sqx/94Zuvjn8Ja7TQTPTLWHLRZ36+ZRPX45At+HwxFuBe4r7jevA397CzePV9R8dznSKcn13O2jU8G2MwFGRYSmuMnZabVseIgAiIQBoISGGRBmg6RAREQARiIMDECDdQTNgRnDHoxoQe4ScDXvYxIGelNZ9M0EsG87FamwE6v7OSLOBqxgb0CCLZx2SXCRbnYALLIN65pnH73OQrsDIqmMdV202m+ZvJL5sz16euzl0Nk0Rn6s8Ej7KdEDRqoEVcHhFQFuHOU90euu9fm6y4CkT7/ODtNwIKC7c6M9Lkj5Wsd7XrGHCjhAuS8MDW7lwmM0FwmYPJk9f5QwOqIrwhz6133/sAgrFli+bPG//i4AHuuH9NesV3Atj6tQVhV6Fi+4V/c4PllatcrQbCSlbY9rTgpeHlRSqTlbwtO3R+jDz9ezzSgQDboefG7zt/b9m4fm00vtlkP9eZ1Zjc76wUd8/CIc23Z4t9CGKYiHJtnZuJLfYdYY0T2qQHugIehfgJpF3gTAREuOOh3yBv+GpU7u0JlnBBg3JkvCUUGzy3TrlBWypYWxEEco8gPKZPoa9wLq+YlPP8u/KdcjVcqO+UDKH9S6hihDJc/0HZ1BmBF8ch6II1G64h6FNwn4e7BfbR56E8gjv3OH0eQg4UQdQVtxXUk74U4RjXDOsUykEoRTBozs0x7lr+YN9ZHUp/yQpY7g3aj2CE830eLIf9bkWvc1liP6XfhnsiXOhQIorcSFYHe/bs4fr49ll+tUIZwr7VPq5AIrWmUPH9cQ9Ml7ISAdNNze9uSywE3Ej1eLBN89BjTTYXCIbNhqJg2qsvjw5XVrDPKYK3bPLvm3BrVLVWnYsRkj1sbqy8BO3Ux+T9fyAoP8mkg+HtCFX0nm7CvHivmlMwFzfTOFYMf2mmCh1b3no95w0v64jgqmOvANTkLRviDoog1N0tEDi/9+ncoXWosoLfjrLIu3yacDDwjoq2oVTALz35CHYeqqzgt3pXNXbKUXMXM+OAmxevcitWq3Ehv2Ohh9992tqxZbProykrOKZp8zb3404Kt19Dn3ki8G4K3YoGLRDjfCc5ASV9C4J7+gT6DxjRjxewRF/C4gHuAcZO/wsKPOkvYEgZbmxEn+PGOVxHvjvhvlOKupX3Li/jIPoW8tI/cG76JPZjneCEquynr0Nxh3UMfQcWfc4NIApvBOnUiRX/dS2VsEQfTN/DOI8+kP4J5RAuKTnfq5aICUNfjmKavsrFI6Gu9JVY53BP8QzynnDKEPpD3FTSd9BPIsDH//5S+2Sjr73UEm360X7nOXEKEsrmuL0mAP7L9lEv3hVu/IpVhuu7g8Ud+HjTvjUM/9H+dsw9duVYbj9GtFL1Osh+o41OmRGaBdZOOUabYI51I+8E3hfOBRXXjfchrPmN/ass0V7uO64xx8e1OXdQKyJYIsRVYITMjCXZvWbFkkUPdH/iGfrfxx5ofaeftV5oUYyrcSHKb8+byze/PowFO849IGNgv0VHvG9c342rwPBqN7BYG/yG9Qdu5mJgwPPB/ckzgoKS54dnkmvOd54vxgU8bzwf3KturkL53Mf0GW4/5QQWj1lyi1foK3jHM7ZzzzHn4NwcTznuuzuWe5nFK9w7X2XV4o8Y+CmLCIiACKQMASksUuZSqiEiIAIJRoBJNCupq1hyE0kmQJgUIyDAvQIuO5jAotRg8HyWRxsQUDJZZDKLANKtGuZ3Bu0M1hlUF7A02xIDasphYv+RJQR5TMYYfPMbg3wG/AzgCdTHQB13ERznVjQxAXf+gZn0M1nmePfOIF/EDWEKyoqfftj1/T1Nrr7US+ATqYDF8+fOZlUqgp7K1WvVwR+5X/57TIiPcgA/4W+8MpZV6J6bUy6Y9yjPd59z74SgBtcqnPvWlvc+gEDx8U7tWoZO1v536v4VrJF8g6OscAEMcTFF/lYPdOnJ53NPdH8Yv76uoq68SGVef+tdrXAxsnnD2tXTJ08YE95I58f84xA/xF4gbGLnhDIHCeFSZfIVslKPlZQFLCG8RygU6b7lnuceR2CxydI0S6ymY4L7niUmv+xjAozABqEPzxbPJhNehOPkRWjF8TzTKKtGW5ptiRWf7EewhfUDzzHPNArL6yzxLNIvUG6kjcm710YfEHr8zfY3KdKGoIbnn34BwR9te8USdUdgUyC4D2E+7WO1KsIszsWx9G0IhxD64L6FPg3hE9xwgUMAX9x90B9RNooT+p6Ay57g5ly+IJTEkoR7knJwm0VZbqX4CPtOf0m/hXAOlgjPeJZxA8L1ow2UQX0RFFIP2oeg0Sl4qS/XgHw8f9SLc28L5qVtlEn/yjFOEWxf02dDWcHzjgsffI1HKvXPP34LCHdYuRvP2fEjTv5oPse9ynQWFhtWr1iGi6U72zzwCPme7NrxXueeyR1HjAT3HWVE70fatwovE4sJVtfyu59LEfrvVh269CDPhJFDBvopndkfqR/Hwm7b5o3rcY1Szhi8N+21ibFyow64gSI/ygr6+27t77ndq48nHsgBSw5b4ex1jtLl9ruGQRFAjAqs6mZMf/3VqR7vqLPPycu4IMfOr77kvo+40bbOfQYMIdOcGW9P69utYyBmh9tw8UT8Cvf3p/NmB6wCvTaCYeOGi1XadS5rcDX3Ga68iHkSrR4wwM0i+Z7v27NLqLUfv6FAJ+gu12T5Yn9XMj7nYcyBezwEzvSjJMYi9JmMlVDM1rfE88EzfrEl+hnGCSgu2U/f6vp1+miedcqlf6Mf41jGZPRJ9GG1LdFvMPZB0M8+lAS4j6S/gzN1cq6PyMO7IPQ3+9N3u9pjD4oPF8QcYbvbGBdG21BucH6vmCx3ehxM3xeweLGNdyFtYjzIeADLPd5L9K8k4lJstDEBjAhYD3MUJLCij6TPxFUnlgv0k4wxt1nCYoJ3IPm4HpyDewm+vNvIR9/LNUNZgTKE/pj+Dd701eznvJzTWddxvfiba8q7hrz0KZw7VDBN3ej/KZ97hecKTpyDfNSDMsmH4oiyaDsbihv20fcT84FYLZ7WdsH8h3w4hUUa7ne/In1/R+nATlzgoQR//80pkz6Z8yFjlagbLtzIRD/79pRXDrjOCz+wSIlSZZ07qKUL/PuEG29v2ZZjGac7t4SuLCxBWrTr1JW/iR8XpXLw5lozJuE+5H5FScF9zvud54U+knECzyb9NeMF3uVYraK84z7m+rNYhfEDygXuQ/oFxoTcY9w/bpzHPck9y9iK+5Fz8SxyjLMg5DnhvmIMw71KH/CiPRfr7BmJW7Flx2oTAREQARGIkYAUFjGCUjYREAERiJMAkzUmkgx4mSgzCGcwziouZ/5/VUiZCDCZTIWvGmUQzcSYyQmJQTR53cZgmQE652GQzoSc8+GLm4koA2smYgz6OY6yELwyIWCgjlCPQT95mSQy+XYBEBmkM8ml7tTZrUwMOf2hXwkojbsKBBWtml592YY1K5mYxrWhJECYhxClYrWaF/opLDC/N7dRmP7nwG96JLdTCN/I9+svP3kGIHX+y/GdTr4mzVu3wxT+lZeGPR8uQEPQQ55ILk5YpUseAgxiqk87Kle/oA6+wgm2Ggrk7Dz5AuVhyv+rWV+Ew2LSiMKC30cPfvapUPck/Fb38isb1bYg5TCf/PKoYX6wg8oKhA1M7FgJysoxJnUn2j7uHa4zAjiEBtxHTATd/YqQwwnnEB4xaTyw0v9w/UEHFQ0IIALWK8Gy3Up+Z6bPM0QeZwXAd1cHvjs3P85FBc8P9z5McQHBPRwoy+obqrCBA88XXGZb4jkI+O+3fDxfOUJcgnAeVvIz0ee7ey6cVQG8OAf7nCsQ8rvVvK6NToEyyvY56yUmyzyvTIzhwH1BP8I14lpcZgkBDN9pEy4aEE5xb9Nmnmcm5CgcENJF2lw/4gRw5A08Sz4bbeC+8BKQRTlVYDdCovCN1Y4oTFHYOEEW7GgD9yNcYIKwCcESAgcEVTDnutBnYQ3FKlpYcQ04hvuUfQgt6L/cylmOQ4AWWF1sCWZcIwRs/IawysUIoSx3L9rXw99QJOC6A2Xs02YlFa1EW3BPH5zj1NPOQFAX81a+8n5FQiSf416FIYQ/14JRsM+8Ii29+Y5W96FcIYDsB+amL/yYKtUvvMj9hrLCyxVJlaCfdSwn/IK/1rv6upvoU1l9i8Dcr6HUD0E5+/2UxXM+eOdNhPoXXd6wERZ34X2lX9mFLQZHaHBzlN/uXRB+zJlWWVcH2hW+P5eZgJhnrYBijvfNjbe1aIP1R58uHVp7nd/F3di2ZRPPge9GrKYnBo2cAAN8xHe+965bwtvX4v79wkE23qME0vYrsNR5FQNCT9wwovD+escXn+PPPpYbDSsOrBVR8IffG7S/c59nA0qVyS+PHOriQcVSbkgenj2eS+qPVSrPLn0IYytn8UVfRJ/Nb/SRKGl5/lHYONdETshO0ShBef+zL9R1UWjVXL9J/0yf0NLStmCG0L7SWRrwWyQrgjibHVf2ePpip6zgBLSLhKUGzxNCWJR7CIMZHwQsbUPeefSRtJExKn0kTBHo00fTT6LMpt/mumAd4jb2OaE/C24QLodu5GeMyXk5fn3YsQfGF8FyGLOQ2FAqhO934wRXF4TSjOdoK+9f2uqU3twv/M07k2vNu4Vn2Smzwqoa/c8ywfgVaVEURy/94BzFzH8dv6Cs4Dln/BtLGVhEMV4k7xsTx46M1D+GWh0v8VFisrDn4iuuvJbyJr00/IXQOtCnD5s4/UPq+NbkiWM/spgYMdSRe4L3N4lnlXc373/GY4zn3HfmSoz3alvi3uR97hYkFLDvbqEC5TF2YDzLb5SBIpTnlncw9wfjB+5TrCewbHLjAvdcc07uD8ZbjCvYz/j+76DSgnpoEwEREAERyAACUlhkAFQVKQIiIAJGgAEuE18mfyeY0HMvK9bsOxO8GZaYGDGBQ4DBZPANSwinMNVnIMzgmcE3wiNcvTBpRtA52xLKCYR87OcYJosItJi8cj78x35siVWJnI/9rDRjUs+Ek9XmTPo4hn2sQGIwz8akwK0uRBlCPQOC3TABbzD7wR9MXh7rP3gUgqWeD7VtsW7VCueGwDN/pB+XLZw/D4UF7kj88hFHAmE+VgcuvoRfXreKNTxQq8vv3FcgVEMgdPOd99yHWxIvVxd5CxRiUpMD/+R+53MumpyQ7s62+1cq4+M9fJLofLxvtzgbXhPIqjVrX8xEE6HXjDdfnxR6zuoX1r2s96AXsSLIwWpbXLdEgc3kimvLGAChLwIIVstzTyGE4d5zZvNYCXG/4T4AYRECAO45JnwIihASI0xCoE95CB6Y/DMpZGLH/eaUBAhBKJ97jXuefTwjCBOcSwpWuCKsd64bUKpRDr+zwo1jEDggMORYBPOUR10KWOK+5m8mlAhVEKgy0cSPNoIJVj1zf39v9aXt1JdzcwwrQGkrKzkPEUKG+Eh2QuyDLFTsGLaACx+fzSs/WQOr6IPCIZ6/gKIkuNE+BHZOMUNfAEf4UWeYP2uJ5xs+1A1m9A11ggnFCgJs8qLo6BIse17wd/7knM6aAesIJvNO2cO52Vi1fDgb9UMwAHcEStxTMKFfRLhJ3+WEDu7aOp7OfQdt5n7lOO4DykGwQR0pxykZ2M937l82eDnBGdf3oC09rYuuuOb6JoVtZfmPZkGFRQKCdRQUFmt0d7enBo0IuE6a9PJorKVw84awybZ9JjPe99tvv/7KandXOSzU+M7Kd6y1ECyH1z38b/IisEeQTqydaPlD99PHOMXuulXLlgwaM+UdlMCmXAkEUw3dLEzCGS5OA5YDfsL9KjVrB1aL4wbJz/VI46Z38n7LMe3VcaPDrThCz4nPdrfi168fnzpxzIusICbvBRdf3pBYQbEwCBXOcQ1CY3WEH58nfwGeMVNYf8X79ZCtZJlyFVEuoMAhSDjfn+3d9SE/dy1FS5RGUJZjs8XuiFRXrBZ5r2Cx+EjbO5vgXz40P9YVTlkVKM/ei5H82TurQt7b5B/Sv3f3WPzfk/fqG265g89Xx744JHShAH7x+48Y/zpuYrZu2rCOMmPh7/L4+KLH5QvPMP0y7wCedfozxlmMe+i76T9oB/0YQk5+p79gDML7gvcb7rF4L/C+C7X08qoi7yW3IajkXUf/xDuQ9wjvmlmWCljC0gALMFZq0x/z/sRlDwJa+hvOh6ULfTd1ob+mP0JJiyKBRR20i++8Z50LGsp2QnWE/fTLvM+c0gUG9I30dyifaD99JjzcanDejWwwow/G+sq5U3KKWsqjL4UXdWcM4SWEpe3UgzZw7wUUEsFr5vrXSEpev32hio1gdQMfrkz3W6x/u3xwIbn3uVuswhiYd65bEMH7Y6UleNLH0vbwc4XWy/N7qXIVqzBmjGQhFrWQGDLwDnFKTrJjrReLCzfyMqYm1gR9SCTLZfKWLFuee9pc1e3+df2alcxXDtlqXnTpFTzzuIVbt2o5SqzARjychx/v/zzKCgJ6dzd3VZGa5vPcO4XWbrtWjIXcPcqYknEbzz9jSp5L7m36ZZ47ngMXx4ux0IeWeKZ4NjiOeQ/fsaRwCyXcfIrneqwlpwRl/sFzyxiJY2gj4wrqw7s67vskEgftEwEREAEROJiAFBa6I0RABEQgYwgweGbyyUTp2+DEyCkhnI9dXA28ZQnBm5tYMcHlbybnziSaSRam1AzMmUg5ITCDeY5j0onygcks+5msM5mcbYlVSNSBAb2buLGPSRnvAHwVs5LOrVQ7rMF341ub30PgUHzVvvvGawhX07y5yQ/CN79CLjfhIPsmjhr6XKQTseIzd558BcjDxCo8LytrCwbPg4KBOBNMtAY/3bubl5DJYtqiDMqxJUIQwqIl9wuhVi1b9ClKFyxPsBrxMtt3blj8ykPoRVkW22OyW9FLne++v1O321vd/xAT0Bf69nrUy91IaFuD15r7ifsToT7CEe41JutM9rg3uFeY3CGUqW2JSRr3IoJ1hBkIhLhPmMjhVoHfuAevsoQAb5sl3FxwP3J/M6nkGAQ+ztoHgUFAGGsbwhMUQEz+ELSECopYcYkSAWEUQhRWylE/JppuhStlUDfufawP2BAwUTc26sG14P5HMMHkk9+c0AaBEufGhQTl8rt7RoNFZPxHhKCRsHbKDie0o0JOsA3HbSGrYVHMsCFYGmiJfgKhLVx5zkdacisIEWbRT6EEQIAHF1auwonri7CZa4+AwK1OpVysFLBeoH/h/ChZuQ9QrnAO7jHKgC0CAYQdKFG5l6gH98QTlrhvuG7kp55uhax9PcjSxgnF+N1tAUVPlC2qgD9aAfHsR5j8+MARvi42XFkoQ0leZaPAMEOpX1Fy7P3zz4DCBgFVp179BhH0FCVwJJc95SpVq0H+tSuWLfZa/R+pPU45TJ+HSyOUEu+9OfmVjWtXha+MznGRrdJ1yoORz/f3tIqgX6p9yRVXcs457789zevcxLdwig/cQUWqn/XRgWcape4X2z7jeT1k22ZKZPpYFLm49ItdYbHfIo7t9QkvjYgUNwmFFPkQyHvVwbWHGCQX1Wt4TSR3hVjPwJlyIin47fV1bov79sdqGvrskz3CV3FzzVt37NortD5+QkaXp6j5jnLfidcxfcpEBHVRN97xtBFFxXvTJrMyP7Dhiqrns8PG8D7DWgN3kGm0rohUB/pD+gwSfSB9DP2Rs3ZjXMO7geTeJezjPUJ/gzBzsiWeLZQY9H8o3QtYog+j/6Rsxgnkpf9jTMXmxkf0nyh/6YN4n1DWS8Hv1In+ktXm9NckFqnwyeYs7FxZ/O3ccbr+b1m+qwAAIABJREFUj+OdEN/N1Z2w3ymQ+dtZmlAubeUYyqDObmEAdXXl0x7esXdZ4t7FhRB9dmAsGYxb8XlwnBCs7kEfnIP2Uj+4HdZ40esEmflbUFHtlNzu+qSpCsRSQwnNwplYrbrSdCI7yBbf5EfZ7Y4fN+L5Z2Itq1bderhSy0Fg7F3ffxuwHvXbKlSpXot9NoZd4OfW1ZU3851pKO0CruDu7dS9T/XaF9fjb5QpPTq2uSsWZXsMbeBaOeVTaN/rnhvaw/iFe57nhvxcV55PfmOfsxaiHBQZjGsYX7mxFWXRT3CP0x9wHBZIjIdRSDKeoY/guWFcktTPQAzMlUUEREAEspSAFBZZil8nFwERSGECDHgZCLsVQEf4DGyZSIYK1RhEH7RqMsjoQLwDH2ZbTGDJSrvQjRVBTqjjJfA7sOI7PQbdCExwfUEFxo94gVWGh7XhSokCUBywQjU8OC3CEXyj87uXu5LQk7PaE+EZv3kJhfBdzgpmBHz4QH962LjJWDO8PGLQIRNB3EQhsKEs3Dv5NdKtgNuweuWyJiG+vr3yOwXIJgt067WfVWz87iaFCMHadOz6OAHBmQgOfLz7w17Bbr3KCl5rJ4AJZAkqrBAaI+hwbpW4F1Ew8InAEkEMAkMEIawI5b5F0cDqfVabkQ+hN2Uw0UNBgQIBKxQEckwaOYbv5EXYg6Dc+R92VhFOmYIQBYUFyiEmiSjqEDCxH8VIqMICgRX1RsiOEJ66hrpYQ/DOOVldRz1QSFAOz4dTyLC6GQsnBPHOqsi+JscWovBwE+hQAUzo9wMu0ey6036XnxXAgWckuKFQ7W2JCTzXgjEj++EMH4RXfLqxpBMEOOsG9zt/hwrWKO8QQUkUhU1SXISt1nfgmgPh8okmvGLlugUtPQFlKa6V6F9w+XakdWj0aXzyjb7JxbvhJ/o8UmijsSZzfzepf2HltSuXBSybwjcXjHWZKY3jhRbqg/2WFm3aI6QaYkpbr3IaXnvTrfyOu6j1Fu/CK0/FqjUucPE3Zr775uteeeqYKzt+pwwvZXLoMa5tWKJFEoQPfabPYygssDbADV+0WCGcw7kERAg/YdSQiApwp9ixsB2eFhEu6Lm7hrim8nNXiJ94zo+Qc/3q5b4WicQ+YSUzSpIRz/V9PJwllj1cP87DCm/qGOn9xPHEmHDlTBg5eGCssaZ4H/G+x2oGKxPilLRo1/HRa2++vQX3L+/Yji1vabzz6y+d8jTeW/GQ/BH6hwA+68voY5zQkXeLO3dAmOmOD1lVT7/He4ON71icBcqy5JQKB+oR4fyhym0/RXcsitNQwWeoJYKfZV44o1CrwNDvKPgDm7WdMSHvSLdSnXr9GTr+c9/D22vHUj/e9wixeSfj798pO8Lrku3+ds/8yqUL52d048193QGrYxbYxOp2lXdMxWo1LqR+s96bzvvdd8Pazi0WiuRa0PXJKLmfGvzSpIvrX30dfQOWcvR70187NN5aWvhEef7ds+MWd3g9h/wW/nski1iq+VtwIQhjVBbhoCThvYyFRiRLorQ0UceIgAiIgAh4EJDCQreFCIiACGQMAVbkMGFG4Jspm8+APtNW/7CqEjccuJSYO/N9/Mof1maLjFH6BDZbTHZiuAuQKjX2uxrBt66fexB3fNVatS/mOwEBd3238xCXME5o9NmG9Wtq1Lnkclw0DbTA2JjChzfCCasQMPkJhJjsodhAePS9nQ9hEqt+vXwbI6x0E0OviacLjMr5/mvL6sZNn73QBVxEudKlXYtb43X9Et6m4IpKhByhgg7c9yCUYEOAQ0Ip5qxxEIQgGMIvMMe9YgkXAgi0ERwxcWeCh8CFslBIYAmE8gVBOa7L+BvrC1a6oehAMcJEGmUfCg8SVhWs6mSyyf080xKKDs7LCn+EMJyP76yide6omNSzappjR1taaAlFB8qMfawmtc/AZpNSJqFYsbBqkTodIrByeVPp0xiETrrdSlPXxGhCtkPcZoWx8fPrnGl9UmZfK1wevfhcP5Q8BzaE1pNmzA8oIns82Kb5Wz5BThHyIJC2zR7zE05EwUHq+NhTA+iPEOibvuPP78zlGwGu/dpWtmKVgJXRskXznQA2ZgxlK1YNHPs/W/LPOXEZgsVCeAH0V+48+Cb3O8ElDa5uzD4sNFjB75XPuYya+e50T4VG6DFVa9YJ9ONrli/hWfbdVi5ZON9ZWdzeun2naAoLLEUItE2BuLaK5l4Fl0/kXb18sWc9nIUFeXCXRX38KusU29vN8s/rfcNxCEMvaXBNgOWAPt06hSsWzIDw2La2qpn9WDY6xdOWjf73CSu0XSwm7lvclMV6ozghJYqRdp17PnVDsxatqQOLB8YMHdhv0JM9OocH4Y617LTmi1XhGbKqnlOF9kV+CoO0VilRj0NZzLPGGPXHOBer8H7kvUrfz7sDBbYEtwbB9YcrIjzr6XVDOAsvypv2auzPLX360UfnCsSu+nTebMZcvtulDRpd73auXPKpZ/9FDBtnudy+a2+swHMQh2j8iy8MYAGNX5yh9OKQieUwhmXMyhjVWVZl4ul1KhEQARHIvgSksMi+114tFwERyDgCTOBwX4PADyEq/vczfNVVxjUntpLdhG3j2tUr/HyVx1bS/lzHnXAC1imBzcu1iVvRtujjjxBgR9wuNF/mZPjIArJ6ZXTCqg1rVixr0rxVOxQgr4weOsgrb6Hg6jaEWn6rfIsFhV9fbt+25fKrr7+ZSeKwZ5/o4VUergTcJHK9WWOE5ylZpnxAOIZQrd/QsYHAt998uWP7UCuPyWqsq2KjMYqi8CK4YPhKT1anuVV6CPjZj9sfJsSsvncui7C2YB+/k1i9jLLAufBA+MGz4lb3O1c/KEZcvAZ3bo5x/qVRZDj3GOHNu9x+uN8SVhbvWBrDOSIIZ7CYIWGBgSuQWFe1RsOq/dmYAEqIHs8MGX3m2efk+dDcufkpK0CEchNlL4n+h6DK/N7wupubIWhCoD98wJM9I+HETVwp8ztOWfEGfqWuTtBdqlyFyihI/c5H4HDqQb/sZzmBIha3UeSbMX1qaCDeg5rgzrnokzkR+3EsNdw7hsDa0W4r+lusLHDFR//u5dbKlZH/3CLFELjzNy5MIpXNtURhQ7+7YvEC+ruDNqzvyMOPsQTDtfgVAQsLcxHvaTHDvrvueyjgCgol1JwZh7rWwi0g50RYiMJgwjtzA5YaFsPbV7FVKCQ21CyL8xGPcLFEUGFz9Y23BvzSc7+hKHmhX6+u0ZQ90a6b9mc4ARYPELsJiy2/wON+lXDWv9sswyGuNTO85gl8grIVqpzPc4DVUUZX09YGBfoM+hcUorGeD0ti8v5g8ZWcBbPfsfUb3dDU7fNbEJP/3MJYvAY2LK0mjRnxwmvjRg7FOjnWOiVJPudqDesi+mkUF9pEQAREQAQygYAUFpkAWacQARHIlgRwYYNrGVzlsBo8ZVcVu6uLWwi+swI4Pa746WechT/9HCg/EMSEl+kELusiuNHgGCw/3CrWWe96m8FbSIr9AThNaFfp/Fq1iV3hp4xw8SYimeEXKb5fCIWLmOtvbd6KFb5+AkRXHpNIr4DZ+QsVwed0YMPVxviRLwx4743JExNkBatbXek+w12cUe1oK/Ej3S7RVvkfsroz6PKDeBy4hkLAgpXHP1FWkvKc4tecZ/YQC5z0uJ9VRvYj0Lztg50vtBgOWHb17HTf3WkhYG7GA/2peZhC+R1xK1G2XEWsNLCKiBS82quQc4sUL+mCL6P4IHaFl3UFbkUaNLrxFspYPH/ebGJteJVXqVrNC4nPwL4Pg/7Nw/PxzkARgXIkmluTyxpeewNKW5QkH896HyVkxI3+FndVVWpceNG1TW5r0adzh9Z+B1h3HYhfgcBxzozIyhACW5MXVyxeFhFOkU6eNydPGIP7qkgVddZ9BDn3yodFn3MJONCsK8Lz4DP+jjYdHuZ3FEx2m2CxloPA4X5BwdnvFCV8f3dq7PGmUGw5QSXv5emTx48Z/+LgAV73SrRrpP2ZToB5P1ZKvOe45+N1G4cbRd6VBSxVsMQCimjv6ExvZGaf8Njjjjue5wmL13j73bTU1Y1nA9bFcSgH8lq8IM63Ye0qXHr6bli9uUU8KM792nT2OfmwgM2xecPa1TfVq1UhneJUpAVJRh/Dc0PMFqzwWIxDHDBtIiACIiACmUDAb2ViJpxapxABERCBlCbAKnB8/TPQxQ1Nym8uCKB5NMH1z2Fvzq2GxZllJf1BG0ITC18RmCzhliLSyRo2vrkZ+1EGIGDzyusmgAijUFRMjODDvHCxEgH/wZEmfS7gNsIoAqq+OOjpg9zEhNbBuZjyK48Ai+Rn5drNV9SqiE/gzFZWHPbFzKQCgv6GncsqzopQBtcX0Tae04ssNbCEX/fQMqIdq/0icAgB4szc80DnHqyCfbjNHTfFI1gKLQzf4Px9bEiQVT/cLg5DNJdJXsc76wW3b+Qg70DaF1xcrwGuqsg394N3pvvVpe4VV+JiLQdxKQgW7pXP5F0ITnN8bf6ivJTSoce4fnzuB+9OjzWQ86SXhj9PGfWuanwTsRX86orQn30I3rxcBoYed2nD/a5SsJjxKq+0uW/id5Qfo1945slIjwZ1Ig4Rebys6/i98a133hMIom4WGOG+5FEs9Xx26BiUSKyCHjPsuaddW3Zs37rFL24G5TpFCdxxnxWpnqH7TjEllLMIbFjzvMK9H2nfSsqKWOlleT7m/SjciBuDS8d4Y4wQ+wprYSwfD8RRyPJWZXEFzqtYtToWZWlxwxdv1VFI5y+437Jhlk9cIL8ynUJ6x+dbAvHh/LZmLe970O3zi0/E/v+dckpgbLX7l19+TmFlBU3k3YGrUe573I6itNAmAiIgAiKQCQSksMgEyDqFCIhAtiNA34o7HPzis5rtSkspLwD96Ydd33OlbdFsICD14W7OjZNXwD98vDNx4xyRBIH/PfbY4665qVlz8k1+edQwr0kVq4BRKpCHIN6Tx48aFmmVXGwWFvuDmVIeVhGfzp1FQGPP7YACZM1Kz1VvtmI2MCn8ySSXh8s0mxyPNROBpT+1xGpQVqiHBp0+CIMpOXheUVagGHLBwLMJKjUzIwiwOrXXgOFjETT3e6zT/ZGClkY7/49mekUe4vhEy1sgaI213lzbRcsbvr9shcrV3G8Lzb+5nwulBtftD7aNMNwv7gTtxrKEfF4ujNx5zBgg0O9GU+acV6lqdRe3Z+LoYZ6u+rzaO9vcJ6HwIY6IO94rnxnYBSws/AKZu2OITVTNXEyhhHp/+uuTvMpyLq6W2urnaEHEC5grKif89+KNQgLLEs7D+yv8fG07detN4GzciBHLiHo55fvOr77E7Y/vVrTE/pgdn8ye8W48Lhzd+4hj9U6K9ynL8vy4XUTwyoIaYsrgjz+eDUGts/jkneoXpyieMpM+b0WzJqMRmaGwKGTmwE75Sv8WDzwbNxODJOASyu+4qrXqXIwrPbd/dYR4QcfYAJt8Xi5b46lXEuSFG4pl4r8wpmR8qU0EREAERCATCEhhkQmQdQoREIFsRwCBKf0rE0KEpe7vlAZhluMEZA64YDot6M4prQ2mDBeM9Z2pkw7xKf5fs8GnbPyIR1qZ2/iW5vcgrEJR8dq4UUO96uNWmrryJowcPNCv3ig33OriTevWBALphm8oUohL4X4fN/y5/pE4OAsLvwDeByaFe/YejmultF6KZDzOKQe3W+VRnuGqLJLCkOcTc38EfDMscV1T3oVbMl7YZKgzyooh49+YgbIUq6h4BOxe7TOXUAEXZbnz5i8Qrf3OVc/m9WsPsUqLdmyohcWr40YO8cqfy6znnDAL4Zyfy6Hipc+r4OI4fGQWEX7nhhH7dv/ys6dbKXfcnW0eeITvWEAsnj93drS2uP0I8Fcu3R/wuljJ/VYUXptzf7J1k7cliDvmxtvuboNbqlnvTZ+68+svD1mdjqKmZNn9MYf8YnuEnt+9e4hJ5BVDguDWBLblPcc5Q4+94prrm9zSom0HfsPdFe5o+O7uAa/6ueOpp1NsxCv0dLE+cOMF31ivhfIlDAHehQhfL7UUry9+FuE4ywremXItbRBwO8fVXbJg3pyMvsrOlRt9Ff1GPOdzz+7ff//jGaMLS61OPfoSY+zAFikmh3VLgXL+tb4gnnokYV7cMaI4RmGHdUqgvT5x35KweaqyCIiACCQuASksEvfaqGYiIALJSwBhJzEsEDCvspQtVsazUhO/2ZjG33DbXb7+wqNdVoQpj/Tu/wL51q1aviTSCi/OxSpUrzJRVDjf3lMnjHnRKz4Ex7FC1R2P8ObrHV/gp9lzK1SsRCl2/GaO2/2EdYWKFitJvci3y6SN77/pvRKX/dSdgLp89wuQmo0mhdFujVj3I4SpYgnTfQKDY+0UzcIJU/8LLDW2hJ/naPljrYvyZSMCrK4fPumtWSg1EVj36eIfNyFWLK6fIcaE61f8jnV9SbSAquHHn2CdZUEz9eJ3FMBzP3zvLa9zVK15YV2UFuyLFOy1bjDYNq6bYgn+7ZSyXudk9XKtupfVZ9+IAX17xcrN5XOriU846STeyYdsZ5yV+xynhI5k6YF1xU23390Wy5JRPq6eYIj1Hyf5eNaMqHE2nPARRYxX3SpUrUGflGPT+jWrnGsw/sZdYrd+z7/I96kTx7z4xqRxo9zxeYJ+6p3Fo1e5ufPkK+BcOM6fHbs7KMrS+yjeOzCh8jM2JR4YSjyssHg/xrOhoMCVFBvKqmzvGsdZbxHrIdLYMR7IkfKaMjhgDbZ88YKP4y3Txdw58+zcebyOve2edh0LFC5aPFTZ6beQhuO/2/k11gY5UKrGW5cky/+r1Zf+3Fkues45kqxNqq4IiIAIJAUBKSyS4jKpkiIgAklIAGVFTUuVLCEwTfUVSDkQTk19ZWwgGN0drdp3chYS8V67ezo88pgT1Dzd45HACtLwDeGNc+8Uas0Qmq9Dtz79TWdxCsqFwf17d/OrR6HiJQ/4Yp5sK6Ij1dcUFoG85h58s295FiTV7Zv2yrhRkXz7Mjl05v1fbPvMs8xsNCmM91bxy4+ygdXPuLhBeYECKtLzR34moAg0cZehTQTiJtDo5tvuGj7p7VkIsBD4P9z6jptYGR93QWEHmPAo4NqH1bGhgZK9ynWWbdYVI2A5sFWufkGdpne1vt+vLvS3KIrZT0BrXAx55a110X7FAUL7D9+e5hnDgf0uSPRys8KI1P9ZWKFAfCeE7O78oefFXVKXPs8GrD1Y6UsgcK964TLqzrYPPOIVpyJ/0E3W9zu/CQQvD99cvCF+d8oYr3wPdHviGazn3ps2eaKf66hS5SpU5liUTNHcQZHPWTls/Wy/dUT4Zh6jSvLbxrWrV7h9WIMMGPnKNNigDCKGhNtH+3nn8Xckt4ZO6PnFti2bUap7ndvvt+92fhMQUnIup5yJ53jlzVICvA9RUmDRxHWP15KQ9+oISwSIZ7yS7RX7tSymD4rkSG4/0/OKFy1VJmAptmXT+rXxlutcBdaoc8nl4Qt9UAy3bP9wd8qcN/P9t/nEgurnn34kbonn5hTjeQsUKuzVd2KNVr/RDU2fe+m1t1C4x1vfBMrPc4Iimr4VqxZZliXQxVFVREAEUpuAFBapfX3VOhEQgawjwIQQ4Sd+8XEPFFhxn+rbwD5dOyEEYQL33OhJ03FbEU+bb2/dvtNd9z30KMewatTPxB4h2NoVyxaTr+4VVwWCu4Zu9a667qYrGze5jd+e7PrgvZF89joLC8zrF8ydhUsg3825b9ppS+n8MrnyEOq9bqtfI5e3XwFiOpWf3eq38PxuUmjzvQOWIKF5zDvW8Xfd27HLMy9OmIpJfzy8UzQvripwdxFwN2Pbxhja+aHlYQXd7GBKeQVjDEyUJQYCKAn6DR372qNPDhyGUuGdqa+Ob9/85mvSy683fRdKV6oSKQ4D+3PlyhVw8eKCq/K9Wq06l7zw8uvv3d+5V18/AXOl82vVdk2d8dbUV/2azcp+9hHg2SlSw/NybieIX2lKhkgI169evnTfvr17iSFUvkr1WuF5O/Z4aiBKXRQo3Tq0usOvrC5PDBjapmPXx5s2P1gpc+EllzesYOWiOFr4yZyZXse7QOXsczFAwvOx8hirEawW+j32cHu/erjrs2zhJ3NjuHUOBL7esW2rZxDck4Pxi1wcE3M3VclZ8LCiu8NdTRrBz53rmGOOCVi/sPkpndhX7DCEnj+YgsO5YTSXVp7vJFxZ9Rs2bvIlDa7BYk1b4hDgnYj7IiwQGSvEq1DFOoN7DKUHruqyvRzh2ia3t+Dy0tcxFkMR4KV8TY9bgHKLmcKSsiJZHvudC0U68WqIrdapV79BbrzIGHrg6Feno4RECeriDnG+SG3hPYBVCdZaNzT7f6tqFBXEMJr47rxlxHJCQXL8iScm82IQ5nFYQrOwhXmH3LOmxw2tMkRABEQgBgLyPRkDJGURAREQgTQQONOOwd8vK9AKZJeJHYKMu66vX2egKStYCfr4wBHjrrrhljvGDR/U/5M5H77n5/O6WKmy5dp36dXPWWUQpPaJLh3aROJObAv8rjdred+DCz+e/aELbHtRvYbXPNZ/cMBFBu4y3nx1/Et+5TAZK2BRDNk/Zfzo4fjljnROF3A7krsNt5Js0cdzZqK8OdzyPnhr6mv3PdLjycrmJ7lM+UpVVy1bTDDpHPh/hy3KCgR+uDPJeXTOoyOtaE7DfZyMh7ASLuBT2jZWhO6O0ghWzzEBZRUzk1LcG2yzFO/q02RkpTqngQCCcFt8+leN2pfUu7bJbS1Yec9z90LfXo/6uQtKw2kOHMJqfYTVJK/gyy7jD7u++xYFCn3gmKED+yE06jNo5HgEU9TLKT7C61K+yvlYAwYUp3NmvPOmV10p49yi+1fJRopLcfY5efMhsCLf1s2RY0KgpP3IzofArHOfZwa3vOmqS1CEcDwKCISBKH57PdyuZaSyFs6b8yHK5FYPdO6BxQD9M1YlTe5s1Y56THtt/Et+/t6Ll94fcJut/rU33jJm2MCnnWsXruvd7R7qimtB3g3dH2h1xy4zMfC7liXLVsCiMsea5UsXRbveWOK4OB+//77bs49ycS1QOjVp3qpdy/aPdEchRPta39Lo8nDrCHhSv1NPP/OsWhdf3mD65IljuabhdSlWar9bmdXLliyMVs/w/XCY+c60KbBCkdN+yc3XuPemxfGu0KJdp661L61/1X4O8Zcfb32UPy4C+yw3Fr8oNlE+kOLZUFSwsv87S7iVilfhEc+5Ej4vll3lK+/vO7v1HTSC5CrNWHefaRP3/3/v/k/7duC7/XbQfvbZhv0afS3KZeIEDezTrZMr85x8Bc7ld57ztDy7jBFfHTtyCH0JFoEX17/6un179+yhv+AcWC53adfiVnc+Fh7hMs8vHg5986vjXhxyb6fufdp17vkU70Usu4hhhFKEcjjn44/cf8/KJftjCSXphnLPBdqWO6gkvYiqtgiIQHISkMIiOa+bai0CIpD4BBASIADNZ4mVndlG+Mnk5vZGl9ZEcHHznffcR0BCEoKT9atXLEP45gQxp5sz3VImhGMVrbukuP3o8WCb5sTDiHSZcT/VtEXb9ufkzV9wxKS3Z8//aOb7x9pKL1bUchwrnXt2uu/uSGUg3GNVHOd67eXI7qAox8WwsPjivooI56JqrClpot2mhYPuqCKVRzBzlD0Eux32ylszF33y0Sybz+ZEeeFWUn+2cd2ah9vceXOkAOTR6pIi+1EQHhtsC88glhPRhCpOqYhlBpNSjss2z2uKXPdMawbudJ41lzyhJ0QYQ7wK+reMqAjKWJQVof2k13k+nTv7AwTJCI8QIrmYF++/OWXSoCcfCwSuDt9YEeyCP0+dOHak38p8lBXOjci8me8FXIZ4bSbjP7DK/+sd233jAbljhz77ZI8LTNCFonfyzIVrcK2C8oG2YhnxVLeH7pv+2oQxkbi+NGRAX6z5sEjo+czQgxTUsOvX/aGA4sJrKxb0Cb9u1YqlCNwnvDNv6SezP3iXvFVqXHARwjwE8j0fureFnzKHvLAuWqJUWb5j/RDtPgh1ZWiGMZ7BjwkwjmUHyn9cUlEmQsVWTa+5zAXZDj/Pyy8OHsC1533x9PCXp9x9Y8O64XmchcWnpuiPVk+v/QgprzBXLyjEXv1gwaotG9evxfWWsy5EODt68LNPcV3SUr6OSX8Cy774BSViAUsoKXDFhkVhvK5tyE9gaSyGiWWBAiTbbigPUEzw7OMSlQUwR+W0/2yAhrXCfhd1B7rDuDn9Hubaz1lXvGkK2LQuTBn01GOd859buChu+1CaukotNauwxx5ofaez6EVpe3aevPlxS+ensOBYFOMly5SriPLDuXLldywDJ9uYetzw55+J5J4ubihZd8AaOzVuQ7Fo0/gw666DziwCIpDNCEhhkc0uuJorAiKQKQQQgDKoRfC5wRI+T7PVxuTt2ccf7TjppeEvsJKrfqMbmxK0FNcjoe5HHBQEQotNEI+QA8VDLLBQMrS7/YYrEcog/HF+01l9OvTZJ3pMHDX0uWjlsEKM1WpP93i4fWhQU6/jWPV7pM1A2bfChGB+ZSPww52V8wMcqQ7OJN9Zh/jl7W7uUIZMeGMGQj0XgJa8+DEeO2xQfyawftYr0Rik4H5cD/D88YkCIqLVTPm8J/5jwhxc7iy3hO/+gI92bSLgRcA8avxJ30OfhWUXfVysfVZaib5msXWua3r73auD1lV+5Qzq26NLKQv8jWsjhGi4/5hg/eDAJ7oHLAS8jitftXot4iGgRB7tE0ya4yw0QiCwKgKtdauW48Pec/vC9tMX/WQdKsGio7WZoK6d772rKauTCf6N4Itjtm7asO6Jrg+2XTgvulCdmBEmxK9HGVjrueMnjx817JXRw5/3E+5xPos/fS75u7VveVtfc+2FMO/yqxvf7OpNex8zBTqT4NlOAAAgAElEQVTKg0htOc0UG86PeyQXhK4MrCPghFDTwpR4jhGmvDx6GEoALFD+sqXZuHQZ0r9Pdz8BYq9xi44Y0v22p1HiX3PjrXe6hQGh9SZALpYdBPomLki06+O1H7cxz/Ts/EC7Lr368k5yVoXcb+9ajI+Rg57uE0sMj7ScW8ccFgFWiqOkYhHNLkuMVeMVvm6xY3AtxbvygDuyw6pVkh6MYvP8omcd98+///wTPv5CuYvy9hgzhcVVoP07lr/pa+3fMfb9mJz2xR5/U3HkzIl2I0cwjhBjSGLF8JyFotm+9bNNWNgNerK7p/I5Foy8u9o2u64+inczLi5lhh57Nq5dtSL8eR3Sv3f38y+se+ni+fMi9nu0+8GWtzbGHR59L+1mAQ3WISk0JkVBR8wXXMFuTcMzE8ulUR4REAEREAEPAtk+WJbuChEQARFIbwIm/KRvxedpn+CEcIJ9vmWC0XhXs6V31bK0PFZrlSxTvqLJdXKfcOLJJx9hCoBff/npJ9wmITiJFNwvUsURzJWrVK2GyWDyffftzq9XLvl0fjTrjLSCQOmCqTv+itMjoC4WEgTS3WhCOy/XHaH1RLBVtWbti/PkK3guPgbwYYywL61tScXj7NmjWYUsPWjpAksPWHrP0t/2/Pk22Y7D1Q2rDQlWzEq6gFVGpGNSkZ/aFBsBFI1/mzQGhWdsRxx+LvyE+8W5CS0dxeqZuc/Ji2DM5PhfRIplwHEEvL717rYd3nn91fEImfxqyurhOpc1uBphVDRhNCttv7eI2gjYYm05lm4cx6pf3gn0b2nhy/EoZ6L1p9QLt1HDXpk+EzdKF1cocjb9cb2rG99kOozCvI/MpdGihR/P+TCaq0DXRlxx2WG7ln768UextJtYH0fbhcIXfLT8pow4KEuXpoH43oENRYV9kFxMgX/eHP3kMQ1ve8itBmbfP3bMPyhVOvd+ZjDWD1zLaOeNtD+3aXsqVKtxAYqfr77Yvg2ljp/bscM5j449fAL2jmOxBe6LnNXvn/Z++z7WkoPvVpcdAS4K0ED/p/dkrBSVL9kIBO97xofVLeEOEIUfyjrd98l2MVVfERCBpCQghUVSXjZVWgREIJEJBAe4p1gdCR6d2xKKi5Ws5E7keqtuIpDsBILPHj4YEMoQEBa3FwE/3VEUFriDwiIDH92sPNVkNNlvBtU/UwgEheUHncsE45mmyDmcRt7Som2H9o8+3g9XT+3uuOHKwykro4/1U1iEKCsQIiOURtlK4hqgwGBVPfv4jf4tR7Jcn4xmmp3Kt3cj9wAxmnBbhkXPRnsn4tZJmwiIgA+B4JgSKzyeG1wc4uo3MJeTok63jQiIgAhkPAG5hMp4xjqDCIhA9iTAgNYF5/xNyorseROo1VlCAL/aCGQQzgUEdNE2ez5328SUvNHiXUQrSvtFIFsQCArQ3cKnA65lkkkYXqJMuQpcrGQIDh1qUeFusKCygiCwJCw46b/4dIsjUFoErCssOYXGXxyXTNcpWzxQGd9IFFdFg/fHmfaJC0RtIiAC0Qng3hdrwR2ub5WyIjo05RABERCB9CAghUV6UFQZIiACInAoAQQIX1tab+k7ARIBEcg0Ak7pgM/hmFd6Z3eXbZl2dXSipCcQoqw46PlKNiF48VJly3Mx1qxYEtUlU4JeNCwoGGvwiaI23O0k14ffUVow53MWF3/bNcRFVMz9Y4K2X9WKnQDXf5slFFe/2vtuT+yHKqcIZGsCKCxY0KJnJlvfBmq8CIhAVhCQwiIrqOucIiAC2YEAbmnwc8qKHPziaxMBEcgcAk4Ix6piuWHLHOaHfZYQ10KeQlSvFeaHfVIVkCYCwWsRep2STvBNINz8FpwcALHEkEgTqAw8yJ4Xp3zIZaf5za5JpBhZ/1p+FLkIq48N9ot/2m9/2XGyKsvA65RARaO42maJz2wdLDuBromqkuAEgpYUf5kFrsaSCX6tVD0REIHUJOCCs6Vm69QqERABEcg6Arvt1Pg7/cwGvBIIxHAdLMDqEWEpRybGtI2hhsqSRAR45g4IZWS+nzRXLukE30lDVhU9iEDRkmXOI0D5js+3fkaA7WTCE1RWMIc7zhLWE1EF0ATctnwoNRBYo7hA0fEfrxgkycRCdY2ZANf9d3sXEmxbwteYsSmjCATiVfwTTIpdoRtCBERABDKRgCwsMhG2TiUCIpCtCKCw2GxJ1hXBy+6jfEDY4vygkxNBChuCSybVfEqIma0enbQ3NkQxoXsm7Rgz7MjwwMEhJ5JP/QyjroK9CJQoHYxfkZzuoHhnOgsLBNGxLoogH25NXDwLyjgQf0R3SuoSkJIida+tWiYCIiACIiACqUpAFhapemXVLhEQgawmgBABv6exChKyur5ZcX6nrHDCE/c3ny6QqLO6yIr66ZwiIAIiIAIpSKB46WD8iuVLkyp+RdAignckFhLHWGKsEdMWjFnhxiQsWuP4nEGLjZjKUCYREAEREAEREAEREAERyAwCsrDIDMo6hwiIQLYiEFzlLZP7yFfdWVWgrMgZFL7g1oK4H27VJ8IUvvO7GWj86ywuDir5iCNCDTSy1a2mxopAKhDQCu9UuIpJ1oaSZctXosqrly9ZmGRV53nhnUksCmJlxbX4DNdQpqDgncqiAN6xuImKFP8iyfCouiIgAiIgAiIgAiIgAqlAQAqLVLiKaoMIiIAIJBeBUEsK3kPHW3KrPRG+OIUFygz3HWUF352rqORqsWorAiKQwydwttx36d7IVAJH5zrmmEJFS5T6+6+//lq7avmSTD354Z/MPS8oGZxrqHiVfn8G36Ucx7tVWv/Dvy4qQQREQAREQAREQAREIB0JSGGRjjBVlAiIgAiIQNwEEJRgVYEQ5kRLrBplw23F6ZZ2WWI1KUIV56ubT8W2iBu1DhABEUgPAnuaHyjlgKA31wjF2kkPtplRRoky51U48qijjlq/esWyPX/+wfsn2TYXQPv3YMXjUvrhGipoZcEiAFmDJtvVV31FQAREQAREQAREIBsQkMIiG1xkNVEEREAEEpQAQhZcUyD0Q1lxqqUTLP1i6WtLuKw4ObiPJuy0hICGROBQtrgENQnKQdUSARFIPgL0W1iB0QcdYUoMhL9OmXpIa0yhoS1BCJQpX6kqVVm9bPGnCVKleKvBPYdSP/RdGFcZQddQHBOwajQFxr5gjItAOfZ34NPHKiqucymzCIiACIiACIiACIiACMRLIC6/p/EWrvwiIAIiIAIiEIGAE/idZHnOssQnCoszLSH4Q5mBuygUF/+zRJBREn/z6dxFCXKMBCwOiAtifuAzxkOVTQRE4FACKCzoj1C40n9hISb3Ogl+p5QpX7kaVUzC+BWOLMoKXELxjkxz/AmUFna8lP4Jfr+qeiIgAiIgAiIgAiKQHQlIYZEdr7raLAIiIAJZS8AJSBDsIeBD0IfQBaFfUUv5LaG4YEMYiFDwXEtlLeEm6hRLKDAC+4JC+KxtUQKc3TgQmZyEMsJ9/499h1EgWTWxrMTFFp8kftdYIAGuX3atgq3kPsKt5k5CBjw7Z1sqYqlA8JN+TFsCEyhXuVoNqrdy6aIFCVxNz6oFrSCcS8T0cGeF0gIFiDYREAEREAEREAEREAERSBgCElIkzKVQRURABEQgWxFwgbcJ/ulcQuH+iYQ7KH5HoO4sL4BT0BJKC37D8gLBe7Z/jzklRZCFC1qOcgI+WKIcE/wMtUhh/3HBPEdZGaRQRYdTeGSrm1KNzVwCKCsy94zpejaneEXpyjOWJ5hQYPB8aUtAAmfnyZv/jLNyn/PD9999u3XzhnUJWMVYquRcQh12LKcQBUgs51UeERABERABERABERABEcgUAophkSmYdRIREAEREIEwAggqWdmJSwviUZxjCUEfrqAQpDt3UeRhFSmKDH7/wRIxLhDUnGHpG0vOJUZKu7ZAMeGxOcUPu1wGFBMIUPkbK5T/BlnzN6zxe45AlTzs4/fdwWvBSluttvUird/SnUCoz/x0LzxzCqS/+tXST5Z47niWTgv2S66fSul+KXMwp99Zylc+vyalLf3044/Sr9TMLSkYNDs9+2ndo5l7CXU2ERABERABERABERCBKASksNAtIgIiIAIikBUEUEQgbEfIx/ctlnIHhX0oIlBQ4BoKX+MIBFFmkJ/A27iNYnNCdoSG+4IC/UMEL0cckcyLuCNeGtcwZ02BAAsWKCJgB1c2XG6h6EFZ4VxswZqV4fD/zRLHUp4LZp6ewrCIjdBOEUhiAihLsQbDuqJAyDOFAvZ9S/RdPEsSCCfIRa5QtcYFVGXJgnlzEqRKh1MN7q3DtjL0Uhwq2PbhXBYdKwIiIAIiIAIiIAIicLgEDnuQe7gV0PEiIAIiIALZlgDuilyQWgR7qyz9HBTA4PYJF1DsL2QJoTtCP+fmaLt9R1iD4t0J27MLSKfogQUWEighiOtBnA8UFfjTh1loQqkBv1MtIUwlL8dhbUE8EBRCxAfBioW8KavlyS43idqZaQTos+iHGFPnCz6TVe3z4uDzhgJRz1OmXY7IJ6pQpXotciyeP292glQpTdUIUTI4xXSaytFBIiACIiACIiACIiACIpCIBGRhkYhXRXUSAREQgdQn4ITugcDPlhCa84k7FVYtnxkU8qGMQOCHZcWPlrCq2GqpWDAvFgHfWcKygOOce6hUJQg3JxyFF8HJ+Q2FRV5LKH7g9IUllA9YqxAEGAUQ3+H0pSUUFXxHieGuAd9hjZsuuYZK1TtI7UpvAvRB6y3hFopnjmeIZ/MSSwiT3ws+o7KySG/yaShvwdxZM96fPmXS5g1rV6fh8IQ6JAVcqiUUT1VGBERABERABERABEQgcQhoxVfiXAvVRAREQARSmkBYDAbePwj22AigjYsitlKWEK6vsITyorwlLDFwu4KbKITpKC2wBuC3jy0tsYRbI3zG89tB7oyS3SVUkJtT8PDpgvzCAg4oK1A+wBFmCElXWkJoWs8Syh2UFCiF+FxqaVeQFUoMhKzfBrlyTeCI8JXYIf8kOz9rgzYRSFcCe5ofUhzPDQrD+sHnEIslrJ9QpqKwoI9yMS0OOjjXiHStmgoTAREQAREQAREQAREQAREQgaQnIJdQSX8J1QAREAERSFoCziLCCdtZ9b/A0veWvraEcH2zJfI5ywIE9AjqF1paawm3RrhhQeiOgBBrgVRTxvOuxv2TayMKHJQPKChQzuAuC4UN1hXsgwH7WNGNMoPkFB742mdFOEyxzqBcApcjTOU4eHIs5XDeVGNpTdImAulOgD6JfmyHpQ3B5xLFYWFLKAx5BnnWtImACIiACIiACIiACIiACIiACEQhIJdQukVEQAREQASyggDCdAR6vIewGEAYj3CPjdgLKCZYtcxKZQTs2yxhWYFFwKLgMcRhQKmBgB0BPgoPBO0I8ZPONZSHBUqo2yzaBSMYoJxAscDftJ24FAhDawS/o+zhWKwo4IOlBC6iYAJ3rFlKW0KwSiwQNudmivI5FusMfuMayZVNEJI+RAACWEWEWVnwjPCs8bygFMTdUBlLWC652DtOAXjQ8+TKkaWF7i0REAEREAEREAEREAEREAER2E9ACgvdCSIgAiIgAllFAMEdygXcOCFkZ8U/LqEICo0wntgLKCzWWcJNFC6hENDXtsSKZawCWNmMIBAB+w/Bv1FwUG4yCtpDLRqcFaQLKk4bsSJBmYNVBXxghSKCQNuVLDnXNCh9nPUE+8mHsgdrFPztf2aJIOcEB0bRQ9wLFB/kRSFCPeC4zxQpfP9XrqGMgjYRCBIIUzD8a4oHLCxwpUZfRV/0ZvA54rllH7/zrOEmKhn7Jl17ERABEfg/9t4EyLL0qu/87vbey732qq7q7qquVi9Sq7UiqRvtEkhCEtgCGxBmGWOz2AFBxIQnPDZM2EM4GGxwmFmMgzHG8lhsYgw2MGaTECAhCdDWAi3dLXVXd/Va3bVmZb7tLvP/3bqneZ3KrMqqyuVl5rkRJ+/L++679/v+3/Le/f+/c44j4Ag4Ao6AI+AIOAKOwIYg4ILFhsDsN3EEHAFHwBFYBgFWI7MhOrAhSDwiOyaDUIecx3MCEv0zsnc255KAGxKd9/E8sFBQnAc5CNGPPS+XxRZqAcrO9zN1q8UCGWIO9SRO/tEGK4QFxAtIUOqOEAGWiBL8j6hDgnLOM9HCknRzfc7jWpCseFrg6cK9CS2FWMH9FyRUOLm6hTqPF3VTEWCsERYKAfF2GeOMcck4Yzyx/YkMryffHAFHwBFwBBwBR8ARcAQcAUfAEXAElkHABQvvFo6AI+AIOAKbjQAkO3kUIMwhxyHZSR6NBwAEPSQ7G7kteJ9E2/c075HLghBHiB2sYjayH8LdyP7Nrt9q729CC8IEnhJ4meBJAbmJcINHBeFm8DphBTfeJq+XIcyAzS0yvFGOyRAoPikDBz6HAIQXBV4phIoCm1fI+B2ASHS+uS74QrjyecqRyMOiDgvlHhZCwbd1ReBfvJ9ob/XGWCDsmYV2sxByK4pnP/adr1rXsq3y4jYWGVMvkr1Sxvxl+WUIuUZenocYU6u8pp/mCDgCjoAj4Ag4Ao6AI+AIOAKOwI5CwAWLHdXcXllHwBFwBDYPgRUI77IhxPESwCDdIesJZ0RYI1YlQ9C/uzkGef5NMoh8CHVWLhNS6k4ZeRo+K0P44NhY5bFYkqPCGsJCQFnOCL6XESqoP4QtYgXkLd4QiBXszfOE/8HnQzJwYUU3Qg8bGEKevrk5n88RFgpvCoQdvC8IUYNQhGBk+TG4L5/DOI/yWO6L5tK+cwTWBwFEB4kWluvBvIwYB4wT+qMlt7Y+uj4Fub6rUk6EQ8amjWHGGmMSoZE5jrnKPMuu727+aUfAEWDeMBRGwyo+JwqOiaDpLeUIOAKOgCPgCDgCjoAjsEoEXLBYJVB+miPgCDgCjsC6IWCJnVl9jNCA4ADxDuEHyYeXgHkU8L+FLoLMxwMDzwGOQ9ibBwHXGvc8FqNiBeU3YhY8yCeBKAOx+TKZhYFCmOE4G+LDEzILAwXRe5/sz2QvlSH4gCcbCYE/1eDE/2BnK78RinjNdTifPWVgv1XDajXV9t1WQ0DEYiny0XKoMC4gHfmfcY+gRr9ERKNvWl8dJ28FyoJHBbkqmLcQBy0PDeOYsYVnGMLGOJV7q3UVL+8OQmBEkFiu1vZdyh5jAYDlyOJ/+42xgxDzqjoCjoAj4Ag4Ao6AI7C1EXDBYmu3n5feEXAEHIHtgADEAgQkYgMEPJ4ACBZ4EkD6QUpy/KAM0h0S/60NIQERT0gowkiRuJtrGMk+utJy3HCibJYsHKGCkFaQsxynni+QIVqQowKSE7KWVdrsOR9Pkt+XQXpyLp8nLBR4gBfJtNm4FveB6AUjsEMIstXrhILiNeGlHmw+A+4c53NOqDag+G7jEJBoUYmgtATwlgSefko/NqLfQqhZHx2nvkoZCQv1ERmh1xBTEVcJx2Zjz3LPbBywfidHYPshYCKFfV8hVvAdxnzAOGQbaD6pc2Yxt2w/CLxGjoAj4Ag4Ao6AI+AIbD8EXLDYfm3qNXIEHAFHYKshYMQCxCTJnwlPRM6GYzJW/EPy8RqvCQj4A82eekJC4C2AUPEF2SmZhY/h/XHNY0G5+A5GgMBjgvpa3H7qhPhAXSFeTHSAAIWwPS5j5fYJmYV6+kO9Roi4Q4aAgfjxBzLEG64NiQO+4MR7iDxcg/e5Jt4a4Mu9KQcbr31lagPGuO/6f7/u62yMJ2tD805Y+n/dru2fHx9BapkV1EuJRcpMf6Uvm4fFuPZP87JgTuI145LxRV4eNnLPfFxGSDYnUMd9cHn5xhWBUbHCBEwEfQuJaOV+zlMQ4cJFi3FtTi+XI+AIOAKOgCPgCDgCf42ACxbeGxwBR8ARcATGBQFISMgGiHUIe0iH+2UIFKxQJrQK72F4ClhII8p/TPZ0cw6iByFZbBunsEajISsQChAT8G7gOIID4gxJsu9ujj+gPaTmS2R4kJCvArEB0eJNDQZc44Uysg4j2EDoGmGDVwX1x1OD6yKQ8JprcN7nZXhWgDEGdqxKtRA2JNt2QlWAbPYmQWLpRp+hnTHGDv2HsUH70c4WPg1Sn7albyFMMW44r9A1WeXP+aPC3rLtLXFjXbcVYsw/5z0hotFCvFCO0TKORf8EnyVtRLkQXPF6Yh7DQ+qPZYxXQraR3J7xOk7z07q2sV/cEVhDBMxL0eYu5jm+0/gNwcZCBhPgLS8Oew91uIaN4JdyBBwBR8ARcAQcAUdgvRBwwWK9kPXrOgKOgCPgCKwKgSYZt3JSVxaTHoKepLWsSIZYJUQUxAPEKv+zahmSAuKP4xD/eGVAxEMSQhBaDOtc19UtxoJ0t9ja4ML3L94TkMeQKIR/QkTAXixDgCB3xwkZxCYrtBEpyNdhibgJl4XYQZ2/Voag82XZb8veJXuD7JUyCByucax5H2zx1niRDEwpA4Q35bNQGlzTPCz00reNQGAZUcJuOxqjHWGCdkKAQsii73xShijBa4S7e5r2JVcC/YTE9YT5QrCgbyGE4bmD8Md4spwv9C1I9rHzXGhWRY+FOLHKvmCCBZ5Mn5G9TXavjPFG2zGe/0qGaOSbI+AIXD0C5qlo3hXsTcBljPEdyvhivuR3Av/n7mVx9UD7JxwBR8ARcAQcAUfAEdhoBFyw2GjE/X6OgCPgCDgCl0PAhAlCFyFOkMsCIeNzMrwsINgtjj0rJS0cFOQrK5jxzIC04PttLJJuSzChvkY4I6SwGSEMuUJIKMhmwjtBrkAiQ6xAbCJgkDybuiLQfJ2MfBUQzxAyCBLUE48SW12Kp8VtzXU/rD33YHX9XU05Pq09K765PkQO7+FZYSvYXawQGBu9rSBWGCFnhBv9mrZFtECg+6Zmf0x7RLsfbPZW/O/WC1bxk4gdrwtELMSpj8kQNhC8ELPoXxDrHEf0YgwhjpmQEal89IsVBYP19sDY6PZYo/sxzhnLbODOfIaoxJhlT5swh20lIWaNoPHLOALXjYDlgYrSNG5pFMV5UU7Fcf11W5VlxZxoAq8JsXwfdiVaFB4a6rrx9ws4Ao6AI+AIOAKOgCOwbgi4YLFu0PqFHQFHwBFwBK4SAUg7SD1Ie1aDQ7QiWkA0QKiyQdLfKCP5Np4DfI8R0ohjfB5iF/Kfz0BmWKz7zSQEjVSh/JQPkpJjJOGFwKSMCC2sgqcueJiQNNvydSAoEErGPDEQGjj3dTJWz/+W7I0yBAk8MbgmAgZkKfc72ryGxQEn86YAI4Qh7sf5lvsDMrVOUOrbpiFg3jgQbogK5CXhNf0Ezxg8Kugj721KiFjH2OCcpRvj4RtHDiL4kbQeopz+YRviBNf9f2WMOwQNxAyEC0h3+gtj00MYLQPyZQ4hsuJJgchIqDfG4IkGR+YA5jpLDnx1V/azHYEdgsDSkHGW86aVJfFEJyvKKkyUedWOkyKRR+VMpIUCg7xcDFXF7wRpFxVjjN8LzK18B46dF9kOaUqvpiPgCDgCjoAj4Ag4AqtCwAWLVcHkJzkCjoAj4AhsEAK2yh+SFJEC0h7CHS8DCAZWgUPgskoSIgJvAzwTCH0DCcHnIPEtobURrete/MaTYul9LM62eT/gMYFHBeID4XzYIKEJ5wThDIEJEc2GiAChDHFM2B7q+7LmHDAg9BXhnxAdIEQhQiGj8UZ5SAY5ClkNboSAQgyBtPmSjHKBJWIFuIG75a7YTHGnqfqO3ZlHBW2NsIUQgUiAdxEb4cK+Q0YOhNGN41e7jYoVfJY+9SbZq2X3yRDGflfGWGJMkdidfoRggbjB2HLSbwT1ZfJY8K55WSD+ICgxn4E1Y/MJ2VdkNgavtg39fEdgxyIgoSJut9LWVDudGObFvtCOp4oibg0Gxd4yRDNpVZ4uyyjRF9pUXIUzUi0sbwzfk4SGqtzLYsd2H6+4I+AIOAKOgCPgCIw5Ai5YjHkDefEcAUfAEdhhCBhZbuGcIPtY2Q1BCrFPKKOvl0HscwwCFcKe1eK3yAizQggIVjNzHNFjswh4EysgnyEoES0w6kRd2Dj+WRnkpSULpV6QyRCZnEf5eQ/vCUQOrovAwcps6kxoIIQHBAlw4FrkqfgDGfk/IEk/LuO6vEYIgWzmOmDEa/AeixBaKsdO3RCxaHf2Jh4hxr1WhjcN4b8QMdZ74x7kWmAbFUL+H/1PP0MU/EsZohiJ4M2bZ7PG2XrjsRbXt1wxhGvDOwoxiHnNEqeDoW+OgCOwSgRuP7Yvml/oR2mS7FIEqNk4jnfnZXVLVYbJNA175XIxG2XpIwoRdSaKwkwSx6cGw7LIi6It4cK+/yxh9yrv6qc5Ao6AI+AIOAKOgCPgCGwUAi5YbBTSfh9HwBFwBByB1SJgXhaQ6ZB6iA+sNIfIZbU5ogWeCuRiYKUkBD1hkEzEQLDAy8CI1NXedy3Ps5A+fM9iCAXsEVCoiyUPf4VeI2Kw0hpvEULy4D3yDhkCAsl6WX0NFpDX1I0cFxCeEMeEgUK8QNxAnIAYhYyBaIZcxouC6yOMEFqKzyCCgBvl4XzMQ0AJhI3YLpOrgj4CmU3/J08FbYY3xd+4hnIhTvH5tdzIh2Ebnj0fkNHvyHmxoHpZmJVcngY7VrxYwcvCPCgQHpnP8JpiDkOEZOwzTjnHN0fAEbgCAp85eSE6P9+rFwAo/NNcWRR7hkXY20rD/t5ivrcKxWQUx5NRlCSpXC6Gw2JSE9LhNIkmyyrOo1CekqDBYoez8rIYupeFdzlHwBFwBBwBR8ARcATGDwEXLMavTbxEjoAj4Ag4ApcQgESHtIdcZ+U5IgAhHT4vg9yH2GcPeQ+J/7DsuMxiwhNiCcGjq3BN4jWijSJRTayAnERgQGiBjEao4H+OQ0xDuLCa/c2UsakHAgafJ2wUdSF8DCGcqIslG0eggeyk7tQPHF7YXA/SE4w4F3GHUD7kAkGoQMDhfPOoqMNiyOqcFRuIj27nW9POllN8s1AAACAASURBVISd/o3gRrvjNfO9TfvzerXbz+pE+hHtjIhAXhP6CZ42iF30J3JhfEJGH/nnq73wMue9W8cwvIN+RvYXMvphPUYlXtDfhjtZuFgGM0RHPFPubN4bDVfHvOCCxXV0SP/ozkAAseL0ucV2v5+35DUxl6bRkWGojkdJ2Ktk28fztNylKFDypaiKsgx7kixt9YeFNIxySmktyMf9iAYaz7/8TmDhgIdj2xldx2vpCDgCjoAj4Ag4AlsMAR4sfXMEHAFHwBEYAwSaHAjMyzY32x6i3cj2ryLdRTSPQemvvwjL5ICgYpDqrBSn3ngQsGd1MuFxIPkg7xEDWOlNHgeEADwGCFWDGGChoYbCaV29CJa0HyIF5YYYQWxAeLBQMAgsrKi2JNiQzNRrt4zPQaRANCPCEHYH8pdEy1wDDCC5IbipL+INRDc5PMj3ASYIHBzDwwJiGlKGexgharkH6nAYLlQIhQ3YlvGsoB0RsRCM6Mff2rQxAhbtvJrtXzXtSj+hL9DH6EOIVPQF2p7+RB+kf3AvhD2O453zehlhxqx/XemehB3D+2PpRl/9t819/kx7hIxnJVggmvkmBNT+tDdtAH6EhiJ8HXgyjh+VMa/V8zteGr45Ao7AVyPw3z/9eBLF0aS8JmYGw+J4lsYvXuwOX6NwUPviUM4s9IqOji9WZVXGSRRaaRKGerMqyyeGRXlR4aC+1B8UT0rNwOOQ70rmytK9LLy3OQKOgCPgCDgCjoAjMF4IuIfFeLWHl8YRcAR2NgKW88DmZva2Ah6ya3Ql4LqS72PSDBYaysIWUSyIeEhXwhqxohviH3IXYpTzTcSAtLUwK7zeyM3iYiO2QBSzap6yUg/EFYQU3oPktSThCBCUl+Tax5rPQaSY8MLnIDUhpfks26dkeFDgscFnLaQQ/4MHRDWkDPUHMwvZU5Oi6y3gNGX03VcjYOOcPkE4L8Yy7f+3ZIQIutJGImzCop2Q/XLzedoYUYpQaJZA3cRNE0GZQ3hNP2Sjf3G+5VdB7EC4oC9BrP+PMo6NbggdiIO3LjnOuPxJGQQ8YkXt+SSSHk+PgXta1GjRzuDHWGTP+Gf8Mm4Z0x5Pf0mn8n8dgVEEFL4pPnX6YjY91Z7QLDejRQI3D4bVlPJUdHp9wkDpe6+KJMhXM5r8WnFIWvKy6LSyqF8WMe4VT/XyspMk5aAo6+9Dviv5Pu7q2ivmcJKY4Q3hCDgCjoAj4Ag4Ao6AI7DBCLhgscGA++0cAUfAEViKQLMyH8IRQpG9GSSmhe+pH6plPFSzcdy2jQp1tBmNZ2Gh+L4i1I2RqeSsAA+8CCDuESog6FmlDAnB5zifnBHgudFuKEYSW7n4//GmTJDSeFNAVkNcUhfIE4yQPYR3YvU1IXzwtEB8MC8TCGD+h+TkOi+TQXpCflpyckQQ+pKFnAE760cIFdu5v6iqY73Z2GY80wdoJ5Km/7gMD5qVNvrJP5XdJ2MOIEcFfR9Bylbl29yw0jVMqLD3cwkKjCHKxDXwvCBkEf2FuecBGX0RYQUvjHtkCGiMwaWChV0T7wFyWyAo/oaM8FN/pPuQp4E+uGLf2yFeBeBKO+ERhacV8wPj2QTXldrOjzsCOxoBCQr1d+pCdzARp/Ge6Xa2S1/yWW8w2NPr5XNyqJhKoqRTlMV+nTgbR5HmtqKQc0WWF9FQ3hax3Aln0igcL+L44SQu5XBR8T3KvNhzD4sd3b288o6AI+AIOAKOgCMwhgi4YDGGjeJFcgQcgR2HgJHpRmZabgaId0hoYp+zAhfjfwv1Ahk/XBJKacuGjFohtJWqV0F0ggkkLcTtS2WQ8pD3YIY4wf94WoAZRCvnQw5CBK64cnKdeprlsKCtEFFoJ8oDSY3wQPshplBWyg1pfLcM4hoyGAGC82lL6sb5hPxhRTwhrrjujTIED64PBmDDca5HnSkD3/HUvTYXKoTC5m60E22GQIWRnwKB6j0y2n+ljTb/PtnvyehD1t/ZX5enVeP5UAsdEhUYW/Qh6zuIDHhLmKfT1+s1/Qyh5S1XgJL6UeZ3yf6L7FdliC1cf6fmajAcEXPe3rQl45354REZr7ftptwDo3Wrv/NeftOsi6fbtsXXvGK1Z1qvn3ei0N8/7Bd7JUIoslO1b1iVs3FVDRAtBnnRyvMyZEmi30ZhUd97U4qamSnfRVu/JXpVHE1r/8JYB8qqOKlzmPdSCSIr5rJwD4s1b0u/oCPgCDgCjoAj4Ag4AldEwAWLK0LkJzgCjoAjsDYILJOjgQuPhmthxS0kO6uuCakCOYghVEAAEloIcotjfA6CyzwzuNbzQv6sTanH4iqQsqyCpM4WBgpyH+8DCNA6aXSDERhyjP/BDXz4f6M2C/eDGIE4Ye1DmyFMWLks1BcxtMljQEgdiBNWpCPQEIPC2p1VoKym/4yM69JHWFmPxwbhedio49KV2tYf3Ktio1p/mftICLA+wZh+gwyyn1BL9N9Xy+gby22/qIO/JmPskxeCMcCYN6+j9aiVeWmYqECf5bcihmDCuOO9t8rIufEDTd9jXC63UccfburwU9ojxkHYX9bbYj0qNibXtLBwiD4IkRbirbfDwmYhVGy019uYdAEvxjUiQH+ZUv7suWiQH0zSeHcnTaYU4qmdD/KW3CWyS2GiokmpGLyeUq4LCfWhkHjRUl6LWX0ZR/K4KNTzbkij6Bm9eUa/y5i7+K7ltxVzq4to19hA/jFHwBFwBBwBR8ARcATWEgEXLNYSTb+WI+AIOAJXj4CtZmY+hsAyrwoIPV5jloAXYhMxgwdqciPwHiQ3D9zsMbbt9tBNfUdXZeNVYHkhwAlRAPwIVwM+EA+sSgefelXzBuZrMK8IiEkEBIQEI+csrwbtBGFNmWlTys3yY8I60QcIDUSb0u60JfVlzzHqTbgoBAvqCcGMt4Yl1bZ7WTkQK/S2b5uBgMQK2ty8fQirhJfC18hubtqMdsOTgfFs2+80731ce8I0fVH2tAht2nvdthVCMtHvuO+gCR+F4MAYI/QafRWvCTydqNf/dJnC4VFAP0Z4Ick0OTjo+zuNHKS+tD39AsERQ6zciVslrwsT7PG2uC5voZ0I4E6rc5rGURKHLE2TRCLEbFGFfUqufagK0UylXBUK8ZSmaVQo0XauARbr/baOdauyiOI4TGTys9D34byiQ8VlWR5QcMTHmrEIlJGHhdppPcrr6wg4Ao6AI+AIOALjjIALFuPcOl42R8AR2EkIQGQxJ0NksTKfVfSEf4HIhiA0bwKIeLwIjJiGuIaw5hjkNQQoJNB1h4sZF/Abwr3USkjzGACTEzKI4FFRAGIVMcAS2JpHQ6TP6jIbkrvBwr7QZrQBq+oRGNgo6wGZJd6G8CW8FRsrrmlD2hci14hiCBUMTwrqxXUhfhE5OIfzEUdGBZ2dRgI3EI7XrhErGMPkdaAPvKbZM7bpB2yflpkgyf9/IXt/0+b0A7wRCPO1rmLFKpGzvs08Q5k+JKPfMs4oNwLhj6xwLUJh/WBjJAr/32XmJcTnd8rG/I7HDBtzFXO9iZrbBoNGiFhtyCe+rzJ9hn6Ve5iobdMNrqkiCs203Odq1V1qQ67v8bwqy8X+MI/zotojCWLQypIL+o5fjCRaTLXTRCeWSl7RqvKC78y0lcWLUYjrUHoSPE7ol9YT/UGY16+C0+FSyElPeH9NreUfcgQcAUfAEXAEHAFHYP0QcMFi/bD1KzsCjoAjsBoEjFzmwRoCHkIaEhoyG2IbYpMHbWLc89rizD+q1xBdrLhnlTMkmK28h9CHHLeYzNuFwLYVuAg04AA+EH5gRp1ZpU7IHIgvSHyIiM1atQvmtCltAkGNcEGZKC/l5n/aGMIaYhpCl/IiTPAZ6sL5hIEiJwcbhDCr8SFXqP9m17Eplu9GEWhCQPH7CjL/oIx8IySpfrcMLwtEDNteoRf/sWl3zvuw7Ldk9AU2+tE4jl/KhIhCXhXGH9s/k31E9ksy+upK23v1BkLdr8v+QIbHBeN3W+e2wINFfYM6IjgyJzDPz5ZRcn6YTOT/4v0fXuoK9bx232Jx9FdLAFv/5vy6z0i4cNHiMoNnB79VxXGU50Wp3zZRrs6SZWm0qFQUT8vLYk5Cxr5EUsWgKKphr6hIth2FqCWBosDLIi+GCB7TChM1Q44L5b6w0JGjfXAHw+tVdwQcAUfAEXAEHAFHYLwQcMFivNrDS+MIOAI7D4HRnAcQgKyyh8iGsIR8h7iG4CLWOQTXy5tjeFyQiNnyOkCAcS5CBmFkILYhwknKvZ0SLiNAQPohBhipS6/hOOQpxCdYQEbUKyc3yLNiac+FBLGwULwHGcd3LmXHYwIRAuKa9iKHBR4TnEMiZspO25G3gjZnVTZ1oW6Wv4Br16G/Nql+S+vr/9NIl/JVIEgR5ocxelyGaEFOkjuaNgcrBCfCAeFd8JsyhCtCBTFuLZb6WGG6Qsio58K1qe702d+Xfa+M/Bb05ZWSib9I72HUFby+rM+f0H7FxLcr3H+sMFpFYRjbzFPMBYMiztJ+OvPUE7N325xm3nHmzWKXHEfRatnqWpinqwjxZDmKwIR5nVBRhXtarKI3bcNTVhDmKnleyKOiVNqKWB4VcU8qRE95LBaUu2JWXhI9eVl0h0URKTRUrIhPURJVcRZHi7wsyzCjL1El4A7SLqr9EiselA002BhXfLeO5Zy7DZvXq+QIOAKOgCPgCDgCjsCqEXDBYtVQ+YmOgCPgCKwbAkZuQ2LiRQHRiYcEwgOvXyYjBAvnQWzjQQCxSWx7iFFW5/OaOZ2kuBifh9SucxmQ8HsbEdvU3wg9SwpsORuMeIAEW+0q3/VoWO5P2RCbLM8EXhW0C4IF3jSUmfaG2IWwRJjg/RMySwIKCQyhglfJc+3ZfJZybxkicz1AHqdrinBn/CE43i5DqMDzAI+KFzflxOMCkYKxSy6ID8oQGREeEacsD40lvh6n6q2mLPR56kBy7gdlCHH/WPa1l/nwj+s9xsP/J/uADG8x5rrN8oxaTT2v55x6jFdRPMyjVjZMJ7tfPPC24RcOfgPiJUI1ggbn2FxAX9iKIf5iiQ7VqGih15fDLW9CQlFvy2vhc9v19LRt+Fl5RuTykgjdXp7GSZS2quRcWwm1i6raKxuq4yi7RaywUVVHOSqqoNcKDdXVe6neG8gb42QcVafjEH+5VxUP6xS+b12s2IZ9xavkCDgCjoAj4Ag4AlsfARcstn4beg0cAUdgayNgxDvENGQVyWzZIKoQKywnwz16Tcz3R2ScC8mH14W9D+n5ahlkKUQ55Bd7rgMJJM2iKreRaDGaWBwMqaPhNrpKeTN6h4knlBGvCDZWkVvCYoQH2gcxwzwl+N/Op90QKSysF3VbmqeCazqhtwmtK2Fi6WZeUkf1xmtliIiIUBhiI2Maz4PXychJ8QsyS8ZNonXGMBveNFtVrAjygLDQKs8KozrcUVO3f6D9t1ymqQiF9QMyC5WE+AouK3pbbEKzX/ctG++bTh63W3nSefzMxM0X2sXCUf1/7OzEzXjTIUrSL5gL+H3OfMAcUL/WCnMTLJctyxiFjKIOlsPnanCzebMOjYWnhntZXA182/7cehHAYFhIh4iejuOE30JHirJQAKgIT9JhFIeefuYECRtaoqGxpGQXUirOKwl3e5gXiX4FsXrjgqJGoWd0ZcxT/O5iw4vjq0Aco3G17RvYK+gIOAKOgCPgCDgCjsAoAi5YeH9wBBwBR2DzETDimTkZMYKV+KywR7CwEECQoRChkNl4WfA+G8Qe+SvIjfDGZs8DOAZZDgnGan5I0W4THmq7rF4GN/OiMI8KMBkHotPKBgEN9pTJEqIT+okV1YgSvGdJ0yEnaVfM4mtbPo7tJDY1XXdb7Oh/EMx4E0C8W44KBETa/AXN+KSNES0IAUaeEoQL2huSHo+CYUP4bwtQVBfqfkYkPTktION/W3av7PuXVJB+zvzE9jYZnhl4jH1Mhihrgt6Wx+Wn3vQX4e//2Tf3JFIsLGa7Zs93Dh8t43Tfmcmj8yGOS4WuqecBVoJr8mD+2CtClfB2tgKcvsbrcRcq7TtraU6O1bSh5xNYDUo78BwJBwgKfB8qrFMYyNHiGQkTxy65JkZnoiS0lcJCYZ+UuSKujmRJpETbUVGFKs9Sjoehzr+oDz81zKuBxpaNJ76HK66/A2H1KjsCjoAj4Ag4Ao6AIzC2CLhgMbZN4wVzBByB7YYAD9LLbHg+GLnN25wEiXeXjBXa5oFBcm2IIMhuQsvcLyP8TP2wLftGGd4VPNBb8mbyXUAWIlywr5/t65WIUbTlRIuV8GvqjwuJ4cd+w8mHZcpXl0HlgmS0lfPsTZQw4YL3aRsTmixnhdVh1JuES/o2HggwVi0MG4Ii7UTbIlIgJDLuLMTNbXr9BRleNnyGsFCIFtu6bSVcDCRakFSbUFgPyz4nQ9z5saYJTazgX7xR/r3shOzfyX5VRqisLS9aiGiN7njmQ/GnbnxvW/vDedw6dHbqWPXM7J3l2YmbdoWsM6dQNYdEsGZiW59UzP1eHIVWFMoTIliZGyw3is0N4zx/U1ZLxH6tidTr70T3shiPiW7cSkEuiqESZ6ujnVNoqNNRkpwv8ypPWqGtATKt49FwiMbPj64oL4riZJoyruRdkZdfKasS4RjPN7572basZ9u4tY2XxxFwBBwBR8ARcAQcgbVCwAWLtULSr+MIOAKOwLUjYIKFJR+F6GT1NWbEJivyWbWNNwVCBMQoK5ZZoc8xRAxCJOyVQQxCfpPEl3mesAesAme1bh12SCT6ZiWjvnaUrvDJRjDYcKFilRUCd9rCiLxRrwvzDoGYtRBezxGS2yiM1yqhGs/TloSCsjBQjL1XyEiqTSgjxi7eTu+UMWbxoPhTGd4VCBbmIWV5Gsa1v65ZI0i0GAo7hBrmIfbMS98h+yHZcvktEDT+mQzR5+MNppbDZ83KtVEXQqzQvaIL7YOtdj5/5NTMHXNpyCfOzN62cH76WKff3n8sjtEp4mfSJNqjFeFHpb0i1CyWZdxXxuCTCmPT0+pwyFVEzqFWg4+7YGHjY9UwL5PjYtuPjVWD4yeOIoB3xFPySLok8FdKqB2FU2UcMsV5mlF4qPMKG3VGnacnAXC/fuvsVt4LDbBqXuPqSf1/Wlm5nypDwZzC4o7SvSu8gzkCjoAj4Ag4Ao6AIzB+CLhgMX5t4iVyBByBnYeAhcGwlfYIFeSnIAQUxyBAbaUqhDbeFm+VQYj+uYxVtxwjpAjJfsllcaQxVhJyDcJIWU4E8ikMmpX/KBdODK1jn2vwxZHGEmuzt9AutrKTNrTV9r7ac5n2aDxolr5jbkuj+1EsSTa/1uQuohO/n/CquFuGZxOJ7skxgycBYY04h7GJdwEkPeQahL0lUbcxv449b3wuTbgriRb0ecJhIdrcICNMFEnn8UgZ3czr4pd08NdkeFt8Tp/HS2zFuUr3GNeNvpl1s13ZQmvfrk5+MStbU9kgmztYZe3ZMuvc0m6lcbudzolQ3avl4JrXkxNRqE7pdaTs3BODQc7c/YAMwaKQCLI4xqIF4405LnEPiXHtkluzXCNhoZR/oiwkWiirdtgVR6VCP4WzSZRMZ2m0S9m2JyVqTFdFtVjFUVeCxXnlrTgv0eJB+Vw8qc+d1edcrNia3cBL7Qg4Ao6AI+AIOAI7BAEXLHZIQ3s1HQFHYOwRMAKTPYQrpB5iA+Q1JCdkKBt5LRAcOA/y6s9kCBvEz+cBHHIMEpCV3TW51fyPRwaEH54YHGP1Mvt8O3pbjGlrj4b/AfvRGGGeo+LqGq1etd4YuDJmLNkvYoElKEYosjwnayHOMaYOyiDZCdkG8c5YY0U8Y/ajTZnwqjglg3zH64IxfNmkyVdX/S17NnMUcw8EPPMUYgS5K96+Qo2+Qcf/qwwxFsGDz221MFq1YFHEWdLN5rJnZm7bnaXpXNmZuXFyopPF7c6ekEZKGJx02ml6tKwUBKpSv6nCgd5Ac3RRHC2TSJ528cW8KFkVjrdcLtFiMMaixY4S5LbsaNyCBR8RLfC00HxQZUVZe1u0+8NhLLGCvndWsRgPaOZnzj1ZlCVz9Je1fzyJ4/n+IPe5eAu2vRfZEXAEHAFHwBFwBHYWAi5Y7Kz29to6Ao7AGCJgoYxGcjBAuPIA/hkZD994TxyrH8IvrbKFBIXsY8U2D94YxyBRETYgyCx5LV4YEKuIHBB9eF78pYx7QHwZseSr+te5bywTsso9W64OcxMo+BT9F/HAcr5YXhCOk7QZcpuwW/RrcK6TmGuMIQyt2uNiJAwU92G8EM7IxhMChY0jxt2XZIxRvCy4B2MO0eLidkqofXVNtuzZrL7H6+R3m3c/oT2eFy+UvXnkE+aR9C91jPntf5b9ngzRAhHoWvMjrEEVVneJJhwUJysPcDGtvqfV4Arn15mcSSembpqcTBfiqjfZHYRhNDF9KsviuNNRt64kcOTlbXlVFnlRPTOZZNFQL7u9cFKiBaH/qDueFmOXLFihnSp5Vrhgsbou4mddAwIjogVCRHeYFxo5EXNCojme30WVXOtyeVZ0NXFfKKpqMYnieXlZXFA+i0Kf5zeTb46AI+AIOAKOgCPgCDgCY4yACxZj3DheNEfAEdiRCFg4DR66IVnNY4LXkLB3yHgwt1wHEHyIF5Cjx2R8jjA0FjoKkhWRgvn+PhkP+ISYIvY+hC6Jf1mF3heZ5qLFjuxy41Hpy4R8GvVEQSDAkwICGzGOMYHxP/lbeA/Bgvfo33gVISxAoEJSEQrtWvK3cF3GEHlgKA+kOWNnV2OPaU/YNTwuuBfvk9R10cWKZfsX85zNbwg9H5bhlXJngyEfAm+MtmQj6BPeGMxhtCU5fZgLx1b4g1j9tX/zk6GVX9Q8HM3NTx7ZOzm8sCcM40OL0wcOKC/wyWxqclj1htPtifTpJEkWJlrJjHwsbhxGYWaynQYRrYuTnWxioTvYm2XFVy7Md/sSLWrRbVxj70u0KBAtEC+WbX0/6AhcJwKNaME8UOf+krcF8zFzPXO0vhOqc0rLnUdxICTUsE+W7kbou85b+8cdAUfAEXAEHAFHwBFwBDYAARcsNgBkv4Uj4Ag4AleJAA/WrBiHhOWBnNdflkGakmibh/LPNf+Tr4JwNL8jI3wK5C1EKccRIFjJDHkKicsqZsQM3md1OqIFK3W5HqrFQEzu2K9avkos/fStiYB5U5hAYSE8GAuENZuRIcZdSrx6SYSjj/MaTyP+R0CAxKKvE0qNsVCLcurrxVV4WlAWE0hONK/JFUM5GJOMGTwpKA9kOiQ6YY9yFyuu2PkgtMHsg037fZ/2Pypjnltu+zkdxMsCTzPwJyQe89eqvWauWKI1PAEPizu+8E9aWu596InZl8yem7z5/GS3f3Zm8Oyt3eLodJVN3DjRaRUT7VY0qJIjrSw5VCqmjSSxbhyHXpak/XSyStutRNfICuW5SHu94ZGqGp6WqHFa12e1+FjWXWLFWJZrafOOeMHwFv1xVCB9TnARzmvYM/xSa4FAI9gRHo2+Rtg95bao+M5oPOsUXO2veyFjxRdlrAXwfg1HwBFwBBwBR8ARcAQ2AAEXLDYAZL+FI+AIOALXgAAP1pC0kKBsxHCHmPu4DC+KT8lYeUzuCohYYsNDlLJC2fJUcAyylhXMrDTnf8QLQtpwXUhfrmuE78LVhsy5hnpt6keqD9YhfG6Lvq7GJOh/8hGc1/89vWaDmCYEF6IOG3g+qPed6NjYloM0pK1MsDDaifbhvUMyvBnoz3hS4Hl0jwzSimTY/L5BSHhR06YQjwh2J5rjPTw6Vila8FkLLcU1H27ub2Kfke4Ih3WuCgkVHnJkSX+5TFJssD2n8Fu0IyG13idDgP0e2a1LLsPc9YMywtp9VjYrYyyf0OeZ38YmKbfKEz39qe9OiyibuNje27rh4heOT1QLd07E+e1zxfm3lHtvnYjTXQpZMxxUWWuYJVk3TpIsz4u41UqSXF2/G3Il4i7vnF9QUJuqaud5eaDdjv8yirMLC4uDLSEILGm/Tft3iTBBOUyYMO8p8LTcQrzH/1stX8qm4buZN25Eu1JtbAsuTPB+LjTZuHojbSZufm9HwBFwBBwBR8ARcATGGQEXLMa5dbxsjoAjsFMR4CGbB2/IT8QEiFBbQQjBfqwxknLfL3ujDI8KvCtsQ4jY3xhhayBZWWVOgm6uyQpwiBpCSSF08FlWrxMyZ7VE7ti2j8QH6gKGiDdg9mIZZGe9yl7vg8VbZJDeu/S/CUOQnghCrM7/QxmC0L16HyzB0DxUIFZTCRlOTF9nLxjJ3WJXol8a4cTvFNoI4QJxgr3lpKANwZ+2eImM0Gf0dc7B44HPmncS7ch1aV/2HCenxWrDQ/E5rovIhzhCmRC1yFfBeFJS5LocTiJfe3+gLZm3yG3xd2RfbC61VLRgDN7dGG38E02bIuDWYb+uvQjX/0mEiqY8nYPzX7wpj1uvnunvCmk5+Mdn+0+/qMgmQ6vVClOD02ExueOZMuko33aatNvZvDp2UYZ4l0JDzeIFlLXifJhHE2laHtW0PJcm8dNxHH85iaPus8rFMr9At/QNBERWrwTEqMeEnWOCKHOJjWuOASh7m2PoT8wX/O9je8y72ogo4aHIxrytvHiOgCPgCDgCjoAj4AhcCQEXLK6EkL/vCDgCjsDmIGCruiFJINkRLxAXiJXP/xB2zOFfkCFWWBJu3mfFMauVIeoh7H9fBtlLmBVC5ECyctxWovMeZCvXh8hdFFnWXeXq881BZ8ldJShAMiHGQFhTh1GRAnHGPE8gsiG6P90cg+SGkDK265V6bcQ313yFDDIafBE9bmvuU4sXui+kNaQWIsdJCRhOlFx9jwB/tqVCBVjSnmCO1wsiEmQ0q+ohp2kbwgkhJuFJQSgoPC9YfU8SbFZLI+iRzJm2Y7xwDTbarE7Y3XgVLdtuI14BlYhoBDCELcYkQ1Cf6AAAIABJREFU7U+/om9Qpp7OHWtCUzkFauJ2zPMKgDHzE6GffkXGWHyn7AdkhPxioy1te69e0A++XUb7Mk4/KcOjzLxiRk5f35eNWIFXG+Vgfn1VUuXfNjG8cFuetPakZT+U8XSoWpP9VlydG3SmLkSdzu68qtKyCO1SLdSKY0JCqXdWPcXel1qRzERJpEg31UmFiXpmOKzSYZ7P7prpnHXB4q/bc2nIptGE5zrLhE76iAkYzCEcZ6O9mH9YBMAx5hv6EG3J3DDU9SxfwrKdyENGre/Y8qs7Ao6AI+AIOAKOgCPgCOwsBFyw2Fnt7bV1BByBrYWAkaiEgoIUtUSzrOiGIGe1N+TtJ2QIGpC0H2oIFlaBEz4HMpd4+3/evOYzrDaH/GM1KcZqcbwsIGcgCPHoGIrIHYov2yoEPIk2qcc/lEFIQUaBCRggVrBHpDkWklY3FAO8K2qPEhlizctkbLyGrIJsRNiAvAIvzuU9RBFECu6HUITYA0Y/K0MM4n/flkFgmaTatpLZBAtb6UyfpL04Dp6IEnhQPCijj9J36f+89zoZ+VxMUKItbpfR5nyGNuK3DmIc7cNqfUQHyEj6ua2kXk0/p69ApnNviHXG4diECpMgsVK/M4K23nPemIsWYMpYo33B+L/JSLD971eoIHPdZ5r3ECJ/WYZ31CPNdTZESJJYYZ47zBuILG+mz0VV9ZpYU3ciNULJt8Og3B0WOgeGw7nDJzutLC6zNCmHRTIsi91pGvfk39Yvi1LOFPGkcltIBSuLVBGiirzcXYVKHihVf6Gb79J4Qpz2bWUEzNOFuZvvA/5n/mDuZiPPDXMD4xphlDmH9xAheY/P0ReZfzjPxvqG9Kerbdhm/EdjPravtlp+viPgCDgCjoAj4Ag4Ao7ADkXABYsd2vBebUfAERg/BCQOLFcoYpcbQWIJhpm7IasgyFhVjpAByYLYgCDBe5BmrDqHBIaE4X8IfUKuQOpBCpO4FlIGUQPyFkKX8xBBIGXjy60+HwcE5eFAfb9O9g7ZzTILBQQ25h1BnebD1As7IZ6cDrtffzgkU4PQ0mL8wblhyGZuD+c+ciqc/+Ri6D9yrKk7jQFpxfUttjlYmdDDNUmETluA/z+XParyEM7mg/K0AGffvhoB6+S20hkSEBLRVkDTnxETwA+hCKLaQpdBLHLs62V4EdHWCBVGQprwgajExniA+P4TGeMDoeJYc308MbgeohZJuK8YGqpJoI1QAYE5dpuIyufKNBqv/xUvOlzjcsP+GUQZcK9Ebhr5Wo0pwUlZmaMQB+kPjDEEi78pY75aaWPM44EG+UzOEoQLC6235uJS41FhRDh96pgMcYy59t0y9TlJELUuRtrsbugMz4con3+0laaPDNLsiLwn4riMkyyKZpI4JFWI5d0WilSeFWkcF71BXkj06OVlOS0VY0YaxxMSMvqzU0nxP3z9HWNJnm/24FD/p88zpzDmMdrEckIxh/N6Fw4sGvvMNTQQcz2eecwnvOb7Fg8t3uPz/M/4fy4vwmbXc7n740k1pmN6HOHyMjkCjoAj4Ag4Ao6AI+AIjCkCLliMacN4sRwBR8ARGEHA4mdD4EHe2cpQllTzP2QsZPprZYS/4TghjvDMYLU5oWsgdzl3dEU55DCEMEQM5I6tGocQRLyoPTvGSbSQIAARifcDdpcMUQZyCuKOlfYQlhb652yYuvNw2P0WMYUHbgitfWmIxV11v9wPE7dNhngir0WM4TNlmHxBFKZeNB0ufDILp38nCan4qXwB4goswezS6ul0z+lQ9vaHchEiHNwgJsENEQgiDJLynSonobo+L2OV9yMk9dZ+R26NZ8Vo2Cfaiv4Gvkb2sgIaxh3S13JPEPZsnwzhAU8KXr9KRtguNkhH+v3fvgyweB3hMQMBiXCB4MFqasYD7QVZyXUum7B5qzQcQoWEiXhmqh2du9BLOu006fbzqN8fspA/3j3bQbxUbueY+tb1FsFZjinBacQwwhJj6T/IGE/MTz9ymTb5Wr33dhnC0r+WnZD9qcQFhFwSoq/Gm2a1TW7kNn3srU1//KWmjJYXR9GdKnJYhGg4fzpv7/rS6d0v+Ex35qZ0OAxTaVYuyJuikDycoW3Iy6KjUFCIxYOyKoeJJAy9P9OuwgW1m6JHVf3Z6Y68LuJYbRer7Vy0GGmtRqxjfjHPCgshh8cOx4RcNC1RaL+apRHzo34jWmpOqIRx7ZHB+KDP0I/4LmSet+emDQ83dqUO2QiWa9m3r3RLf98RcAQcAUfAEXAEHAFHwBFYNwRcsFg3aP3CjoAj4AisDQKN5wWeFlwQ8g7vB4h7SBMLWwE5Rux+QhvdI4Og5RyItDfKWGmMsAHZd0xmIgjCBDHhOY+8F0Z47NVrEzi456YSIRIAILwRJ6gb4X4I7QPZzIpYyorwApkJDouhc/zGsPet7TB1t8SH3XMSK8qweH8cotk0zL22CNnBOOTPDrS0fhCmX7U3dG49KCGiDAf/Tisc/18nQu/BPJz9eB6ilvDNJ0M0UYbOzfMhPz0TBk8/GyaP79N7N4VicRDO/VFP6Zs74cIn9ob8HF4ekOSU4w0yVnl/SeUnbNcXJFxsW3JxhZBPqnbddpa4FoIXItBWNNNHWb3Mnvf4XYII9HIZXiyIUvRPRAvOM7GC69L3r7R9l06AcPyYjJX3CCL0GwQnW3HNdS4bn/5KNxmH9yFq52Y6aX9YtJPeYKKVJVqIn+Td/nA4M9mOkiSavrg4KEWIS4QMMWKGSG/wzkV8dzdbtBjJF7IUztrbQoLDp7RnDkNw+lPZ/yFDdKLfjG42xpjTflzG2KMP/VvaXdehrREursnjogn9BG4Ix8w/iMTc0/KtIAT/8POLVD2iHr8YV/mwmNzzm739d10I7c5taSe9EFXxU5InpuMo7siZrqPKxjLJFJV0i5ApAXceR+GiPC7OKpHFvNru4SzFLyMyEXAcut9YlKERK2gb5l+bT5g3aKu++r7Eo6jQnylhvF+4yuKqlFBUlmXQd+1Qx/WymlB78RqBFG8uRH82BA7EvtozyzdHwBFwBBwBR8ARcAQcAUfAEVgfBFywWB9c/aqOgCPgCKwXAhBj5iUB0WoxuFl9DkHHKvKXymxFKEQwq00xBA1Wm0L6sbIdIockxHwWUhei/VhzHchdzoH4KVBLNjKfhQh+iEjKQhnJPUG5WcEM8USdKBvCzS0yCyFEPbph7zfuCu3d7TD90onQ2rsr5IsPhGz2YJh9+WRo3zgRkknhly6G6OUitKokVINeaN2s6xYiMkVhhUIeGLc8HqZfs0fh4tvhwqeeCu0bdoVS51VHLmgB7s21AJLPK3DL2Sgc+o6JMDz/srDr3iic/3ih82clbDwQqpI6EF8fbxC8Xz6keuGxAVmOOHRCAgZl307baFwziyFPH+I1RB/iEkQr/ZM2xfPEPGQgAwntxUpmyGkEKFbLgxVtjUh1tZvlaUGooH9YjHpCDXFfyGs2LYKvLKfG8+6xQqi2qy3HdZ8vMvZy16g9KxZ6wyxL4ql2pnX7VbVHZS/Ew/bPXuiG4VD8fKVV/HFoTU20eCOW18W8Vpt3O610MBomarkbjYacuu7KXNsF6BeseKftmKvwsmB8IUqMbsyDoxsiJwKYeY39mV5/RcIDfYNrIlzYvLqcMGv9mLnWPCroT/Tl18vIVcHqfeYm+uty241iwz9YJa3f6B16yWfLvcdmomwypFlHeSnUt8tql/a6djTMiyKXGjFBhECJFErGXc5r9Hw5iaNH07S6IMGip7br5jkpun0zBBqxAkxMsLDXfH9oLMi7qgy740zCUhlPlqE6KkVIsl3U0RjplFH0uDxaHpOgcZvaYkKYa56u9N1XC1K3yQibSL+rvz+VZPuqRfzL5ZnZbMHQe5Ij4Ag4Ao6AI+AIOAKOgCMwTgi4YDFOreFlcQQcAUdgdQhAlFhICvas9oTQxXuC138lg1CDhEPUgMBjVTnvQZjXBI6M60AcW6gMI5bZ46HBuRC6dTxwEbrFeosWIvT5XiIhNiuiWWFvniSU91EZAgXHIBoJ73NChiBwd0hnHgyHv3+PPCGmFOIpDf0nJDQcbYXJmb3KWTEM6T7VNRuErMNq2WNNvVTPFiSkVtFm3BushONEGrJ9hJj6isJIzSp81NHQO6mwLele5cHQ4ue8H+LpVijmJIB0opCevzG0FmdD2rkYZl/9VDj7py8MC5/thSH81nM5RghTg0CBeARR/4TqS1v9oYQL6rPVNwjCUQNX+g6YsqfOJIAHZ8QI+if9DA8gCEHCaHEufZpzyFeARwXE8LVutCFEMvdCBGE80IcYL4hhzxMt9P9Vk5DXWrCr/ZwI0mU/AlF7+7F9yTAvMyzL4qnBsNw9NZnNaaX4wVYaHxjmIbmw0JeaEV9st7O+8iL0er38yaKsLk5PtaaLydZAIgYEPthfk+fB1dbnGs+nffD4QlD9Axmr34/Jvq1pz5Uuy5z2r5o3/6H2f0sG8czn6WuIGfQJ5kn6KfMefZn+wvxIH4S4pn8SLojPMHcylxKujO1y4uOvRFX5L8ukPZiaf2QqU3Ltfnta4eWqM5pXh0UpT4qoPCJ2fCjBqaXQT+qv8reoqq48Y1TnqBXHup80NTww5FuRtzOFkfJtKQImzo96X+GpcqN8K16gFs3KorpVIkQljHfLU0VeMVUkMWhxWBSpju8T3p0kCl2EJAkZzBvkueC7kHkEYb++h8ZddbWixWVEv7Gdd7yLOQKOgCPgCDgCjoAj4Ag4ApuBgAsWm4G639MRcAQcgetHwEQLC39i/0PmsSIdUgWChVj9CBUQcJaE+HG9JmE0RBsrlFnxz+cg9TiXlaR8P7AindcbEi5H5D2kI0TT98t+S4Zowf+Ul0TK5OOAUKRMCBiUmW1RYsWXw/GfeGu4eN8JCRYzYequqZC0z4SJ2/shmX0oJNlrmjqxwp7rgo3hRP0gzCEgIdm5HwQlAtAtYeJWBI4qtA9/OpTFbaE482TonsjC8OwuZQOQgLFrKkSn50J7z/mQ74/C9L2Hw9Rtg7D4aB6e+k9fCIsPkBga7wCuTzvRDtyTleI/Jjugug8lWvxqU58ttWs8E0yooL0s4S0eFOAJlvQtCF2O8T75KWgL2hGPIEI/QQbzP2IbQgWhda53e3VzATyJ6EP0e4hnrv9JGf2AMm5J8rdZVR4jVMxIeFAsm30iXe8QIX5E4qLwrG6PkzAh+jvVe/N5rjwI0fD8IMQX+sM8FmGusGehuDDfl4iBC0aoHn3yfHm1ROz1NtI1fJ7xg8DAfPW/yH5e9k2yd8pecoXr/ezI+z+n14gOlmAZDw7zVKNPMwcw53DO18gYy4TXI/wTHh7MK7YhgC230ecQy05FWauQR8upas/RfYrZJWeKalbc+d6kqBblwibfCsIShTmlsECwGMah6up8ggEO8rxgvjqdJkk/jeLFlrxiPH/F8+C2OagOISZDDEWcZL49IED3pHE0iUkImpEHnMZLMkFekFjZzrOqOkR+EI0bxYxSHgupFVI6BvLEOK1Z+xld1LwQGScejusKg8zfdgQcAUfAEXAEHAFHwBFwBK4HARcsrgc9/6wj4Ag4AhuIwAqhaepoTSoGK/RZCQyZApF/nwxPhJqskRFr3Vb2Q8CxQhkCBlIHIoz/+SwkoIVJgYDjWuu6+l9kPXk3LnlJXCILIZxYdY8HBWIB5CAEka2GJocFBDQk+ELY+/bJsPsd94TZe6fCzCuOKBSUzk8eCbM3vkqCAnViaToE1gkZq6Opr+EEaQ5hjfcGWPG9CDnJ+Xh4UH8wIhdFW9d7LMT75V2xa0/In/7z0D8FIX5naN8k4jvbE+YOydtiQu1R9sLcmyYlduwL8596IDz9Kw+H/kmuR124JuQ5daSukJ7nhQOkKQm6P6v9WG9NvgoLSQNmFj6MPocwQz0RJ+iTtCMbxC248j7CBMc/I4N0/obmMxDR5CpZ640+z/1weaE/gz+r6ukLtD/l3JLb3l2TSmcQWpofdikvxeHF3vC4Dtwo74rDWpu/N4rjRfGxqVbop+1WWom4neh2B7MKESWuPOx5qjf/lDphn2X8c1PtvkJL0R4mBo4zJowd2hJRlnmLvsM4pu/RnwjXdKXtB0ZO+O2mf3yP9r8rI+8J8wxhnphDyK2C+PZDMpKAI7KNbs8l2W4OUq5fkH28KV8vn75h8eR7P8BE3JbNxlGxoHQi+bAq+2qLLE2jWakT6ovlgsjy82LMaZdM5/aqOMmrqHoqScKzSZIyjrZtPpwrNdoK71t/4G2ESMSKeyQADTQ2JPTEh+Q9cUCCT6bJqp3nhEdjOIRYYl5b50yBvS4y1Gf6+sKZU6aQI/qmOKLgW9Izqg/rXOYK+77lO2TNvhsVLmrZkHRW1zEIyXaNzeIfcwQcAUfAEXAEHAFHwBFwBK4eARcsrh4z/4Qj4Ag4AmOFQBOmCeFiNKyECRgQeAgTkGd4TEDqQdojDEDSmhAAEQNhjygAuQvph8DBuWwQZJclVK4GFJHzkHvfLIMAxCgbq5tZbU+5IJIg8CkHxBCr7tmsPqzWn1GuiUfDsX9yb5i8TTHHO60QzSgsUx3aCY8JPk/5qRvl5x7sR8O9cD1W8kNGsnFvBAtCgEC+Q2rzeYQJvAe471l5bHRCcqNyZdxYhOGFE+KtXqJw58PQf7wfoukkTN81o0TdaSgWng2Hvu1YmHvN8fDEfyrD2T94RFoGOFI26sj9jsk+Kvs67ids8HyBWP91iReUdxw36kD/MG8K9uCFuEPfA08LUYZQwwaO4AoZDpn8nTK8HegLtC8GQbyWG/2ZMFS04wMy+hM5DBDCMNrAPF/W8r4bdq2pSbSKqLPQHUxKpNgnR4kXKezNoXY7nRBJm5EfIU6iIkvSiwuL/bYaTnkSqkxhoQ7o/AvyznhIjUdC4ryXaa1/VaU/8+v3nVOC7uE4eVqskJTbSOpcOSkQaRnPkNWMcfrnSjkllmufd48cJJcKxvagjPlkdFsqVvAeHlMIw2w/LfuijHGOuMH8u/jQ9/9xTZDLEIUWJCY9Iv+JuVYWdxSeS55jyUWpSHMKX6R5JMLLokvOChHnZRpVi2UZPSV9mr686N4VyzVhfYw5iHaocx1p26++fUJCxaMKqHWzIm1NhjguE83OeVnFeVFmOqeM47iQN1JOiK6slRUaR8TkmlYwxDNFmc9o3Nyizkbf4juAeSzGw2mcxsiKiPgbjoAj4Ag4Ao6AI+AIOAKOwBZDwAWLLdZgXlxHwBFwBC6DAOSdiQoWHgOyH/Ib4ps537wtWJEMWQ6hD0GPQaZBKkPM2+pRyDWua0lpr7sBRMhDGpPPgfAtkMWQi6yGxaODVfkYx7mnrWCFbMYbgnrdL5sOB77l/nDLP3tn6BzdJXHgQYkICB+UnezEeGtYrPub9RrikDohxnAdyGpIQwsfY+FcwIP6Qnqxh3g3bMALzwDEHsgwwmn9lRJ6E+5pIZR5FqKp6TB8+NGQ3qBy5rPhwHv2BfGMoXNLO0zeejEM/9Ed4dGffjyc/cOBxAxLAg35xbUg7MEb4YgylsLq9yRa0FZjsYnMgwSmXWgHykqf4hi4UB9rP46BERvHCMPFnrYn+TsiEWIFxkZbQAaacLRW9cUbh4370vchGwkpBolck44yE4+2Yhz5uN/PO4rBPyvi9ZCSbR9vZ8kNomkn5G3RkxfFTFlFbTGvQyVwTqphrnj8od9Ko5miiOd6w/JZfZb2HCRpoig41YLUDOUfjvA8KUXIFluIkGUeMW+L/6zXn276HOPp22WWa+Jq+9ZSsWKlz9OvflPG/MBrPIoQMZhrcgkuZfh5hkAotJqeueQReVE8o7Y6qnG1lyTbapvTaoxpJX6ek3BRC5sSLxCcKyWuOBXFVU8hjJgbt2QIs6sF/irPt5wjCKCMZUId4jmoeSVqCdxYiA4VdKvI4khJ6WsU+9p3NAmo75cLwnYo3OMi17ll0LipppQv5GTj3ciaALBnvuB7aU09XDzp9lW2tp/uCDgCjoAj4Ag4Ao6AI7CtEXDBYls3r1fOEXAEdiACRrqawMD/GGQexBdkDgT4QzIIcohcSHoINM7hfyNwIZ0hxthf9ybyHbaOUDzkqkBE4F4IEW+WIaggWkAEITooB8XU+TBx23RoHyzD3OtboXOkH/J5vCpmwuQLZ0L75jskUvA5iGdW8SMyQEDjDcGe+yFEnJBBZkE2mVcA4YF4jTDA3nBiP1pf/gczysVry8tgyV0JFcN36QUl5H5Gdihkd+3X2t2Ozo5CebEbot3KcaGgPZ1bJkN5fy/c8qM3hd1vWAgnf6YXeo8b+UXdeQ2BT+gR6kBYm7uEG7ktTkq4oJ6bsomoM08KE7XAAmwRAdjoSwhGljOFFc7UheOcR5vSBrQ3x98wUhHq9ccyVrSPJstdq7oiYJHQG/LYPG3MgwhSc8tuhINK0lhh+eXOkyr7u15kWdItijKV7deq/SkxsZGIWPVHRSsLUabg/Fo1rvhQSVK0lJmlSqKs086OaDX5oDvIn5bIUUi4QNizOWSrkeMIlfRD+pWJnO/Xa+aIN8lGc1isVdvj9fDrsj+S1aHdZIhjRS1ULL9xvPb20laLEoQikljxhEI/aUV/vCCPgBm9R8g41UW5oeOIuiGAtCR6MFbq/EIiu7daG60V7kuvA6aIn4jMfM89SDgoiQ97KzlRaGpfiONqKGFoRq1CGCiBGjrS6BJhz//zEvgUpaucD5FCRinMmj50o44/o7wXNNRAcyFiXo37FhLz1gtvv64j4Ag4Ao6AI+AIOAKOgCOwLgi4YLEusPpFHQFHwBHYdARGCXgj6yHsIWgRKCDgn5CZRwb/22p5yBjIMI5B/tQ5LZrQU9dUMZHuENiEAYKIh8Q2IYB8BdxvIbQOHwntA4+H/e95NuTn94XW/ukQK9z45Av3hFgJtMvsi2HP7YdC+xBEoOXkgBhktT7lxDvEQklRRwhqCEvLgcH7rOJH2KDenAMRT10NLz6/VLAAN85BrOC82vuhwcUIdq7Ja8SNLIhF1l4rrHcdDMPevNbvZiE/V0qAmVNIqDxMv7wXbv3JVEnCnwpP/Ed5XpxGwMEThs+BCdehjMdkxNT/c2H4EYkW1GnDtkao4H7mTUGZIAPpK5bUFmKY46wsJ2E5K9IRJRAHIG/ZU24IYwQOvGvwSmGDgAXXl8s+0VyTnCZrtX1AF/qcDJIXEp6+Zu1vXkQ1oXw9/XutCnu115FgoVA2CrCfxEm3n88qMTOvezoo7xbl1C6KC8ppIceLeEYrx/cUVTkhEWM46OZql0pOFXFL8oTyJFSndVyfL2nLXSJvDyqMzlD/5/Ky2IrELOPUVsPbHGf98e/qva+XMQ8R2gkRjT5Hv1jNBkaEGiNUFHvEBsbE78gQgm3OLCVWrOS1Mzo/Q6yT7LkOXyfsVV6Ic6mEUYzHkQmwjC28yxhLhFtDIKQsn5d4AYnOWON/6vlV990hORDMI5D9cWFJ+16MomqPcmjfppwVe8phNZNHpdo60hym5NpSk5tvQVyNSHGuHBax5t/qrHzcgvJXKKIa8bmUqPvSdwPzRZ2gfjWd5VrOUXvyMfotW32fHdJ+1wKXf8YRcAQcAUfAEXAEHAFHYBsi4ILFNmxUr5Ij4AjsTARWSsoN4UFc7gYViBZbjQuhR84AiHwIcv6H+GJDpMD4nHkXXBOwItoh135EZvHdLdE3hNvJkO66M+x9564w89JB6D99TP9LrDh4Wl4IuvPpJGRHnwrtw4S5uUPcEtcazZvANfguM88RBIlLHg+XCElIalb4Uy+8GCDIORdSESKI0C1c01Zic23bjDDimogJJkrYynMTNiAKjSizlelGaJUh63QlWChu+uG+CLB+SKY7YeZVyrmR7AlT8saYOP5sePzn7gvz91EG6kMuj9tlrBKn7LQB3havEJb/RqIFYU42chv9rQAWiA70CQvhZZ4qlkib8hIeinNIVs5xiFfCXuFhA/ZgRlt8RHaPDI8XS859ubpB2hLi53Ibghb3JKE3oZ8QLGhrVsEj2HEfy11hIcfWjXy8Qlmv++0sTfoKZ3O62x8+rddKDB9NV3k52esPci3Jn1Gy7dawLDuJlozjjVGUhTwugpTARK+rljwrjg4GRVed/QmJHxeU/+IxjbWevCyYF+rQN1tBtLhMjou6bZXjwjwv/lD//mlTt7dpT9/8cRmCAaLjd8jIr2PbCb14n4z5ACHuF2X0Q/oy10Y0pU8zl3IPwj9dtj8R/kekdC0Ey5iDGGOMf8rANVpylmEMIYQw5pjP6M/MXcxjiHyEO3tY9kkZoe2YM8jPwlxEWRhjNqcThqrYAXkvbG6m7pdyWDAXVdUhhYLaXxUSKvRlqO/Kofq6dDxlrYhKeSQpqYVi+sWaqKM0rpScW7leklYZlY9JBEwIE6Xr7FGjWlg5E/R1i7XfECca0YJ+9DzhYu3v5ld0BByB7YbAK1/3ncwb/DZjj5mnn/3GHV2kU33qo+/fsr+BtlvbeX0cAUfAEXAE/hoBFyy8NzgCjoAjsAMQsNXj4mp4aGEFLg8tkGUQbRBldYiL5hhEpZFd9lBz1Sg1ibVJessKYUg4yDMINwzipxdu+C4F4jg6q+TV8kLopWHunmfD5AuyEE+qPOnZMPs6Vj8TEgUCjhX6lJnPQ0ZB+NlqYrwoSLgLwWcPZIgMPKhB7hkxbeE8bJU9ZKWtmuVzRnjZqmzqDQbmpUHoLBM3jEiCZOQ15WJjxbQJPhyblNCiRN3xad0Jsl0eJKp/tXhRYa4UKupvzypc1EvDIz/5uXD2T1j5DhkKGQkxyeptazMw/F7h+ufaf2y9E3I33hVgglFHcAR3jD5Ce0CS/pUMAg+RAHIVTwneQ4ig7Ig4EK6cw+doJ469SfYu2eU28l2Qj8S2y4kVrD4/IYPYhey1fAbgyb1pewsLRV98biX6VvSLrPkRAAAgAElEQVSuMEDmF3rFRLu1KHHihISL/XKc6LdbSX5xcYg40RHxPej3B4uSKTpRERWsFi+qSOGfhqk6rTQO4vZfGh9q80Na2f+0hIyLEizsNyI4rWm8/iu0+bq83YRmWpBwwRimbvSJ35UhYDF+mQPpv+Sh+JCMuYc+Q19G1KTv/lcZ44+5hX7PBjZmYSWxoiGgR+vGZ7gv+Jp4Qb/EuBfzEt5WzD+ENCOsFf3avMRqYUP2yuY4YxRPEfo9wqcRUHgX8fqiyvCIyHA+tx036mieb2AAfkfUn+/QG4irpxMJ3voC6SdROC9rl9Lw9AlpdBXJ5qUnV61IMaHiJC7SNMj7KO6S00Vj4VkpH6d1CmIxc/Ka53ZZpn9Y+42KFuvWbhIlR69t3212rFL4q3W7t1/YEXAErh0BiRP8RuO7wIQJ9nxPsGiH3/IWwpQFG/z2thCweMXym2he16jF9pHvjecVSILGtRfQP+kIOAKOgCPgCFwjAi5YXCNw/jFHwBFwBLYiAg0xm19aZKrgF5c8L0yUsDwDJl4YeX/V4XJEqkOevVXGCmZeQ/LzsIRAAtF3W7jhe28Ls3e/ImSHJ0L7SKywSOdCcaYbkpm/Ci2FhkpnIbNJ1myEHuXje4sHM8rMax64LLSPiQoQSrYqGXKdhzMe2BA9eICznBSWnBXyHDKe+pqnBM27dGUr71uoJnufclg4LSOWzCsCTwl7H+8CCP1LHh5pNgzF5CCUE6pTLwuzr9od7vi/Xx0e/d+eDad+44UKicV5dQx2mRH9iAOQmRCs08L4QxItqNt6bmBN21GnYzL+hwwFX+rG/7QvGJJkmHBQtAOrziFXj8pGPVvAkFwVEL6r2ZbLMQEGeG7QN/5Exv/cD5KSstDmELysXAdH+g978zLiuHkabelVhQ+ceLbav2cq5HmVtrIka7XkTpFlNyqRthaGV48uLg4uKHVFTwTsnnaa7iWRc14UqcLbzBdFpehRyn8Rx4v9YbFYFMVAxxYlVmQiZkdzlqymnbbMOY2gMJRwwbhFPEPQoo8ztk2YGRVxIXToP4gXJvLW/cbECV2L19eycR2uaUS7zcUcw1OIPs298eagn+NBwfZhGf2c/o4hwFJ+BD3OY2NOY1xaCCnmDcYd1912G/kkRLqDH32X74VJ9eMTEhpuuvRlJ50uVH3FfNolhwl5VES9pKo68p0o4yrovbhQ/KeuvCqqYb8qpOwp/0t1s0JG4XG0qNdPNaIFc64J4GuG4xVCPm3EPGXfd0v31NGwrV8vV2kXNNasK/iFdigCEg34rYeVEggQGp7bGo8J/rfxyXkmRPBby0Kc8juH7w+ECb4X+C3EdwW/l/me4ffZ18hYCMLCmA/KPirje4YwsfZ7yXLZBbwvuL97YezQjunVdgQcAUdgExFwwWITwfdbOwKOgCOwWQjYivJGtIB84SHIVt4+t7LzWlaei0iHMEKoIHwKD0ysToYU5GHprtA6tC/MvrqlZNpJ2PWG6TA8q2D73Ysh2/PlsO/dc/JGOK7zXiuzFWOIHJD9PJzxmj0PYFyPMD/mcUG5qQMPcogWvMe1OA8CC+8LI+8g4Hkg41xe84DHd+LoylITIMwbZVTAsPc4Zg+ClIv7c28IdepvuR64PudCelKWXAnDz6gmk6FSou681w39k6fC1Ms64VCrEx5/nzjlAeIKBCTCBd4D1J3/WeULWZ8I69+UaLGeq9/BB4HC4uOTL8QefiFGeTi+V8ZD7qdkhNrBs4LzP9vUGXEDXCg3dcHrBhyuFN4JgUlxwb5qg0ym/mycgwAGVpSHtoTkxTODB/WbZbQVJC3vQzZaW9QXuJY+vkyZNuUQJO2/++3PF1kW95JUgfez7MmsJU8e1biVJvd14+jOyXZyJC/TtlIJD/rD4URZlLli9A8nWklXIfqntYCcNBgQuItlVdZJ7EXMnhLZW8MjGw2Ttin1XM1Nl6xQ/6oV4ksJ4RFPCOa/eYkOFiZutN6gUItrnK9zoiuFe1qprJchpGuRQuWvy0y4KPqo/scrifFEvhf6MWOPMWOeBJQXG90+rX+YN5l3IKZM3GXcIdTVyRG28QY2l3IiXbKn1I/Vp6M3KDQa3nT3aRzcqrwUU3FVtodl2K/wT/X5EjMKKfmZ3g8KmaYt6ikj92Jc5mcl6p3LQ8n8pfmjwrtiWyU5l9BjYWMshIz9Bog7bTTNqMySpDx/sVfX25ONb+MR5FXbcAQaMYLfp+btW+oYv5tYsGG/7/idy+9gvqOZ3xEc+G3NawRtvseY5xm7LB5BsEakfqPsPfqhk2uQkxqJRSX8hrPtzXrx6zKO/2cZeZnqvEoyFt0sqCycG2vP7zrmCpv/nhMv3QNjBFF/6Qg4Ao6AI7BmCLhgsWZQ+oUcAUfAEdiaCDSELd4WzyP5roPI/XYhAaHMCi9IIh6OII86Icomw/5v7Eq0WAhz9x4NRf+p0DpysxJsnwnZXoh8HpAgkCDbeDiCcIMwhDhnFRkPbZDP9qDGPTgfUpUHNAg5Huogp+v4+801ILEpiyWM5oGLz1Hnh2UIGyZCPCfYNO/zPyKEJV3Vy+d5Yphnhnl6jMaX59qIDJQF0hHSizIek/FAelICTRayydkw98ZbwsTh82F47+EQTVbhsf/rL5UTlnuS+4PvazC0HB1cj/dYVfdLFGgtt5Fk21Y3cKbc1MdW9bEajzaiTJSHPSIROCBKsNF2xBqh/chXYQ+6hNVh+6GmDggJPCjT/rQ5K/+OjdSJut8nw1MF8YOwU6we55qsDqT9uQb9g8/zwM1nKC91sNBaXNJWseNmtBErl0eqsfYv73npTcWDJ073Jjrp2XY7VUbt/DF5TOwSMzGTZvGFwbA6PJTrhNhYuVMIKKUQFjnb0m6QD+VRUSgwTlUpfFSZ0u5aSQ4oCD+MIUu2XiffbrB7rhJjuqrayNfniY8SAKpGDFi2EZYIEbVosPTElcSKa/SueN7lR8vWiBcW/g4yir6MeDc6hpZ+nv9pI1uZu1TMWPvON2ZXbLwsmIuouwltFzTilctG4Z9CdFqD/kwSV5pjo5t0XIJxUIoXxYWSspEkcV9OSIOoigt9+FFl436oipPHFEnx80L2aY0V5hzz1Bqz2l9XcRgr5smXp2ncVhisaXlqzadJkijEXKb/y+nJFnPCQHPB0EWL68LbP+wIjCLAbzwTovmtx28s5i8WizDm+J/QhIgP5OTCa5XfrObRym9sfp/x+1LTVnSXftu8Rfu7o0gfrQqlTMuUtSoL+aCnTD31V/mXtOd3Fr+X+M3Odpfsd2SIFdyTRSj8hmLO43++W/htdULGbz1+i63ngpmmWL5zBBwBR8AR2KkIuGCxU1ve6+0IOAKOwBIE1oK81Yr/t+uyrPxCfIDANhLkFfXDT+vAYmgfOhjSg50wcetsGDzzRJi47VyIE8h3Hpze0+ztYYjr8DBnMdkhpSFT2UxgsFVpEHwQ+Ebu83AF0cdDHGKBrVYz4pXzIN15j2tYuBfKwms+C0FFGbgv1+M151IvKwN7CB/Kw/3ZUxce/ljhBjmPiGEeHYgxPITygGmJyBUKK50OrdvKkJw+Eg5/Xye09nXC/GfPhzMfmg/5Wc4nVj3XpWzmtXA3mMvL4vea8qzlDnyoCw+vPBBbvpM6ZEFTZzxW8KSw3BIIVQ/J3iQDK+pquSPAkBXihLXBM+J1MvCyVXuE52EVOPU8tqQitMP7mvfBgjblIRpvCzA5IUOMsjwikJbcj3OtvHW7r0U/X1K2Tf0XovsDH30473bzi0qe3RoW5SmRi93hsJge5mVXZGtPDhRRqyUaNoq7CnbTUej+C3mRnwpRMaE8F2S2WcxLXlQD9WTpGTVmECYQEiYAbGo9V3Hz0VXiFtrNPERq77FGCLiscLGK+2zEKSaqMa4RapkPmfditfdzQorqY6S8nb8RZRvre4yIFnV4FfXpTGIc89e89MmhdIlHlVW710rjqUKKsGJBzSl5C9m5FTlNjkYaA5L3iqiMzsgV6UmJFBc0NM5J87O8N9uGoGs8K2hPGycSJ9K2vK4OyKtiVnPl+f4glxdW0ZpoZ/N5Xp4mPNau2U5Pn63JShcuxno4eOHGHAF5LfB70gRy9vxWRKS2UJuWs+ilOvZajT9+Ux1nwtJKg7txCNMiBMLdTejIS5WA53gstzGGdNJqhaytrw2dm2SZkvUUoXvuWe3rtTpSMHTjMq8FjEselRXzJL/BbcNblrCb5qnHnMqikvc15eM3teVs2/KLP8a8q3jxHAFHwBHYkQi4YLEjm90r7Qg4Ao7A2iIg0hzi+J/KeKBh1Rcu6ZBskG2W6Hoq3P7Th8LknYmekM7Jy6IfJm+HYOaBjYc0yGpWc0HIQT5D0JmHAgQ1/3MfSHLLoWC5CGxVGhWDrIYsR3jAs4IyEVqFa0KUszoN8olrQbTzoEUZIOaN3Oa6EN4WSognPK4JscP18RxgxRubkYV1IJGRY0b6EjKJcrAyjvtSfjwF8BIhIS57rq8wUekXQ3Lw7hBPnwkHvlU1eFUcdr9lX3j6l46Ecx+1RIncgoTAYEdei0j4Q/7/hIQLi18/UpTremnhsNhzP8oKbogStNkxGYIDHhi22o8HWtoKvNiDMR4OtCHl02rnWiQyLwweksETD5ijMtoWUhAhxPKLgN8jso839+E87muCipHVPEDTZrZC8Xn5WLabWKF62lYqOXA3L6KLWh193yAvFgfD4mtFOh4WFZtFSbSg5NqFmI1FiRoK2F9cVK6Kx/v9AuwVGacS6RAhJp0RwQuudZikZl/373EgJpdJTGz1p3/aKnGIHgtzZ/MCY5utzmWi69Ti1eU8Lkaw3cyX9OX/Lvt7Msb451X2j1Fu7ann35QhfH5C/zOGnkcaXSEvwmbWa13vTcimhoyvvawQ4tQ5JkTc1SSgBAiR8KL45F1BuCO5HfV0TiJiXjkuojN6h2FyUYTgOTkWPCZQaQcE23wcxsEag2die0tY7Ms0UaSJgsZF8Wn92d0fDHdr3tit0TWUV1ZHOOXywjrTytJnB8O8i+fVNsRkjSH2yzkCKyLAdzDfS/xeIkQlv69eLc/bG/T641pN8CrN6ryn7+dqd5Skr0xbnQe17xbDwYs1Tl+WtjvyXpbiGifzcZLW4U3zQT+0pmZC1rm0vkdznu4yqI+lmU5Pklv1+VAM+xIw8lDI84L/6/OaeJD6GMLJN8jwfv0jGb+7+K1HyFbmQ8r9Rcom4YXvH+69rHDhIaN8BDgCjoAj4AhcCwIuWFwLav4ZR8ARcAQcgecQEFnOiq8flkE4Q3LywAKxzQMNRDWixRPh2I/eGIYXJ5SzIgqzr/uIlnxBgPNw9jIZhCPu6XwvQZh+UsaTFrkJWMEFAc0qLwhvHt4govg8ooDF3bYQMFzLVsGyRyCALOfBECLzhAzy++tkkH2UmetY6CVbwUzZuDfvs/ofoYOHMsQGxA+uiSgCKW5eH7bi2QhUCHRIMkh4Eh1C5hPOiGtzDch8ymjJsxEgkpBOLYb4eCt0v7InRGkU9r9nT8gV0/7i52y1NZibaAMOHP9Haov/U6IFZb6uTQ/KxDo2kQK88RQBf/NwoZyQeBwzUQcBB2EBscqSc4MbRCvtRV154KXseJ/QP8CO8v6qzMJ88QBMfSCZf1sG7idkiFe0ISIPG+1Of6DduQ7txGYxnpt/Q7GNhYq6jt/6ulvK//B7X6pjWE/GLfB4THX+Qr2wMo6f1croThnFu7WSUnGgcvGwwo6Y1rFWked1ku0Lau/TMrBjzFp+Esv5Mc6rJ0dDQPF6Qqvi5WhSdZWIfEbeJuJXq0JvJKpEC+8TDnVa6UAkfzGOogVCQyPOWDgz5hnmyX8gw2OL/s5cyTjBq+2dsp+SnZA911ZcY6eKFsLB5lX6xFmBcr+IuJs1Lg6ov0ug0JweRdMi6Z+QSPFYr59nEio6Wq8MtoqbUj2imeUBjR3mecYEYZC2jXeFTY5Nf1E0rGhSySqmW61kuHtmmnE/eW5+8QVFEd+VpXFfc8OMyNFbJYg+qf+fnOy0evLKUjitCnGIvB7jPEeMVNdfOgKbj4AIfn5f8duQxRt9zUW3R3FQwphEr5N3JGnrZnlL7JOI8Ha5fk3ESfarEhOyOM3uaHWmF8p8cG/WnniB/pf2kGm60tQURTP6X/6USWhPa9qL9TWvi0dK4IMQkcrjIo5n6/+T1oTWDcnHTIZg0Zs/G+JsGPJ+l2w+jddFvVaBEKssLuG3L2Xlu4jwhPxO4zcHcyNhP/EGfLCeO1cQLTYfdS+BI+AIOAKOwFZDwAWLrdZiXl5HwBFwBMYIgUaseK+KZA9frLgyrwlWZ0Fsfz7EkzeH6RdPhKm7TobpuyFDXi5jRTciBw9tENo8+LC3+LmWHJk9BD/nGWnO/SCWzFUdVMzTgfdshT0EE+QrhPiLmvIgYLy5uR+CiCWR5lwIdwh1rn1Chihg+S8QNxBVKKcl2uZ5kAc4HtIsHBHlsFWrrEbjXMpJmXj4Q9yArLck0BYSgHtxbcozo4fNU2HvOwZhePpQWPjiTeHCX/RC2X8sLN5PGagj5eGeGNhw7L1qk19eC9FC16ItKSOeMpYfhHvRHmBEO5LkF6w4h8yMvPcVGQ+21BFhiFjLiEEQq3i4YIgLeEvwmnMRK8CG9sCz4oQMoeSNMvCkr/CeJXAHJwvbZX2A8phgRJnq/rDdxQrVsd7+3tvvLCRahHaWSHwQOV9W96sXlqr/nBJyz4rAv9AbDHcpTFQhAqQXV9UFBYFSPy3B79nGswIM6/BJ2sCQ15AS405GMt6oh6JelKVWz093ewPlUG5F8jRJulomPjXRUlz+MKF6DkW4hvmFfh3ySqR+Xb9xFC5G2oHxzbzxzTI82RACGV+Mge9uzsPbAiIJ76fniPWdKlogLohIp41pX/oxieSZi8HsCXJWSLk7nJchk3D3OHHQdGiiKspdeinvgvCYOEATrJkHIeYbqJ+/G9NcLsuW1Q42HigmSiN8IaAfWlgcvFzC5tlOJ9P3WnSzRIw7NPj7mk+GCqm1T4KF+hZB8cP+llwx5M21cMP+Gb63vyrny2UL4G86AjsMgUakYMzxG4/fUHdoUcHtaTs6p/3bNP+8Kk6q2XQiuymUsUSDcDDJJqclVoQiH36XvrNbEleDxIoXy5NCukYqEaItoaGl4UgUKP3VxFV/Xet1LWJoWpPwEUncuIS27XmdXHIKRrSof7CqALwe9vuhv3C29rogv0/jcfEunWK5wLjJCRm/QQnXyvzB9xO/D5lrfS7YYX3bq+sIOAKOwHoh4ILFeiHr13UEHAFHYGcgQLgjyExW0fOgAnnPgxhPRzwNPSKxoh8Ofc8g7HrL4dA+APEDWc05POSw4p7/LYwPBDYEEw88ENlcG+Ka/zmPBz0MAo+N4xaKyUhVjpmHA/dg1dfflfGdh4cDIgJeEhCyiAQWYorr2L1I8Exd7m+uTwgm3qN8EKOUm/pC1OM5wIMaz3xGFJpgAdFvsc9NUMETgdVqJIvmOrjXc23KjEcG5eM6fPajSka+GFo3zISbfuhAeOoDU6EaPhW6D4Ef5TORhM/SBv9FRpuQOHEtNtoCMYY6IBjQBuY1Qv0hTqkX4hR1Am/KYsm3+d/yftBmCBzUmzpbe/E+90GUwFi5h2hlCdJpF8shYr9bTDSiDJxLm1sYIMN53En2tWif510D0UL5LEQulqeVRviiuIdntIJ8z2J3eEhgTIu3v0Gx+EMi8lFhXp4i5zjUo96DmLVY1OzB1UI+jHPIF/OuSCTEtAaDXCtU40mF9jkooeLAoOi1yqJMpF3cMBxWUZZGWmSaFjp3kRXjEnPmz8/3FuZmOkWT32LFFfQb7akw4mUBKfSLsu+QMa++TWX9hWb8EF/cNsRf5jqEw19r2nDN+9gWuyBzgHlf8XpG7T4lLk+eN8wbdSi0GRGBhzUbETZqQZzd49o/rP8fl/cAY2FBgoSJeFus+lcsrgn7UyI45xT6PhUhevMgL+8qF4eK+hR3ZbjbZTpeKv82ovJdUoH3SKiYrYrq01mWnLxwsd/30FBXxNpP2OYISJBYrobm+cvvRn5v8ruO34AtzUMv0q/Gd6Wt6O6JuehwV79qFL4x7D+q7+hWmS+eSybnn9W0xQoEfXNFrY7WsVxKn5ZOaMhqj0ARx5fSjUmYqN/THMdCDd6z78fLIs/nskmmRoWDLAtlsZlMpIqEQkLIoLugUFH1+g+Sedf5fuqbhfBW2cMy5kh+k/ObjgLw25nfi/we880RcAQcAUfAEbguBFywuC74/MOOgCPgCOxcBLSSHzdxVs0T3oenKAgzSGtWWu0Oky8swty9nwiTx+8Ke971dEj38J3DgwyeDmw8uEHAIQJAOPNUBPmPOIAXAYQ1ZLZ5LEDQ89pW0fMwZuGguJ6dZ+9zDDKbh0OOcX8eGNkoL2WBjLdE2ZBSnMdqUa77PhmkLYIGHgIIAeZNQVktrwb34HNck+MmIpiAYTH1TUgBH66DSEPoK3Cw+r5Ar3n4gxiibC+RnQvtm0s9LD4UDnzLsZDNfiI8/csvDotfoT514lMZq9wQCb5F9nm1zXl5WXxMr695a8JC1bH+m/tQR9rLMKR+iCuIEmDMyu4vyPCwQBCiDoSHoj6cw+dIco7XBWIU1+J/2ptj4MNnEEV4CEYsAjs+CxacS3l4EKaNKI8JFTygb8dwLari1W2EhxKhPXjgxLPFE6fmiYkNMXtB+ymRjs8oNlJLgkasYBDPECFKMfrpj+Br4dwQpMAYG2exwoChH7REpBDeR2F9yikJFO3zF/tZpyU6NQ17BoNyTrlHVb9q2B/mrelOdlor61vK+3FKoaFSnb+ovc1B49aPKBdCH3HEmQ/eIftFCRpdtTP5YDj2EVkdA13b+2XMDYgcNWm0E7wsVvB+YO6yfCyW30eJ6AlxV9Hvnxav91BZ1d9dbJqTq6f0/5Oa9Sxk3XZeLcwcrpwVsfKLR5rLoxl5UJyVqHlI5GULvlNqxaT+zqIEEmJO780LvzLLooFi0czp2MJEJ+svdJX1w0lKm5N87wiAAN9NzMv8JrTfuxzj994xxWv8scndVditTFOtqeQZRYPak7XLbnu6yvuLE7vyflSHaEozeVIoTUWqME6EfEI0YI8HhTyf6r3ECea5mteRl8S8vC+439Vs/IZSrKh0qAJGcbsd67dBLZDIu6PxV63DhNrGYhvmTX7jYXhgfKPsv8nwnuW34AXlrthxC0euBnQ/1xFwBBwBR+DyCLhg4T3EEXAEHAFH4KoRECH+N/QhwirdIkOk4AGFnBCDkO76Upg4flto39ANsy9LFQbqcSXa3qMHIYhA8jhY3gIIfowHK0hrvpN4AOIcNo6zkh5y35Lncg0j6i08EUQUZLh5NfCAxIp880DggRFindX73O+YjCTcCC4WjgmyHXKcc0xoeL1e45Fxj8zyNeC58CoZZJbln+BB0R7kKBv3trBYdi3uA6HD++ZBQv0I8WK5G6ibeYawGo/zLuWISLIjITt0KpTdkxItbg0TelZ8+CceD92HeVDE84FV2B+UIarQJt+qNtov0YKHx+vZKAP1QVCgLGBk4WnA0rwZECnYSJwOEUh9McQKhIcTzXHEH3BDcLDE6rQ9XhW0PfjQP3gPLGgPQnJx3JJAm1DBeSao+ENx0wDs/n/23gTKkuus87yxvS1f7pWVVaUqVaokWbJkW1iWbMurjKGNbcA00Bgw2AxLT3MahmFg6GGG3qabM8yZ5tD0YYYDNOthaWCapQcMpjHGNjTGlm3ZSEaWtVSpVHtmVm5vjRcR8/+9el85lKpdci2ZN07dei/j3bjLd5e43/f/Ftwb4VdebpAkn88Uw8NJ9OEGuIOCrvqvX8jKQBrkZLdA83y3gNsAYdcdTTdbOZSCcEuYGlR7/cHERieVFZKbaHfTnbKyqMprTa3Xz2qiwQ65iurK4mIsmG4Q1KLT7w52yYVUUKsmHRWQKOYFMS2uN8CCcWEf/Dml/360LljzT9NW0eARhlwJ8GLk92MItrL//azSVha4l2b9eb8yjw3oZA/h+1krPNSKR3uLuYsCsGMdDN2hEcD7Uiq5gfMoxHbQIUWh21VN4moW5TvkQm4mTbHHGsa4qRDjQ/hFIbOLlraUnXEsL/mSp8oD22cVfHugmBa4zNrYBvS6gYfaN/1LSQECS8vKwqwa2E84x2CJ0NP6SrXVcE7F2vcr5KXJTeyquPnbMjcxnxYyaJgWOBCNTXeavXbXVeoDeWyKBUaEri31jbQ7UGq72vjU0JJCvg8FJihGhdkXj8AK+qcYFSjRXO5l7uF0QhBuESZFHvaDSqM5BEQGcg9VCsZ9puwgQFEAt68ozMAHoIyEW8K/UMIKkPMnZ2V/eQp4CngKeAp4ClwRBcxM8Yoe9g95CngKeAp4Cmw/CkgQ/nb1GssKBO4vV4JlQng87sZe0XWzb6265t2Zq9627sbvRDnzWdmvo3FPPhg4mClcCPFpgiHeRwiuERbdo4Rw3CwoEHpzIYwzKwoDJ8wNkMWUMOEUf1M2z/CJ0B1LjoVRO/gdQThgB+ACQiyE7mj4cx/tMIs5cVDfYcRoB8IrNP4BGcxlEYLBsiso2ko7EDKWLUS4T7vNkoO6ERbTNvqBmycE+lgfGG1oO2Uj9J92WW/NdZ864dqPTcst1Iw7+BNtly7SF7NMoDza+HdKgBgfEGjxgtxDjYJvw8zST+gJvbCoMAsK7sG08jsACnMBrW+Eg8wRAIpPj9rDswAaCFl5rgxWGa0MHKL9WI1wmTDRhOgGlGBBMMriPzZTYOSnHtoZ2GTxTphvzD9bZ/zNnGPszB99cb0H0h25cQql3T0mMGJvp5veotgUE9UkdK1O+rK2AIx6EqMQXi3yINJCGkgI255sVo7EcXxc+qSdZr3yjDIcrlXjgbTLO7K0gA7EtLiugAv1lXX07aO1xWUdpEYAACAASURBVB7yT9RG9gcsKFgEBOXGEqN8sS5xE7Wdg28P6TFaC+zprAf2HvZK9nRzizSMZTJaF+zJPc3/LevWpBTDoi6gblJWFrfIHumVSq+VBdYrRYiqQIv+IC0aAj1THMcpX16N5H1NP0qm2ReAcUj7738TrPEJWSk9pvW3KJqxh/jLU2DbUWAEVrCvcDbiXXuTDihfIeOkPUIRXiXTh/uGDhh1pJuSk8a5AxVXaShwzmRf+jyJQIjIzd2y7nrtoLV2Immtnoh3ci/rJW715JjiSUzKyqI5BCq0RnMBE2WLhzP0LorP6sw2o99kRXbll6w0+oNuJxikvSgb9MNUrqHSDtjDmSM4gbqJozEM3F3IseSZH0wRFsth3ju/o/Rn7Kne0uLKx8I/6SngKeApsJ0p4Ln87Tz6vu+eAp4CngKXSQGBFa/WIz+khMUCQh1cGHVcbd9jbufX3efm3l1xnS/0Xf320MXTH3HNuzB9Jx9CoduV0M5HSGTxGhCOmksa064nLgLa9uRBaMjvgAS8sxBgI9hHYGeBrHHNRPnkQ8BkOmcGMFAObSiDCjyLsO/wqCwE55QNYABXRluwrgCQMasO7gNcAGZgdYFgE405mFPTwi0zkLQXoT0XTKxZTFA3l7nPsn5yn3KoB2bXglkjWIb5/OTo/opLT8y6xT8dd8d/dd0tf4h2QlusFAB7EMYBHEBrwJefFGjx8VGdl/1RAixMY5A+Q1vaSB+YC9AD+kNDgBru0S7Gl34hSOU+muEAG/g+ZpwAPsgDbcy9lXHF5oqq3Obnaf17wOLCQ1oSTJpFE/OCsQQQMusK5hrzlc+UgMWXPVGu0QMS1keKQzEt9zUEDN61vNLe0Wgk+6XAelurM9g5GLB+sx6yHQle52RV0h9rVHtxHLQU1+ITjXpFYFq+LA3x1Xot7kRR2BJoMQwcej0F4lY/WV8/rPQ+JayocMHx/hLZGT/Azv9F6Z+M7v87ff4zpfxqx+C4RtPhgtWO1gJ0Yv6bm0Czshs6amfcodd2sRQQTZIkjvZqeeyVa6fbRJx3DPL8zrwImpKthrKgqOgd0NY+G1XlYA23UPKQn+leRwZaG3ESPqy19sHBIP+4LLgOCTzsX+9A59WYm6O5Vq6K+TYE2j19rsYIXN06RgG12Vc4qz6ohAJMJGuIb01qjTdGSfUVAhn0lt04FIbZ/ltf23PTewu5fIpcdaxwYzNYMcT9+kSaKvD2+vqpaO1zH2wmjenOvom5It5YarrTx+YFDoxnYVjRnlVovwrOBLQoig8LGGHv571glyn3XCkhTudZ+tCg15rIer1b86xXT3udsUFfL1SBFblerEPgZOiWanhcUBCNINUNc7MKLbBk/kYlzoW5QIsb5lxxpUTzz3kKeAp4CngKvLgU8C6hXlx6+tI8BTwFPAW2LAUEViBs/l4lLAss+PRTrn7rgpv9mle6iVenrvfMuKsosHbzpSuKWQHzhEAaZoXvCKJNEwtmyrS+EV4j/L9VCSE4gATMvQEPZbc/1E0ZCF0NJEDQhOCc8sgL44YQHME9gvByYGoLBg4IwPMAIx9SwuLDLCzQ9Of5B5UQXMIUwoQdUEIID0MKILAw+p22m+YuZZplB32gnbQJ4TB1A5ycYTLP0NFcRtEe3sn2iZUB5RI7g9gNBhK8TN8PumT+mJv7+l1u4r497vH/cdYt//lndR8aUyfurSgHgIC2fq/G7hmBFrhruuxrFMuC5yx2BG22mB2AD/QH4IcL+hhQhFWIBVi38WIuQFuL6wGgYi68jJk1l1nW1iGNPDBx4aE7jw9/HjKrI3OhZa7HzOc89DWa3wgxK84SYmRZQMDtot3tpwIj5PopEEhR3Jnmxf7eIG9ImCJXN9FGHEc1CVWnlHVDFOl1u4PJdi/dm+XZkYlGvSbBC6YYS7LAWBVgcT0KVtg7cLXBXvNtSl+nhPaqWQEwzoC9/1Lpu5XYTwA4yMNzW9210YUXiH4dCYpxl2YAHft7WXlrOO7bRaD8RTCzAJuIZSkhx/iuqvU0JYCvK8rIc00g5zPSoNYC0dqpDmNbuEKuoAJ5kFLuOJwRqHFzlrvH9RzvKgN+LjoeWzFDCRSje1GjluByq5hoVobKDHI/5/7w488M5K6vWFphSbv83W88cD3uN1txeF5wn84TWJux5TzHeeulSu/QmD+iOBJv1Oc7BFi4uFpX8Gq5eqpF+3fopFZtRvL0OZDrp7w3Np0H43ODuMjTKIgKQMFafWIw25gerG+ccq24WsRjM4NBlBRPry9W9qS9ZIcMG5a1Dk8KJJD1huKVFcUOfT8zj4pCRlAFbt70DiBxq8AaijPywkWIYOeDw1Ecr0XxWC+ayuUxMSrCuH3P6vFGdSCLj97G2hCoUD3aHYbbQ6C/Kd8UcqjmHrXpbUNA5Yy70KFFoL88BTwFPAU8BTwFLpUCHrC4VEr5fJ4CngKeAp4CBHtFII2QB0H/Djfz1tA1Xzbjpr98VUGgq276LWsurEnQMYagGgE9QncE6QiF8HNbfu8ghEdgjZWGCbEBHkyQiuADywcsGMwFFIJ489POPSwiAA8APbCGoD6eQajHd6uPTxPc0n5ADBLWGbhSgZkCqAC4wN0TAIMBKgj+ARAAAgBD0HQmvwkACRANsEB7Ed7TPtOmNG1ec2tF20xABmNo7ki4T9/M2oLPoWsaJawr+JvYHpQPvRbFh37W9U/Nun0/0FRg83vcsz//8Kgd5DWgCLpAY8buV5Su6BoFtM7F9AI6WYBm2mzxSKCNaSrTP+hDvdDaAmSb2yGzguFZc8NitLRxPmtJgbDnihq9zR6SkPVCPR5qjkuYxpwz//1luqL1e0MKtOWGJpQP/aomTk2gxGSlko8lUSjJTdBNhGDEUdxBsKLJW5NauISy2fhGp18o4Km8RUkBNgxixRXVegoP67GPx1HEWrVYHtfT3DNAgrXNfvSPlH5KCcsqu8jDHvqjSv/X6CaAxcsJ0H09WYxcy+VpwMW1bMN1VLc0o8OOrCQqejNJRhkIdwjacl2j/Vl2F4GTM3v28aKWawFp/cgVTSAhvMu0eNIw1L3U7dG7YZ+e4XzQ0z6zLa0ISm7HIsX6UJxyVxGdGnKlFYqGsUCdJKy5TFYovBM7lUqU9ft5LgAjvXn3lL0Lzzk1vIXUtV8x5wArTHmDsyRnwFcp7dOZ5T1hXHFJXW6chq6TEgEWDYETDQEVsatPLbr1U7NFFLdak7vaq7XxbDIICXL/xT4S/ro+kadJ1T0pwGJQWw0EqGfZ2MzKqaVD4XJrZYxzKHu93lfBu7ROcf93pgSAibzoCUQ4rYDZKI7Ie1OiNR1hlXexa6gbEkbZSxXNZk5r+nhzNlfIp6xda6YfaEwmb1o6XJ2K4lnXXV8dxrbgAVldnavcRHd/FMsL7Q9/IPpxRjQFpLP5if3hL08BTwFPAU8BT4FzUcADFn5eeAp4CngKeApclALS0P8BZXqzElpkCJrX3a53t9z8e6bExyQuaqZu8rU7xTT9last7HFRFXCCuAX7lcz9Bs8hbEMYCFiBQB4BPEwWYAEgh1lWUA/Cce4bk8PzCBMNiDArCQAGyoSBwwqC59DgRyiAAA8AAWEs1gBc5gYHDstiUfAM93mOC5dGlEl9lMvzWBHwN4IF2gXYwX1ADkALnre+wpSZ8J1P+gBTaywp7TJwgvrok/1uLqkAhSwOhIEh5CXfm8XOrriJ1550/cOnNQYLrvNM7pb+lHxYW2ANQ18Ai2Bk79YYTsrK4qcp4EqvkbWFaXQD5JQZUPNhDEhBLBJz8WSa/dbfcwV0LkYWFNeTgPhKyXTdPjcS1BpwsSU0yTVvArSV5e6pJj/6NQXNSaT+jZaq5mcwoUDcu2Q1MS4V0V6aDpphFFbkr18Ow1E6LeqSzjYFejwe1YPFVtdlki0OJqUUXZrb19N4IhAGoPiuUaN+TJ/foVSOG8Ce9KtKuO5jH+AC2HiX0lCl21+eAiUK5AL00iKMuthLSLAuU4CgJdMKYRGBArkUCZrZWj/oUkv6Snx7xeQNA4W4KJI0zWPhgoplL9dR+fCdwzthy8b+ON/MKYEVwkFDnTmKSjVJdoqOaN1ncp3Vcdpr1tvpmDagpaAYtCSU7skN3Xq9mnCW2Th2aj17x7033ZDA8TZcUWVLU6yC36T0LXrnvOkMQFFXvImqrBAUl/qMJzDhBVXJ7qdcv5WsZYPKUn0qrTVn2y6qaL0UUlhhiX3xDNrRAlzU/Pltxdi+rT6ZJ/VVd7K9Eu+rT/YWe+3q2+RCCmWWHQImWLs8r8UZcl4l8PZYlvZPCam4Xa6bpPQTXFIgbq1tGVPk3VA7gXRFOnElixuT/VhRK06MzYafFmxSqY6tveb00Xh66VBt6BLKCawo+h0XJuorygECaUYXFll3qMSfCRWjQxvH+9WmNR/PYhuuFt9lTwFPAU+BK6SAByyukHD+MU8BTwFPge1CAQm6v0J9fUAJATqC+Wfc3Lv2u/lvvdnVZHAwWFp20eyES6ZSV72pJ64MIbtp0WORYO6fyjEpABO4zN0SDDvCDjSHcc3Ed35DuM1lzCHCEL5bIrAf4IFZQ1CvuVniWSwM+A0rDcosx5gw4TiftBNAw9pIOVhZGJByRN9pI9YcFjycPLixOqREDAlzSWWCe7PoMLDiDNf6/MDh3DOtbj4BWCweh1mCmIWIPc/fTRfV+q52a+56x0+7uW96qQJxP+LajxvNEE7igom+MXYPaCwfFWjx5/p+xdcItKAO+m/0NIsSyrV+G31N9a7sDuxs/d7V0xUPxRU/uIVc3shzTRBL47vW6WaBBKiSFQaVdm8wLW3wGbm4qfSzwZhkKPWxsWRNPvhrEukIswj7G+1+W8DGRiwXON3eYEqWGCe0+KYEWKwL/GhL6tiXVQJxLK4ndy2soV9Q+nql1ymh0Qso/AQa2GqvzQnWPdq0xL3hYg//Pv3+k8rnBaJXvHK21oPsA1hDaA9OZTmxoji+vWolXpWQdCIbZI0BLmWGbqAU7zdkX8feTX/If5TyKraFvNykwUScBG19V2D7gvcl70oD67cWwdSb87jes/OJzLXCmmg4I8HvjIS1c5Ln7haykws4bSs+znyW5rujSnxooLggvXbabnXSZ2an3bJA01zuo/q//dGn+i9Z2HFdxc/ZcoP4wjvEeHM+5czIme0dSsTxeqNeLnKupmUzSCW4rwi0qA8tLSIJ8wUcFIN+FPQ7ebMx1Vb8Cr2e0mQjcP01wRktif2xnuV9Q6qHsZuvxMXX6vuiLDC6U3taC63V8XTl2MR+xbnA9dToCnr5oLcmF1SJ3m9drdKhW079uVdLljyc1bjHmeycphDDbEGxFkYyA6oOPqJcY3FlMDu773SvMdWJWqcbDeGTtyjbp2du7t6+87bexqGHksnFZ6KJzpoMOjI2CIWuq1aHVhf0/+xVFNOCNH8qiJJMQM7v676dUV/4SPgSPAU8BTwFPAW2NAXKgpst3VHfOU8BTwFPAU+By6eABNx36ylcET2iRLDpOTf+yre5qdcfcN2joeserrlkl1SnZI1Qu/lvBVZgov6QEu6JYLoAOBCQWYBs7hH/AvAAwTyCdz6xyOATa4UHlcwVFL9j6cD7ysAEWCvqwQ0RjA9AAn9bXASEdZjB45IIgf9HlLCGMKF6WYvfGE805ABahkGHlbgADXiOa0GJPENXDkpoOfNJwkqDchDUUIcpA9j3MthiDKMJQU2wMwz0qgRgg3WCtcHib9AGA2lglI3pbEqVLnZTb+y6sZdUhhYvZwKDA9CgXf3gqH2MHWN432hMR926sg9ABoALJcm0hqmP0GuU+JvfEIQZwMLfdm/oQsDSlbXAP+UpMKSAZKRFpv/Wq5XwcLWSPBEnkXx7a88JZE0QDq2tijjUPMyKephEzEmFBc5SaYRrnRZzEs7ulxuou6XFeoc0nu+sVqLbBGhg4cU6Pqdw5xrTnj79zKgNd+gTgdbmdrLu/k7p35Ta+n/qO25L/OUpcJYCuIITQNeTlcSiAL5DvTR7XGtjRetqVW+kriYSqaXfhWko2jZ2Fbn847tgXZrjG4IvEgnmY/nUb2q9IcAtv7O2E6UDuaRrJEk0k8ThHgGpr1Dn94l294hWb4mC+HXSWX+FNqvb5cLu7l4//bI8z/YING0q5s6sqLqnVo2bs1ONeHW9Gwtc9Dz6dTZ7Rq6LGBfOqiiCvIExVnq90vtk3RBUGhOuNjHjKmMTAi6EHwi8iCu1gcAKne/A+/RiWqmHaycn4rWT463VExOZ/o7TTsK5FatVrOg+pIRbTc7PWEac1AbPWXeh2ui9qTnb+trKWF9HvzNHWb3TqgrqPStrCs5/AidkCQWgEgyDcnN+xi1gObbEWcpSRhjnD9cmOn8/Ob/+eHOm/dHmjo1HZ29ebs3uP91PamkS11LN52JHfaKXHXj1iZft2L+6OLO3tfiSB1efnNq9kU/O91yloeM3COZA7Rq26bnTV5YXOxXE+9tEh52vf/v3W3y662yEfXM8BTwFPAU8Ba43CngLi+ttRHx7PAU8BTwFri8KvFLNQQgBg3ariyfX3eTr5lz9JQquPS/v1jOyfR+XYHDSAAGE/AjxYZwOKgECvFUJQT8MF8J93EKZ4N6YKPNrawJ8yoHR4nfq5j5CfP62OBVYV3ChOfZqJZg0QArqp17axDPmDsqEelZH+ZNyEPLTLoutQHnm1ohPXCuhwoy7KKwXzCqC8gEaLE6FxaYoW1RYfzdrnnLfYj/wnbJ4N9NH+m2upeyTdlo/EAzBkCJcbbmx+6uutk9t7J9yT/84zC7jBg1herEEgRmGNozpoxR0NS4fg+JqUHnb1lH0eoNUQta+TC3q8lvRGmRFr9vPQgkAJRxSylH7lDuMwPXktyaUC6hUAbqbQ/c1ulcM8uW+G7RkmaGMyZq0x0/o2Zbc4lhg5qtC3JJ1xLnqOwtIYPGhvO9Xpl9Seq/SP1T6ZaXTm6wsaP/vKP3zUoH/Qc++R/kuyT3IVem4r+R6oIDk5sWG1kBXi2ZFLl5OKQQDbtb6kkFGeivKUX0o8yVJQmWgJMFkX4Hs28DRQv5iReOezovgaf3JvLqeLJKuFm0DuXaSsZZrCKhoCriYELCzUK9V2rLYSja6/SnJrWtp5hr9NJ+TXUqtUo2h+UBxLNYBgFY2usFEo/rsxFj1Ke1nHcW52NBa7fu4M1drCC9ej2IwIIVHMYazFWDx25VuUvpqLBkAKAROuKQmiwq5g0JoL0H9GsoaOrZhfTS8AC367aRx+sjU/kEvfnpsun1Cc2cyqgxORvEwcDV7t51j9d4K17I0inqtyrF+u7JH3/tFNlQGGbowlfXChurpq35Z9gS4Wx3eHiXOiZyPOSuevbCoAKwQhLKhz4P6s11p9KtTu9ZWknr6eGetFsrSoiaQLe61qrKcSI/IBRUxWW6q1AdH9e5cbM4WB265v/8XvVa2cPgzjdvWTsi31SB2qeBM7QkCL2RlMrQ0Oesi6s2iyTfo2V8ULVveNdTF55zP4SngKeApsN0p4AGL7T4DfP89BTwFPAXOQwFp4mPiTiDrO5WwYKi7qTcphOSdCs8535U7oknXP37MJbMrLm4gpIB5QuBOIOz/qIRwHw20tykBVCCY53ezFCi7DCqDCcZwld0g0UpzuQSYgZYxQniAAwT7WFEQPBsQ45ZRW3CVgmXB14zulS0ryr02MMFcpcDY0XaLtcB3tOhoP1YLtNW0r/kbcIQyjCsrB9ze7DLJgIfyfWsLDCp9hH4APgAuxOQwV0r02eJwWJvNPVXTJZU1F4jMu77zZnfy9/qu9feAEoyfATaUCc1ixlauoT5WJoL/7ilwo1EAYZ6Eerk0kiu9frZTMYH3dnvZuCwqBFoMtC8EHfngX5YT/kR+4uN+milwadHWas2lCS2vLLLOkO9vCV2dAl8IwCBMt4wwnr9HXSvSlC0nhvsm/R3tOb+iz3uU2Evu0P2PA2aUg/PqHvsf7kp+Tok97BuUfkb3P3Kdubq6VvT19ZYooLnf1lJY1xvuiSzPaiPgrkiSMJNz/JbczYBQzErQLmmpXELpXKA7LeXry9piRWuJ9/HwHUdMhy3keu4sldSn580Z+trpDoKZybq2lUje5YJmP8BVm4TPQTgpGs0LwEBxQJG4g0quU5RAiiCJ4pcF0jwXOHG8koTQb0LfBa4GR+QeCvBnwHr3oMW1X6YjsIKzJ2coLIIBKu5V0oSQDY1wvChRaKR8QPwIszBoZWnv8aETwiiUu6cAy+HhBWiRdmO3cmyyf/LJHT8/uXvtmwVEJLKekDVGIWvV4hEBCacFGPTbq/X9q8fHd20sNgcCOiqt5Ua9u6H4EZpIXCq/Sf1fLHtoYdEWeMHZ2M6jnAPPZpJ3JoEQAyewZKk61itq471jM7h/muzcp/ruP/743KmkNuiNzbQX4jDb6GzUZrMsqk/vXs317H61ryZ8ZnrnbVlPgMnhmZsHi4c+WX1tr1V3G8sVp8DgAiuGZ8+zdaqNVcWwuDvvZa/RfWLcoejjL08BTwFPAU8BT4HzUsADFn5yeAp4CngKeAo8jwISaMPofKMSsQ9gss4Ewd7zPS9xtd1N1z+97hIJx+uzHRcNFccQVGBF8Skl3DER6wGtrn81en4zOGGCOBO8m3WBBXGGySoDG2aBYSCGASTkgSlC2E8ZBCE0YATA4StHbTP/vdbXMnhh9RiIwHOAL9RFwvKCOgBSsFigbjpt1hgWaNuCZptmG3WRtxzfweqCoeQ56xd56ANWEHw36w7AC8ql/dRvwbfL9ATIgJGWD4Jkw1X2jrm7fvU299mvW3e9o2ZhQh78I9MPaPSNGuPPCLSgTn95CtzIFCjkG75XFIMl/G5L0zmU8G8saUd39LMslruVgQSqk4pZ0ZTGeK48ioUbtZEsSojIJtOPw3BZwtgjEsRqvRSsfdahAYVXhTZ//OHP297gbt8/6+QaZuhSTm5iCgUVL/vXMB/n7LX/jxLuSNiznue+amSN8df6DeEQgAXXTyixLwK0+stTAAowp2RNURyXhVFNzp8kTnUNebjREsln5UhtIJFsU76jakNAQ3lkyaR77jiWGfr7qF5Ih4dg4PXpRu1LOsqT47VQhAKtGFP8iinFz5Fm+kC+54r9og+u52q9tNA5Ik+Vh3duUwSfjKXd3styia1dK0niY3JHV+2nwXitKlsXuflRPjsHnE/Z4kvar+1YuICJc3WbvZXxAKiQAkzwdqHaDwgpwA3mGfeWcUVWFXW5Rhofghe6NmRNcFTxK5r6Veev4LDuWay0s3XkWXDTkc/tumPp8PTTlXo6ddPdxx6RG6anZeEwFyfZJ+X6qXPssfn/TtYVO9srjXHFwNDcEhiQPW+7P1ummqP3WGAKMCjgmMtRAw9S1ZELnIjk/qkr0GJqZu/KLt3bRewVTrYz+1Ze3l2v7pe7qqbcQU1121XADc6jJ2Xx0YzCDEvjThS5alY4WYYU4fiOtDa1J711uqM53Ejcs49Uo7yIFBpD71lcRCkCuWLjfI/QGs6ivyxa/xfoJEsLH1dpOy4232dPAU8BT4FLoIAHLC6BSD6Lp4CngKfANqQAQV0JJI1g/nGlvW73P75J7p+kMVgNXPOuzBVZ6pI9sSIJ/qV+h3vCZ/PTo+9/rE8LnF0W2p8Vyul3AyvKVgfmTgmSl7WzLNi2DQWACvdgoIjNQF1mCUEZuG+C2Tf3UZtdMm3m9kwggCslGD1ACoT8gDWAFCTemdRppvXEmoA+1A0wAENbdt10vr7Qh+eY5486RXuxFEE4CagASISVBd8BJNBGw6Jjc19o65n2hbHak7Vd4/Yx99JfiNzD7ySvuZyiP/hHhjaAH4zxb4zq9h+eAtc1BS7gMqloNirdTi89pZVRjYKwoagun5SrlW57Pd0j9yrzWgAzckwhOUkRScXZSTCY4qqlX+D2Ke+5sJBctkg60m6WD5djimmxJhDkRQUszhOsF5oP9yIBFJG0qxMFAEcUFa63+/IoI33sIAurFQXciIYOy9lTaBfrnb8/oMS+g1XZk0oALZsvgIkfV/oqJSy40G79FtHzF7zm9nU95a9m4wx8X9U6+IKElm2JzDek8b8i3fBmNij2ZEF2lzIp1naxpnWkd1+h92SxqDy8+5Z0z4B53mP5VrSuON+A7JwdC9odlOJdZTDI9mjvCLVeN3BPJzd01Wa9Amja6/Sko67IXwKFItFRgmC3UaTFugTCE91ef7I/qEzKUgU6KhCzOzgY5A3tV7iAS/1avZrL4Tl1sT+zb/KZSvKOXcMDuH+S66dEcSMEHmhL1s04qcrKonosjJK6QIw1WVrwHPszCSvjoQunTVdTAMA3d1ZrTygV64tj5LlPVhZ3KAB2LQjzw1qPUb+TVJRvRlYV5ypjVOTQelBBJIZgF2dGc1MKUMI1POdqog4Ut4Lz7EFZdRxR3IpY5e7prMkOsZrK8VN28/iOjQnlay4emlmX2yq5LQvXehuVTyjgd3difv2uWpzP63f5vXJRlLgva0wVrT13ZX15fzrca8luKHWzayfD3ctHKmIV5BpLG8Wwev4VQ+vtQ0ofVzo2cg/lQYtrNsV9xZ4CngKeAtcvBTxgcf2OjW+Zp4CngKfANaGANO9hstDaxaUQmlCvcPWFwO382j3izHIXjYcuFD8UTa8JrHhMv+OKCYDiT5RwP/LVSpjLw+CVNYMNFDAAowxe8N3uw7hYkG1oYL/x3YT1/I7QDkABBs6CX5tlhmkhA1igFWdllNtUtu7gPi4bEOqjJYrrJYT6MHyAC5RhfQEY4Z4xg3w3YKDcXvJvdgF1rr5wj+ehGbT8pBJCRvpH+3lXAwQRe2KHkvk4Lgf3tkDcfY2JfAWMHXbjr9jndrxz0S3+Mb8B8PAcoNIzSljAvF5j/buyskA721+eAjcqBYaCfAkFs/4gW88G+YletweOzwAAIABJREFUVlQqcsyi/6paWTvlV16ubvIIAWIlidYU76IrIANhrFQ/wzUpgHbjJGxLO7onICMQUDD0w/9iCgnP50pG1QSTzVrU7qYNta0hz1Wh2lmrqZGBK9JUbqzWW70iiaNcv+sKu2oiIKRZZX1C3wE3WePPAyxGbrMe0m/vUmKP5sJFFN/R+vXXNqcA4IIANbNUJIj2aQnVxzT/pgdFwHsD12nSGNd7tJAVkoSxuoebyGNYKGkBAqbzzsLKctsJHrXXBDjIkgEXuvXVmYnG9Hq711LsikzWW50wkpZHEYa1quDHLJvO0nxcj9RE21Qk3Z3KJGN1I11vNtKToi3gTyrRsaS+hQJ5+9jb13h5cs6aV8Ka4j6Nz1cQo6LanNRRK1E4kt7QFRTy+KhSSfXWGVdg6aZusCY4m3K+O+NS9cy58VxB6ZflIuop/Xa/AIQH9BlLHWhKT37FKL/KG7qiusglMwZFllMmzqYWf80mkMVaoy036Z1XyA1VKBAkUmwKAQ061BfBPC6nAEYEkKQCKhqKmZHqd7laLQK5r/oH1UbaHZ/bOAo6p4vzKF80s9W5erEaDdznFMPiI62loFWfSv9tcbjYnQviGW4dI8BCj0ADzqK4KeXMHQi08JYWFxte/7ungKeAp8A2pIAHLLbhoPsuewp4CngKXIQCP6nf0eQnfgIMyaLb8XX7XDTWFxMWu/bjx9zEaz8vbo3fYcZgtLA2QCCGVQYa/2Z6XrZkMMbJBPTmOsneRWWLi3Ig6s3AB83nHgwZ4AJxGrC0QNMTwZ2Vi6AFhsj+NldRBiJw32Jq0LZFpYNKgCBHlbBsMLdN1Gnt43fTdgZQoO8widQPY1uOYYG2qQEaZbDF+mAgjgEmmNkDWpRdQVHH3UowebTXLD8QDpmrK+qkHWcY5CiRWtvOgZv58kiABW2gb+SFXowbfeA7Y/39NMZfngI3MAXyei3pry31VgQ4hBL6jwVJMBUncavT7R+RT/nT/V7W6EtlOU31Lx3MK1umZ9YkFFyR2vjRWi15IgnDVbnB6QsgyMfHqrY2v9RkCTs9xd5NwvE8d1PSth6T66pp7bX5WislNsDkuKvNCb84Le1tgp2uK+AxewqAJheaqoCQa9LEDs4FsoxcQ+EWqnx9k/L/e/227QTMX+oBvRHL3wRaVLUu+hJCYpHHewaAgvcLa6LmcrlNU9BdCdaP6HWT6vPkKN+2DObeqCeuVkkqivvRWNvoN2XtdZvi5TQVp6KZ5oNKp1s0BTRWBDT2pfMhK1UBkbniE6dpLOuVeiSwtBbkTe1DRwoXrrUHg/F+P2tg6dLrD7QB1OzMdCNOrRumzedwB8W5inMXsYJOydXT++Ja48H6xOwwuHYgf0hJreEGPXlGTaqZjl2pLC/OxGALAqzeUKThnMXZE+UeAnUDXHAuLV+ML6AyoIS5I53QauMcznmPc/ilXJz1WKuUYQoznJOpH0tpzuZPCBxJ025lh0CJjcn59Sfl+olz62sFujSJrdE63XCVWnq4301qyjOb9aPXC6yRNUmxGET5E5WGZu+ZMzhnbMqmTyuar0dlcFJUm0V34f7BXllaPJr33ZEjfx/fl6XPeZ3SNuJ/EEftZ5T+q9JHRH9Az+e9j+Qy6lL67vN4CngKeAp4CmxBCnjAYgsOqu+Sp4CngKfAlVJAGvf79SwCCpich5Ve5aal5DV+76wLK8tusFZ38fSiwAuYsb8bMRcIv983YmBepc/NrpGM2TbwwuI2wMHwHjKGygCNze+mMqfDswjqJCgZCt2xiniZEgyXBfxEyxiGDZN4vvNJGTBz5lrKQAxIRb1ow1HeghLAA22A8TQLB9oOI8VvCP5pA0wa3+kvgABMKJ/URz0WA4M67NosBLV2mLUJlhwwp8QOoW/0k0DiuHGC2TSAgn7RPqMZY0Z9lEPbZqQ5/qyb/ZopN/2Hz7jTHyH47puVYJrpE1Ycdym1GHNZWSD09JenwHVLgXIw6XM0kuDb8lcjFyxhsS4N5rzXy05Js/nvtfRPFVlwl6wv4l4/n5BQcLkSxwfHFOVC+IU8tUhLXPErut301CCKlnWrJXcu2ZcasJBG+9CKTFYdFcWpiGU9MS2h0IFUbmAItaFA4JGAixn9vatWGci8Inqql7u2/pYjjkKYTNSSDQbrnr2AvY1EUO7zAS1o1n6r0m+O6Pcj+iQGho9jc93O+qveMOYO72PehwIimFMFbg8B0ht46leGOQEUe/R9Vb/rfVcwB3nvIVjl/bit3EExQoox4wQouk43XdMes4TBhdamthGJcHNXl//MBkEpBEgqoHKwLhPVrtZ2RWu4kMcnuX2KXKMmzfwwqlcq4bTAjknl78nKIpXBFWPSxS2UPp+3ti+yL171CXQjV1gWjI+CbAMMs6/eLgDihwRKvLk2Pi3Pm8kwEauiKAheXXsojCu3CpSS9dEZt09aG2ZNO1wTSljJYkXLd86OjCXrbI8S5z0USQ4q3anEWRLlG/Kale/FSMv5lHcB53bKXVAyN6DUy72XKmEFHSoWhjv19Ozu9VPNO2VJEU3uWpOlReTkFsoJoJAFSe9Id6O6L+1I96UYtmM5SqOn6xPdT0dxRh85L/Pu4KzLmZd7k6jLVMeKd1XqxVqWBofu+dr0E91W8Esnn4y+V7+jXLT5+r5Rm9lHDGS5WsoCF6Op/91TwFPAU8BT4BpTwAMW13gAfPWeAp4CngLXGQW+Re1BEI7P29YwJkLt5l3yTCIhdzDl6gfEydwiJcAIl0IwKAjREWbAYJ1La6wcv8I0p8zdk7ltMmsMSGGMyuZPAzt41kzeEejD3MFQmiYcwngYPbPKMKsGAwRgikwzjHcgDB4CGrRHaR/gA7/TJ3OVRPkGDtBnBH/GTBqAwu9ohxkAwSfMXDnYt/1W9vFg7aLvABW0HwbXaIRmH1p50AgtVgAlLpjFoSn9qA4LCE6boc+Gi+JZV1tI3a5v2+lWP3any/vkxwKG8imHMUbQxJgTiNdfngI3LAVGro/yY6fWN3CbJGuKzlilshKHyU7JCtvtXjqjRTXZaFTlEip4VsLCSIunIQBgQ1rMB3XvtASHa5Iypu+496arZXWQEFxXQsm6do55aWjfLWHwuAL0BqtrnaUgCmcVMnyP2reidt4kAeg0AbiVf0PNx6qC+D0Ivyw4b/cCAsyBhJ5/Nlrz7DXscW9T+oMbdtB9w19UCpSsLHiv8b7gQosaEHxW6B7vId4ZK5qnvDvJxyfCUFN0uFpr50Xt+5UWhlUTz8pKqiv3T2vSMD8mv26HiyBora8XuwpBjfqeyrVTKPduWsLhIJE7KAAOxbNIO2kWxnGQ16vRsqypUgEVnbFatS/l/Vz7WE37EfTflpYrVzomL9JzdtbkjHu/0puxqogVWFsAhXx/ma8uLYkoudMF+Vql2ftYXCneLLdKs4Pe0LC2K4sFzoXMEYthgWIN5zTcjgJWcHF25jzGfo4yEGPOns7FWfNSLtqLwgtuXDnbUg9nZBrC+ZA+nD17KmaF67eqsg6J5RQqTxX0O9P3CbmkGtbVXq2jxIK1L+fWP5ELqJqAioHcRVEu51r6ZC4IATUBLQBEcDOYyTlVL6oUByfni/D17+u1//Qn6/+ysxb83vMht2F1X6n0F0qcTSmTvecsaIHli7eyuJQp4PN4CngKeApsPQp4wGLrjanvkaeAp4CnwBVRQJr2aPFjqWAgw4KrKnbFjrfvdJX5rguTuhQsHxFzZtYE+0YVwajAsJhGmQnbYThMY2roE16XuXriu1lekAdGxeIwlLWrEH6U31WUA7MnzWn36tF3nkdoZ1YGZasF2sYzBgTwCTNIXSZwIfAfQAWMKYFrMcs3KxGzzrC+mNspyoShpG0wmwh0YOTM9RJt4lnrF3kNEKHv5asM6hjwwnO0h/ZSN+PC3zC/9JULJhRaUDf5+RsaAKrQx1xjNnDjrznupt6yxy1/AGsNBJW4m1pQsrGZZ+xlZYHLAH95CtywFBi5Q8pkvZDfe9eeol5Jsr48cQuMWJKrqHpQjXfIkiGXy5Y1aTGjAp0mSbQhf/NL441qKpdLvXc8sN/2qqtBh6rq3NHpBzW5o6pKWBlKwDUv/+I3aXUuyfUOwTTmev3sZoXbWGzUK7KwyDY22u5zg8wtKXj4QMnccrC3phKgZheIvYEA698o/fSoc7+v/FXl93FsrsZo3wB1jEALWsq7h3c0Lma4mCMmpDRFAN5p5XfrlrauwIrrPFdB7BtF+6hEQbjc6vafTjOBO0FwUkGIM7l3qgrgqQQuVFBt1+xluYwwAoWqkZhbCznNo7g7yOb1Zyrg43OTzWpfOvxdgZnrOjHxfr/Qmr4BZtWN1UQJyJnnnGkR2L9e4/jNAExClnABVSiYdlnpRJYWQVMeoZ6YmGsv42ap2ujPrByfIGhDU/9pHF1PO/tJgQSfVzwHxUwaxoUBsChfnNvsHmA07qDsjH0+Appg3+K5ASSg4MI5ERARAKMcf+055chyohBA8X4lFFg4FxIMm/xcKAOhnLOktn+0Uk/vuunuY8dn9srzU1hwBuWMbP3gk4v2A3R8XunL1O992jHqCsg9e9db049+4a/jn26fDn9A8TmGMT9G10F9Lij9OyXOqFgA4h7LAJvntNn/4SngKeAp4CmwvSjgAYvtNd6+t54CngKeAheiwBv1I4wHWv3DQJtu93t3yv1T7vJuKg7jiGu8HKEFWlRm1o6A3AT2MEvGyCFAL1tOcN9YFAMh+LQ8FufBLA4sL7+bv1zT+oQZQ3gPs0Y7YSzNjy6f5vbJgohSN88AJmD1QF24Q0LQAkOGZhsm+QQZRyJxTAktNwMGeJbL3EEZUDEUEI7KNuE/IAW/U48BI1hG0N4zIMIZoY9ZjFCuATcW74J7MK/GFFp+2r3ZKoV6DEzhdywvaBP3ATCedo07G273t68KsIAegCq0wxJ+hD+jxNh7wOLMOPvrBqcAQld1of/+Tx3JFk+3OvIBz9oYEzixjBsWmV8EAgqcpIa9sVrSrVcn2AsyWVZcTbCCdS2/IkHT5cEu7Vq75T5coSwUlzfPK/00PyBwJVNMi2Hw3TzPZlrtoNGPw5YrerVGo3LzbFyPiyJsS7AJEMF+yP7M2j+nljvxKiR0/eCm4X257n2aOBc3+LD75r8ACgjkKz9dVhpgTgHu824sKyAgsDTLHvJvabDiAqQd9l0WFMT8WJto1uJ2t7+e5K6heBV9BdlWgGJ3kywrEsmHlTeQl39dClyuoBaFqyaZApyvy55CN10iAGNM6/m0vmvn6q9Ukjr0x+WdnROe0xTvEuoFTPpzPDoCK5CPIPj/LqV75KrLVRrjAivGBE6E5bPbmRIUgDovwl6UZMW+206dqE928u567diRz+3aKLLwMblbqtcnu89sLI0dP/3s5JjcLt0u4CIXcMG+zTmPhMIQIAVnP+bUmTP4me/nktdgycDZjXzmaoq8nEux1GDevHXURXMbaGDEb+g+70QCXz+o9DdKnFGH7qxkTbGhU+lnNUl7UZQvj820qvtf+ezhnbcuNmWNwXmfMy1nScrAcgTrDS475/MuQskGK74lka932+sGlR3785NP/m38Z0ceiV7d3QimBMxzkYd4ca9Rgh5/qIRVCed17xpqRFj/4SngKeApsF0p4AGL7Tryvt+eAp4CngIlCkjD/s368z4li/PQcbV9dQm7Z8W9SEDWX1Eci1PyTgtjNGRqdCEYN5N2wAqL/QDDZACECTjMVRFMjr17nqOlNirTBPrWujLQgUAdJsisGmCwLG4DAkcEKAaAUA7t+ZASbk8AHXD7xD0AFzTYYN5MS4zfFkblAVaQz8zyqQNgBjCCTwNp6DOMGcAA/bIA3sf13VxlWBkweUYT+maWF2WXVUYX+kJe+9tACuoox62gHHNFBWhjjC0CS9pKe253UeUhN/XAF1ysrIMN6EP/0Mgz/8OUf5/mwBOysvgwhfrLU2ArUGDk2in77Y8+lc1OSdaPQxYpQktSVCx2JV8UDCs3N/nuufH8AlYJXypSDC3BhE5UekWqIOCVpFGPlqRlLQcxoYJu5xMuywMF5FWEXgXwlW/weuwkzCz2K0J3RX0hKGtdgq+BQI3jEnICtLJ3WDDu87WbODa/pvTeUQYADFzFnfpSddSXe0NSwISFQ/Bv1APexyY4Z64NBA5uKxdQ5xnJ4TuaGAb1WiIA0R0SCHGLRNsSYTuFxgnHda8qk4qlahzWWt2Cc4Fc04VBTc6hXBEsK7bOM9VKZb3SSNpxGLQrstVoNioWQ8HT+OovIeY958ZE8SkW42p9R1KryxtqLtBC0JNcKpFYDUktJUi1W3jV4ZnmTGsPaNTE/PrtzdnWpzqr9Ycnd68+GMX5a7RXt7trtWef+sT+U+uLY3f3NmozeXYW/1gY7cGAAebuk3mFMs25Ls6vWCQAdhAbgvMo8wrLClOWYd3yO2dSzo8GWLxH339Z6Wb1paH3xyvVr25cHRwmLo2Cay+NzbQfygfh0Zm9pyd333lyvFLvV5WXcyagCtYYgAtmmfFb+k5sDDoDT0BcOfKRn7yfqNSK5o5bsn31yaI9uy//0ON/Fb995WhYU33GT9BHzsk/pPSflHBVCB08kA5l/OUp4CngKbBNKeABi2068L7bngKeAp4Cmyjw9fobhgf/twiuFtzYnfkwdkU8s+HiqcRFU7wzYC5giAAuEPbD1MEIISCHSTJrABhsAysAAwjQDVOFRQMMmLmGokxzibT5WROMGIhxQHkxN6c+s0ZAM8uEKFYnXbNnAGLQ1DLXFTBZMG8I7T+rBFOF0J/ysLBACAMogusk6gdYgOkzt1UIBWk/pu88wycCQvrPdxgtGDYYNRKabmiQ0Z6hJuaoXAQRXNb3srUJ42AAiQmNqN8078qalrSBeniesqAr/YHRg1a0dber7D/ixu8/6k5/CNrRHvLz3EEl3B4Qk4Q54AGL0cD4j61DgXe/8cBQoGj+5hVQ273r1TdfM+1NabPbXjfcDwSaJHIOvjMvkkyAhPaSYiyMohkt0ijr52hob0gbdbrXTaWRHeEqZqo/yJsK4ntoYtyt1itxoYgc7AXDPZh+ng+AGVlZ/O/KZ4AF+8A/0DMInYbCIa+1vXXm/qX2RMDDubKeBS1GFhhlhYKhEN0sM87z/KVWf6Png05Deii+TJKfsZZ4UuFpArmeG+RJWBvIvVuCTr1uVpJ8ViCGSyrhQCsu0o11xalBsCs3b/GpNFPg7jxEoeDsu/4aAKo3+phcdvtH1hWcoRhLzoPD86b239vzQV+6H6GrNXuuMdVxrdMNlw1CNzbddrXx3jPjcxtdART3af/eKyiDc+KU/n5Avx/RPSn+uDuIdhHPtu7d/8rDbvHg7Mbxx3cm3fWqgtvLyu7MGZPzMGdkgAXW2oXAZ86DnN2YJ5xX7UzJmY8z/KeUFpQ4I2MtwpmSPuHylD7eLouQU+pPKOuPp3YsLH1KYEojqmTV6T2rA83U2agyeHR8R2tSYAbKTFhpAKbcrcQZkrM0AAOgCZa9nJ1pC79zH7etzF/qOqZvXyZLi/HmbL4+d6tbqjSKX/zYb1Zem/aCV+n38vV2/QFQhKvWL2z6zf/pKeAp4CngKbDNKOABi2024L67ngKeAp4CmykgzfpX6h4MGiAEjBNMxpgbe0Xo4oZcKddmFMPilFTLLEYCLpQAK4xB4hNmqwwYwLxwDwH4s0oLSn+ihAsiBPIwMeaj1lTMTJPKgA4DIiwINfUgXOP5P1V6UIl6yq6ozG0UzJUJ7mHU8HcB0AKAAVOF1hnCPQALyocx5J5ZXSDYp4/0id9JMGAwhoABmKybdYe5jrIg4AgviIXxlBLMIv0z834sO9BKK/cRQQV/Y1pvAgqLvWG0KVtiKNtzXErxt4FGfKcsGEjcXtH+0xq7O92u935OgAVxP8w1FXVgpcInY3+auSAri09TiL88BbYaBa4Xod8oTgBrWtYRQVvWEqck4byl0+3vlNuqUP7t01A4hgRlAjLycQUDb8vaImz3B0l/kE0J+pxM5SZKz8iNSPDxYqxwCsZdqCzWvgncLgTIPK18/4fSj47G+Mf1+f7hXqELX/0etNhqs/+F9acESFwzoO+F9eCFP32BNYHLJnMPmcvt3E4ZbglYDFOBo1Wt4eXBoHhCoIRWt5tSvOaurCrWG5V44OQCbrxZeSbt5QrUnS+zHyi6cVeABmeZoTuoUXrhHfAlXIwC7J+c51A++UdKP8bfRZG5pBG68bk1ARYyiJG52/jcuku7idt954n18dnWZyX0f1zAxAOjCswqIpFVwlfrHudgQIQx/b1zYm6j19uoHlVg6z0KYl302xWL6cD580Elxh5wgbMr9zjPnevCMg6LubI7UfoAkEEqX5xnOed+TmkfwPjU7rXfkruq8fEdGzsnd62/VBYVUVJPpwVkQAPOryeVjzMoZ37OvB8bfTIvSbwvzHIDF1UAGrSV9gBkcEYmDgfunjh3r+gNNRify4/3W0FaHXeZVKI2Axa0mTMx51RAmecE4N7UJ/+np4CngKeAp8AWp8C53HFs8S777nkKeAp4CngKbKLA146YEIt9AGNxTNYVp1w8J9Biuu/CJmABwn0YMZiZcswJc1nEO8XeKzAaWDLAdPAM2rtYOnCZEN7y2t8We4J2cBmjbi6mqIfyELC/RWlh9LfVC5N0Bmw5A2IYgILvbfMJTNuxrqAsrElgqHgeZo5nhm4uSuWa+ymYMJhDNMvMR/xZW/5Re9EqQ5ONNsIsQi+YOLNaoU6eNzdXJvgxC4myCw6+G2AzKv4smGF0JA/tph0GNBngwae5qFoY/j7/DfQPqxIYTEAktADpC8mCiTMX/OUp4ClwdSggi4pgVWl5GGBXa1mWEvIUE8pVVS6hZaBwG3m20UkbcnTfEEIRDbK8phx5rDzaIGrKMydLi30SirJfmGu8zXvTc3ozilfxH0o3AVG/cbSXXJ2e+1o8BbYQBUZrirNDS6DDqSiKPi9ri0fGGpXjzUb18Ymx2t9OjNcfm54Z+8L8TOPR6anaM5Vq8rEkDj6mEAhPRHFwUM8phcsCMDtKCKtZz9fCXd0WGpnL6gp7KOe2r1L6QaU6EHBS7Q8tKWZvPu7qk4os0qpgVZHL+mBVn6uVRv+ArBA4+yGw33wJvApeMehH75fVwicZ0zDOpxS8ujF3y1Iqa4bxKHlefGnAAFygAkY8fIEecKYEXLmYPOcg81KJs+i8ToyPCDj55My+05/b9ZKTRyd3r23I5dO+2kR3Z5wMZNFXHFSKlQATOGtTB+d4zodYEHPGBUjgLMl51M6S/AaIwbwlLhrPoCjEOZr3G+do1eFur08VS3O3ZF9QW7Bi2Xx9v258uxJAB2dcf3kKeAp4CngKbFMKeAuLbTrwvtueAp4CngJQQBr1AAswO7hrgpmC2Zh01b3PuB1f99UuXZQGYO2o4lnAoOAqqQwEmEWEuXcyl0doR8GBYc79ISU0xH5T6YdH9y1/WahWdiFllhvDJirxrrIYGOYWiXaUf6N9CN3N1zNlkIe6+Q2GChDBtLbMVN3AEdqEEJ88fIe5oy4DAAxMgRGDKaM95gLLgAGLS2GBSAErHhy1E6YODTWznCgzmNQBk1y2urAyyxYWBmgAjNA+LsrjIl/ZQoV7tN9cRe1w0Th1MCbQEwYU8ALtN8aL8mBOn2FOyMoCRtRf1xEFet99tjFn3YSUm1f9j9dRY31TLpUCmYJ/Z1KvJWjvuqJrZHnmgkrVnUwHxbTAiXFZWxTddNCuJtFinMhJhxzhK+5FR/krAjEmJD7DP/6RajVi37kc7XcESR9QIsYP188r4Td8GMvCW1lc6hD6fJ4Cz9ubOSdkAh8+L+hxEUupMAmSah4MNcf7RTCh0DRVF+ZH2r2i3e6lrlaJT9eTuFVJInOt0x+BIJ68V4ECI3dQKI9gTcAYzGrcXH2icDsW2FrXXbUenG5Mn94QuNyd3rMWxbW0qDb6YVKT5UyScX7iDIh7zaFgftRs7e7BDoEW35r24knFssjCOFuX4zApBQmgrgwWxuda1dXj41X9wpmSCyUbznZfOSrrfBTgLIDV78WE+gsUIFBlvdrs/VZjovtkfaqTzC0spQoQflr9lPuyAoUcrCKwwCAYN+0/oIRCC+6ZsDDmPE2d1MfvnGtRAOKsSZ9pM8AE50doiKXz0dGzfGJx3FAJB0XXT9/++sG+k09G/7y1HPzaOTrIiQeehLP8xeIyneNxf8tTwFPAU8BTYCtQwAMWW2EUfR88BTwFPAWunAIP6lEYLYTdMBswHn03ef8Blx5dcxMP1Fz9AMJ5GBWYOa5yQG0DGmBiTMMX7g7NMPIjpEfrDEBE7kuGlgAWnJuyLIaDBcs26wMT1NunMXLGmHHfwAZrj7ldokyYJxgt2kKfLEA35ZsLKz4R1FMO2mL0kbbyCThjFh68K2kf5fIMdDIGylw10Rfy0Qa0lWkfZQCCYNVh5vjUxfNlF08AK1zmB9toQRnQ3lxTGX0RNNJGo9VmmpWFlpRBu6jzje6txcPug8Ff6DtBEWkf5VvQQ/rHXHhQCfcw/rqKFCgBEtRq64m5YECWWRAxxxhj5pIBb4GeN8sgniEPY4vQYAgkCtDIlOc5mve6dzkC7qtIja1flVzs5PL/z5j1FKB3Q7HAj8vv/YLcxtyUF2EqN1CpYoRvJEk4SAdhKijjuAL6TvcC12x1006tEi67Qj7wA1lZKLqvQI9mp5uuKg97k4GX5yWkhKF9gRKAyAZYkPcfK+Eq6qLPb/0R8j30FLg8CgAwAPSV9t1AlhLcqOV5IeUPHUgGLK1iLY6DeiWpLNYqSauXKsyF3L4JrLDziAcrLo/0L0Zu3rO8N4m3xtXkbalYC252vwKNxHkxuTtPG1PdYHxn6xn9NBFXsnlZKtQl7Ecwz9hx9mOAEfq3Bv34VEc2GCqnmXYZ+R2yAAAgAElEQVTjncobKWZEUWvmCrWet3beulib2rMarJ4YV6STfcX6yWYFd1O6AAMAEM7nCsr6y15/roDsKB5x9j57KZC2U0yNfPqm1dfJuqOjevtBmPfCQIZ6wbAe2o8yDJZ2uDflLMx5HfeBH1HCZekbdGJQ8CfZ+mXBw/1u8oFKPf1O3ZfVX14R8EG9nJGhIfHbcJ/1XwXYPCQavUT9B8ygX3PJmSDcC6/9lt7hD/1c7YSA+vlNpxHaQrwNL6sqD6T/7ingKeApsM0o4F8C22zAfXc9BTwFPAU2UeCd+httKKwBiGURuek3fMHNvmPBNV9VdVETgTsWBeYuCc18E7bDmJUtD8iD4B9NLPNBS/6/VkIwZq6UYGosXoMJUM2iwNwgDbl6JX4vgxcW9NPABP6G0aId9AMhrQEvJuxFC4wYDbSN9x7tIE8ZJMFfL+0iYCBAC+0wKwqYLP7mGYTEMKfUb7ErrM3WTphIABLy0E9zoQUwYO9dE0Lr1tn+0T6YPT7td8osBzOnTNpBn2FIaY/9XhY+l8eIOqEvmnh73N2/1naPvheLE5hB3HYR14LfAZn4ZE54wIKRufqXgQ0W4J65iNCAOcQ8RIiAliJjD3DFXOY+6wBhycLoPnOQOY/gZBgvRmAF6wBBhFkmcW9oDeSBi6s/0KMaWW9rcRRInORmJNRcDOOiUknCqkCIlgZ1h+5XwtApDm8xKc1eV4njJB3I8XkRtCQEamuDSLKsqG20+04gR1+ABfvWpV6fV8bfVcJfO9e/Vfr3SkMLruvNyqIEuJ21MmLu6j77JWuGZC4Kh9ZlNrdHeZz+9mDMpc4On++yKWBWEVo7rEPm6VC5IS8KCYcDLdFQMWuGIQvG9fdqGAedwkWhAAuLC1B4y4rLJvuL8QDnKJRDSO+hQNxBVRUfaFy7cK1ZHKuN58sStOvclN2mt+iZ82MwPDMBSnGWQvDPOe/P8jxYXTk2QVnvTDvJgSDKq/1W1a2farblhimPknxCrqEmqmP9Qq6lugIvws5qXXExzopmOJ9d7DKFhc35ngNWCChwcvnUq0/Iy2CS7Wuv1Aq5g6oLNKkN0ljAQrFbgMxJAQtd9Weg9wqKDh8DjBnRg78BGm7We6efDaLxjaWx2qFP7Z3bc9fxx2tj/bvUlzSppY8ocS45KaDmUK9dvfXkUzvGl56ZvnPfy4/ePH/7yb0COLD05RyiOt09O2/N75ranf/E6WfDn9qkPcE7CJdSnHc5c/t9+2Kzwf/uKeAp4CmwBSngAYstOKi+S54CngKeAheigFz+xHL5M9AnDBeMw+uVEHwecbW9627PPz3gkpnIdZ99zI3diUATbS/eF+byabP1A38jaCcvwAcMOv58YcARtuJmCaYD5ge/vFhaYCHAVXaNZN+NbzHLAQMvDByhXGNeaDdMoYETBliUwQ4DK+irARswVQAsgBy0Gzco9BMXSdy3QN/kN7dLZUGgWUlsbjP1AtLQbxhZmC6+mxUF7QYsoE3mxolP8vIsbaGdAB4wiTC/ACnkoQzKw+UAtKRuPnmG58vAhv48q31vfaGsV7ld377hguqUe+Td5oOYINuMB8AU5X2BuaE5ktlcoTB/vTgUOIclha0nA8UQDGD9wlwhcPqdSghDYNoBArGCYV5+VGlJ6VuU0EZkDrxViXn0/yndNyqDgPOsX8YbbUlAD+aRWRo9qjbxW3ldPa+z3uXUizP+5yhl0E+zjtRTTwSu+LvAhU8pdva8BJwbilMRxEm8Q1rZawIpZHwx0BgpIHcUCpiIl3VjudfLqhtRL9Dvq1EcSVM7DBSA+6xA/0KtlmA0lWAVgMIAC7Lj4mOoHXs1r/NYGFkT2NsMYGa/P/tuGIEY7I0AsqwDhIfk4d2wqt9ZI3zn91B/892EwwaUFx7IuJqjvS3qYv8euobiU0AFc1bv8oD78uyWW8ywVGCFna2GZ5+RlcZziHSBgN/bgphfyk6O3EHxjkRBwCxsXaGR6m4EbuVY6HbfkSVxpeBsyz6E1QRnXcaLMyPPcK57crT35AqqPhPF2RsUWPumk0/uqGb92CX1vuuu1RuNqU6mmBgdgQcD5XMKuh1naaTyB9IsiC0A98W6bFaWnBUveAmMUOyNTlWweEWghQJfF7sVYPuhoFKMnz4yWSgA+MbU7tXl5WenD+VZsDh78+lGNggPKT7HYQEqwtUKzgxvEaCxKquRY5212sKRR3bfu3Js8o1yY/V7s/uXu+pDPammB2ZvXjkuA4yVpx/aP3fy6dn3KT7LHULn1p/6+P5f0ecnd99xYloutHA9xVmmiJJi8sCrB49/+njlQ1k6jJdhF2dRrP9QuvgNJc4//vIU8BTwFPAU2GYU8IDFNhtw311PAU+B7U0BCaBNIwsh99croa2NQBPB6Jrb8TWvc0U/dfFExdVvQSiPYN8E6WhtGZhgrqCMoBYrAUERwlDyAQYg/IKZs2DWMHtmmcB3K492mcubsoujzRYW5DcXUNRtlhAIpRDgPjgqn7ItFgbtAUSgDbz3EG5h+WBm84Ao94w6YgGwed76xDMIjBFymZ9e2sr9cpBbA0koA+YKIRv1GOBilhgGVpC/7NbJBBxYqKBZhtAappgyELLBLJvbAe4zNrQTn8sI6XieOq0eusQ92gktGA9AmS9obDtu3w++0h3+KegCw42AkvFmLjAnvl5zBc3rSJ9DMEUAhr9eAAU2CWQpyQAnmyOM5QGlBSXu8Tv3sIDBpzTXQ0r3jn6DmWfMAJo2X7hgMwuhB/XdADMED4AWv6PEPGSe/RclBC1YYDDPEaQ9LwroOerwt14gBeQWij0gk2uodr8/OCWhpoJZZDelaRBkuZvKE9eOQteWcDOMorAiAVoiVzJay0E/UKgLCTrHCNhdrURrcieTBWFwLvcgF2slc4oIKBYl5cP6vqCE5c6LZmVxjvlP8eX9nfluGs5mSQYAAYBrMZSY08zb20adYk8jLg/rg3sAb1y8z5jrANG4J0E4Rp/sPYPlIL9BL4DcZbWPPdXcDJ61zBiV5z88BS6LAgIYhmtb4MMQoBjNPcpgnmcE1tZn2WKU3zYpmV9WlVeceWR9RN3Pq3+bANWckTirfpMS+81+rCsq9cLN3ZK7vS8fnJiYL9phPLRiZF/h7Mh+8UElFAY4Q7GPIIjn3HazhPsqo9ixdnJ8Iu0mThYJxJAY7kDLz0xHAgx2CBAYKGB3HldTgdB5IeuEfnejWgHEuISLdmKtcLH4FcN6CRoud1Ty5eTCpDKgr4sa7TCpDhaOPLo7WjvV3Kd2vknASXPx0MzJXqvaPnD/IbfztlNHBbXNyLLiSVl/VFvLY3P67LVW6i9XTI7Z1RMT72uv1fdWx3pOlhbz/W7lWd1vbyw13qLy7xGgQVdqaS/4jpNPzP1ec6Z9YOqmldkwLDizrooek/O3Zy+rjRefaZ8O3oLp0ejiQfb04flVoFL4yb/6dW9lcQkTw2fxFPAU8BTYShTwgMVWGk3fF08BTwFPgYtTAAH1+EgIDTNgrpnWXLLjJtd8WejiKbmCGl9z0QzC6zfAbCgh2EE4ZPEODGwoC8gQqCPkwoICASiCVhg43jUISV+rBHMFYGFa/2XOzMo0IX5ZoG/up+ihCbmo2zTHYX5gFM3ygXxm/UB9PEN/6YtZWSAEo1yEtrQTYbEJFyiXfAASlEPCUgIm0dw20QcADGubxRagLu7TfuuTgRmmSWnawtYfBBoI2xBiUP5fKsE8Uz91wiDTP/oMnc3aAzDI2gRIgoDP2mHtpg7uMX7QQuN8b+Qmnlh3s++cc0t/zH3KhoaAFbQRWsEM0851gRVDx9z+etEoAF0ZO+br/UqsC4AH/v5WJeYaAhHmEYCUXVhN2IUlxubrY7oB+MYcIsglABfz2i5ARwumybxlXKnH3L49rO+4CUKYy7ww9zrnqMrfuhwKCJS4UPahZZXAh35QBEWaFS7P3dEgGDT7GgEF2e5GYbQhl1ETsrboKpjvWrc3WFcg7qVaLX5KYbsPdXppDrDRavezd7/xwCULdkaxLH5G9RtggcYuc2QIWHwJrvK+xDxln7F5yZrgHYXV16HRd9vjbJ8CjOMZ5u57lT6ltKCEBQXvGX5jDZj7PkA4ngWQY16z3thXSezVB5UAbNlTH1Uif09CXPZT22spy4BnfX3+tU0Eu+fsu795fgqUgAuzerIzj4lmh59Xy4Ki5FbNAELmPecd2rVdwWrORZx5OAuiCHBTGLnB2HQRT8zlrrmjWFcMiFWdjKDVx0Upzs2cmThXoSjzJiX2Td7JGcJ9AQ9PC7CYFwgREZcCwb3AAEcgbwECTvedrBXiWl/+wfJQbv9yfi9UhynDXGxZPcft0zkyUw572IQsHhKsLOLaoCvQYqPSSLsCMSYFLKwdfWw+k8umvtp1UhYf++XKqlVk4WOysHjz3//l7cTXeOKW+w5PC6QYbCyOxYvPzMzq83TrdOP9AmW+Xff3YhXSW6+6bKY1rcn8prbCx6v/Ewa8DEGIIpgTKPJu9f3g+NxGNayl0Buw+WBccccExk+eB63jfQCdmaOX4+7wYvTzv3sKeAp4CngK3AAU8IDFDTBIvomeAp4CngIvIgU4+COMQjhO4GU+cdn0eVfZPS3QYkNuoapiyCouSt6o+whLEeyY2TkCUHORZAJ5mgcjgQAJQAMhFFrgMFQIiaiTuAi8c4ZuOUbfDQAxYT7lmAasCfRNA3GolajEfbtnsR7Qlh1qM47aagG6rVzTQLMg0/yN+b79Trso09oGqGG/8d0CX//RqH9fSUNH/YJZfUDJgiMayMLvBpjw3YAK+lfui/Fo0AnGjN+gNQzxM6N6ECabNQe/QX+ABejHMzClpq1v5ZWFI/TNABeKvEMqd+93g5V5t/AjE27tb/7OpcsLug/wgSsvhNbMDXNtxfj768WhgAlrbY7yNwKSdyghaGU+3Tqqivl6rovxxoqH+Y+AyQQXCHkPKiGU/RolxpR7ZtFEWWZ1xPzioo4fKVUCMPY/K/2JEvPGAnsTsBsByHk1gL3A9jyjNbota4oLZSgEaKRy67Qx1oiPyHpiI3e51l24olgWuHpS6IrwYNof7FEIix2ysjipBX5Qg7G60eqvCtBYbnfTDVlhdKbGa5cMVpQahJXZP1X6v0f3sLj4KqXh2n+hsSxGQlLmIfsp+4pZ3QEIAHDbXs77Bu1fA1/5/mNK7K+fVcJ94ebLrOO4D5hhF/s8wB/rgz2cupjvm9WXETZircb8Jo7Pf1Jiz+VdB5gHcMLz0IhP1oB9UtYNbY2heWcKAMXt+2eD5dVOuLTSPgvOjKyAzkF2f+tyKDACLnjkWllR2DjbeYhPzmuscVPU4NPcU15O927YvGjuq/EWI4rvnF0FMGhTWgoELoRu/o6g1phwzzamilu0e6B4w/mRvJyREbrzPrf9bV2C/D+Tm6X5qDK4f2yqkywf/uKQI7yXmyh37PF5WTx03c4DS07AgVt+dsrJ1ZIsIC7JuuJi9Gb/5FzMntbL+tHuznotkisqWekFTq6bWqrzhOJLjJ18cm5OYApn9wmBFFim0Y+hco4AlHtkffExubN6tteuLPZalb9RG5uKYfEyzWL2xdFV6Kxa1AXAzAm4CBQvY1Egxs1RpSuXWlWXC6gRECJgJvhMe6V+QiDHLrm/qgrQmRFQstiYyifueWf/2EP/ufLhtBu8eVPn/oX+/hslgGkPWFxs5P3vngKeAp4CW4wCHrDYYgPqu+Mp4CngKXARCsCQoKUNaIEFBO8BBJx73dgdmesclDZWpePG7jbLAz4xgYextXgMJgBHAGTWC2ZlAKOEebxZPhzUd4RMZr5u1hM8a66dTLhu7pXKgv6zwhTlt3xWhjHbJtwCUEBDzgARAwb4NC7QLCZoH/exBOEZc89g5CsLFcj7n5UIyA0zzzMI3GDqABpg3BD0mzB6qE9WqtP6cK6+UB95EaTRNuiCUA+/vQj29ivBpDFeCJMBbAxQGQbz1GV9gTllPIwe5XqpA+EzQvEPKz3gwtqq6zzRVYD1u93xX7dgzowTklXK+i4l7gNg/MWoLv9x5RRgnACbzF0ZgtrvVcKlhF3MIcZnM9NerhWwgovxxN0NQlrmCmDWPxyNneU3F20GMpbLYZ4gKMbFjl0Id9+qxJog8DpzHQAFgQZzAa37ayJwKzd8K34fCYYHEiCvN+qVXl7kmWJbLDdqySAJgoaoviQLi2AwGKzlebgia4qDg0GP8ejr+5ryAnhkp5Zblz0+EqZ2BEr8lsoywOJBfef9AIB2WdemwNjsQRa4FRCU/ZP5tqAE4Mp+BEhhcXhYC+zr33OOSs8FVlysbRYHyKzpzicNNECeT6zUmPPk/WslhJOsB9alWSDZ/g79AfNYH+ZO6qwG/SggeHC9BrXXXAtnJuthr59FtWoUnF7tVOWarNaoJx2FXBAOVgx+8QOPDe69a09eErhfjOb+92tEgQu4XbMzEGvRYhtx5uHsx3mC382tJPP4sveQa9TlF6NaO1Ox7lEEGV7Er5Aw/ej+V2bFxFwRxtXiJdoR2B9sr0CADvDP+5hz00CC/y6WFOunxt466EcVCeZXTh+d7EnAXy9TFNBAQamdgnG7fqcytL4QwIGlBVVzTiifH61J1EEbL+WiICzF6M8J1d8//ezUqkCCbkOxMxQge0MBvqtLh2YitZMYWZwzOcPzDCAx1g8ozIRqW/3Y53e+QX3fr1atCFCRJaBieYRupza6J8Ikuy2uZATjdnJz5bqtypOK7H24Mta/b2Juw62dbA77GCeZC+PsvuZs68/V/1D5M0EY1CtgwyleRvEpWbKsrAiuL7mFoq/s3eyzObFG5BZqO83NSxlrn8dTwFPAU2BLU8ADFlt6eH3nPAU8BTwFnkcBrAg48KOVirASDVIEpxIT3V64yfsjF++ouNoBC1ANMwZThrASRg1mtqyhZ241iCGBUAcNVQTrFoQQbTWYLIT7JjSHaQb8oGxjzEy4jhCeMsljJuDmhqoMZNBifkeYRF5AAwSw9AcmyJiasksmnrG2I+CFYUcwRRBrTPkBBmiHAQD02dpMHywAOeXA5EO/d4+eK2uxU4aBKjyPkI7+Ur7RnzLOCrZG9dA2aML99ykhLEagB8PGeCBMpp8APdCEsmDkeI5xMa1ltJHNKsSsUszvMuNA/kU3/83PuFO/t0/jHihmSdcN1hhf+oEQHNCJOfJnShcN6khn/HV+CkiQxJgxftDf4lL8D/pusSnsYcCi31ZiPSEQMWse3DQdVFoYjTVrjDH/KyWEqgieWAu4k2LMmS/Maebfx5W+Y1PrmA+sFX4vAxZkAxzDQuOHlf6VkgXo/kt9R4hhrqI2Fen/fDEoAHAhQTLrd1lxKQbDSNupm5CLKMXidlF/kDeiIFiR75CeXEglAit6RVEkBOV+gfWzl/ypEpYVXFja4GJsKIg/jzDUqrT927SV2YN4jrnCPKRtX6uEMIy+sa9dCJS73K4gbC1bkdnzBoKzp9t75EJlkw9Q3/gjhLu8k3i3sRbpzz9X+m+jPrAeWC+sadaZgRbssR3RbOiGT5/cp9/ntX652hZKI8uKWKBErPkz1u1ljTAKdsZJ1JB/mqUwcOvZoMgEYHQPHjm9/tsffSq9HFdjlzuAPv8Lo8AFwArOD3Z244wA8MfZAQ38P1TiXcB736yGXlhDbryneTcjtEdIz9lxeEW6e8urB0u7X5pVBVaMCcD4gFY572cUBFAAQMmEfYG0ppgPn83S8AG5erq52uwvyNpgWRYLj8pK4f39dqJ9JDhbNuUDUsgxk5IZPeplfGFR/MXACgNWORuwFx5Q4tzA2K7IouKP1k81T03s3JhWsOwD3fVqa+X4xLLAA/Y7U37BNR57NBfnAubNdwhcOKqTwoSAinpcHQSyGjk0uWvt2dp4N1BMi+8OwryG1YisKtqNyU536qbVOxSrokXcjtbpuss3wsWgOmDOjcntVE9lLMsFFkA1tOP8Xc0GweOzN+eH10+GcpVlo3D289v1jZhq7LEv9D33vML9DU8BTwFPAU+B65cCHrC4fsfGt8xTwFPAU+BFpYDiViAwhZnBjB2BNJwSAhQ+T7n6gd2uv7LuarfC7MAc8Y5A4ILwEwG/WVYYyIAQxgQ0CKC4b+6VEHIiqIIRogxYEMo0F0vlGA70k98BBGAEEfaY2yeLx2B1llk68uO6A0CFsnHtAWiBEBc3TZRR9vNrfaV/0AEB1kElgAuCslKOgRW0mzwwfb+pBHNqWre0j3bSF8o0EMSEdvSnfBl4AKNVtr4ogzXUCy3RcKNd0Ie/cYOCUJv70Jj2WDmmPUy9Zq1CWxBeG8hAXymHeAYwh7gvIE/igmSPa9wxcPFk1TVe0nRrDzHOFgCaNjBHYCofZu4ojgX08NdlUGCkbc74MJ7MZYQiCHNfpYSgwIJhW6kIQmHgCYT8tBKgBRdjyvgwdhabAlADIQVjBkiBNuUfKDFOzDnqQ+jAd4RT1Et5zFncUH3jqDyr2z6xsLDrp0rff0nfSZRhbkQ2P3vD/l2KMVEGEs/25yIunV7UfhtoIasJabS6nsCJE2EQVPJBcULfx0MXrNZryWqW53GaZk6gBfst6zx7AS582E//VyUDLBBuIownvs/5LtvzEIqxJwK4vmb0/ZP6ZM4CVOB2EBBs877/YtHNXPJtLq98f/NaO1/dZd6I/dPAacBG9sX/SQmw5XVKBiTyHgJgZp2ybtk3AVEAfCmP99NBJVxP8b6xPfzF6v9llQNYMTleixUPBfo05UpsJ6BFGES7FQzayQ3ZtLTLNySgzLNB1lrd6B1LFC9FoEXHgxaXReprldmUO1iXCIp51zA/EZoz5lg7vVSJwDqcz1jrvCPYQ67Epdy16ueLUS/nMN6hrGlzxyivmYWE7eHetRPhoem9WVMxLaApaxhwA5pxjmbPPKVTHYDGkaQ2UJyh8LjAgD2K8UDsig25UrpFLpWeA1ZYoy8AUJzPEux8/WWPNsUDO/Oy17AHf9toTJfXF5sfevyvDmitB/dILWbN5cFBfeZqP/sX+9Xvj+YIZ072avY85omdT8cVvPvw7a97uitgYkEGf+2Nxc5ntE/sVr87srDIZ/aucEaZFRDyrKw3Pqd9ZKYx1c4JMK7YFo/JtuKw6p8qXFDDSRRlK8/+fa8Y3B5XiseOPBr97aAf8A4pX1j7Ap5zHvaAxflmgb/vKeAp4CmwBSngAYstOKi+S54CngKeAuehAMzVu5TQEEOYiZATwcoZkGHt4b7b8VWxy9pVcWsmCIU5WFDiWRgY8sJMweTBDJvbJQRmWBxgrUE+tHUR9JgmOEyMafAhsEG4ZVYHMH+UY9YFxmyfz4WSdc+EX7SN68uVENwbQwPIYgCHWUqY0MosHYZBEpX4pBzz2U/dCPjRPuST/Bawm09cQZkg2uhiYE3ZuoM80Jo+UYa5zrI+WF6LD7AwqgeawERSNs8CmEA3Ln7jPv3jMnCH79QH8015Jnigf4APgDDQHUH3vOzzBy4c2+uKtOsmXzMjwIK+0gfmBM/SbhhXykSA7q/LoMAIrGCuMK8ZK9bG/zaiP6AaLpe+qVQkYNuvK8GYAwogcGAdQX/GhvG3dcin6SGadjna3rY2KdashWwOMf7MJYQyCDgQVtEmNG7LcQDO18vv1A8IQwAxmA9bBrTANY51evfceNBsVIqNdj88dmp9CDC+ABDgfLS86H3VyRrsq22sX9trmA9LmRZt2uox/ubqhTzkxzrjnGVfIuBC0Gn8hQP4ApD+oNI/U6J8u2xfNqCW3xCCEqeI5xDOAbDSPubVD1y0s5eXAS3g/xc6KL1XiX0KgStgAePFXmnCO4BoAEAAE7P+uJza2C9Zdwju7KJsK5893VxVvWWUgTawPtmneQ4Qkvy08++VeIb1NwSYlK6qgBiwYqxeqfTTQV0WOpNyM7ZPgtObE8VJSZJgUq6gEvmCaqZZFuk39pajnW460++nn282qic8aHE50+ea5GWeM9eYuyg4MBdZy1iDsn9bbBreSbxjcPfIeQZwkf1l21yj+BXsY+xf0OjsJY1/ARbBR/pttxHFbkHWbaxvsziDvrxXzygiyEZVgvjbFbz6IwIr3iaQonbyibl92gjeLbBCqF94MeuJc9G8rKRzMQBjs5Uk5XG+XlBiv+HC3d671BaBCMWcLB12RlH+tNxDfUKxKWq6z1mFvXMzuMJ5kDMlL5aOQJmGXDtJ4aXoCPD4c5Vzp8CLl+v+vKxJ+vo7iuKsL5ocnamlBwVwfEEWFROyvmB/XlKw73m5hzqsNnB+oGyUOKqhZu3s/vxD4zvy3+qsRpw7y1bLgMDM57rGbM27hTrXdPH3PAU8BTwFtiYFPGCxNcfV98pTwFPAU+B5FJCG/Lo05dGYRfiJ1hTCfZia3CXT0276DRU3WF+WeyDywBwAQPBpmv8Lw7xnhCy8PxCwmtDSwAYEMuazHAEpjJZZTRhoAIPI82aRQVvNaoHvJoAvM2nn0no26w7KgtGiDIRElAsjicCMtporELPWoA4TupEPph6tdZgn8vMcjDv5YeoJssg9+kV+nkUQZfE7rD7abVYo5faaUJF6y9/L1iLUS332XqbNtIHxgeFEaIbwyOIXmE/2zVYv1AENoIW1gTFCuIf/dVx0mfVG4cKqyo06buL1Yth/VlrAcjxzxjrDxp25spO5Q8H+ujQKlIIMY/XA/EKoicAIYIw1YtY/zDuAKej7QaXPKCFEYr6xvhh/A9I2O4wog13na9hmQQd/I5TmE+1L6v5jJYCLW5QeVEJYYO4lNpdLjIyvUHr7qK3My7Iw+3ztuC7vW8DhvfMTFQltI9zjKGj1QNYL8rCUR/ospP1Z/OwfPZp971ffbcDol6Qv5wMaRvQ1IIp5Y/se7TBhd/5CQRXFKCC4NmV/nxJB15m3P6T0M3f964lD+mTvYu9g30O4h2ALIZk+sm4AACAASURBVCfPLCjxTgFAsD3sPS+QUAi4EKZincDeRxtYO9zHUoy+s7exF7NP0T7WhO3D7KE8Rzwg1h37KO0HsON9QZsRVALQsPdjdcQ7kf5QHsJd1t/l8kqMFeWwV/8LpQ8p0W5o9SYl1gx1otHOd/aA/mjP2LzG9dOZ60V0GRVocicK4j5TicNmOijmFL9ih6wsav00v6WWyMFL7hrZIJ+R1cVSrVaRILOQQDHMuv0sH6uHx9//qSPpO+696YZd92eJuvW+sAZYD7x3WJ/s6VhWACZ+Q6m7nB+4sBYAHEcQD8hY3ltezDl3vVKatc0ZjzPTF62xtIIRoC/cO/jduQP5q4dWCGfoansI7027dmrXOR4qgPTxx3c+KMH/bQos7QRaaNkMX78KpH3Z3efszfoya+NLcWdXroRnARlQ4inHr+oKKBiLa4NbBTIEY9Ode+JqelSxND564om5B2UV8VZZP5yrtez5WD2cUBDto0vPzGQTc+uZnn+VXENtCPgQgOGmBX4c0uuyq+/sp/NRnO9RoG/KywRotFR3A+sK5bEzNCAJYHNLzxxsnw6eFi336vtzYn7o97uVAIx4B3xYyVtZXPaU8g94CngKeArcmBS43EP4jdlL32pPAU8BTwFPAaMAgpN3KCFMQasOBmzDzX7VhIsme679WOqCKQQpCIlIaKjC0JHPAA6YDRgiGDg+YXIPjsqE6YWxgcHjHYPglfyAFwiBKKccXwHGGWYMxmWozTxqqAla+TQBlIEFlsdADxPem6UD7aQOhPQwTtwvl2tCfpgeBEbkg8E3F1nkRVhFuxBY0Xbrq1mYGCCAUNnic9D0MiBRBl6sTvJAs819oW7um9CNTxhoowljRRvNRQmWK7TRyjHBJfmhpQEy5p+a9qLJZn7UEZKlLpl62NVuesD9/+y9B7hl2VXfedLNL4fK4VXnVtNK0MIEoQZJiGSiDcYIBGb4ZhhgjAO2sTEgjwkmDHg+Zj4bTBhMkgkGCQFCEmqpW0gNkhq1uqWO1a9yePXifTefMP/ffWe9PnX1UlVX6qpzvtp17zv3nH32Xjucvf7/tdbuLijfmLpZGABkQlvNKOEJcN0PgWeDZTAQdxCUz16XvUbg84bK+BWtWwo8AhLQPgC7b1MCJKWN6EsAuyTagBjijDfKeULpaHoN7W39vl/xywQsNyI5+p46aTkBRvDMwGOCa9l0GSv5L1aCYDEvnqyMOPcflX5WCbCLPmb9L3vdy+G7e+fhyaBclA1oFJNqnV5U0t4RXVmhO/K26K3U24pe4TR/8/3P1I+fWSbk0lWp6zYeEHhObGSNf+lQ2BatwsbKIi1mdQmkdf9w4/A/rdz3jd878uQfMTcQWgaAifkKkgsPCuK6M8++lOPndTOEqr2XGAsG6PMs81hgbrN5kucRcol5HMDRSF8bZzZXIiPG2ovB4tfGGyCckfN8sncP+T+sxNxHnRjDjGXAX0hHA3p59iCpx9jeKOwUQBuJA0JyJq3Pn+qTehKbHa8Re49lvePS267MhxF0CjUWB4EvT0rvkHiIV7iOp8hP8ZT2SznYC2NtkaIwUa4bFgpeXabhnn4r+AVvOk6SVXlidERuLKif5BtxX5lmuVK58P7G2ABwl7ULc/v3KOFdxMH4gDRj/HLQz/A+YtzxeRFZcaUKdaPmk3pXMF6pt3kSX9DMMBVopqhNxvWRXfE97br7d9rD4n7X78uVUFqsoQbfi4R/CrSh9D0LJ8e0yXRBwY62WpZsKxXWlLZ2HswI44aN3svZTO29YGE8eedDQO/W2K6Xhzqu9piol0fa8oXw9xGuqTLS/jNtzi0PDPd35Q3xOhEvhK3MHlpDuoe0H8fuxkK1Xij1Kro+GYrcP6yOt0oiISItr+hfGMUwZ6I7MOdiIMFG3exvd0SfkMXInPmXPSlYm0IALSr81tFOyx3XSiS7XrYyIHvmaebJnLDYtgvlF+QSyCWQS+DmkEBOWNwc7ZjXIpdALoFcAjuVACC4EQgoFbwHys7wAwUnXFx2Jt+yz/GLKBMARwA+gOQoCAD3gNhYf8+kv3HOyAuuwfLVXNMBtwBdUbpmlVCwAH9QnPgNhcM8FAxIMk8FPlGmbV8G6kZZjACwuloIJgPn+eR5FioKJZznrtXxxbAefYuv9FrqiXJvZeBavhvJgYz4O/ssysazqAMAAfkZ0WBlGzxHfgZ0GgmTVUQtJA2fyN/ys7qZRZ/JwPao4O9BosfuJR/bewSlkDojfxRePicdt/gJp3P6bscrTziH/uWoc/znqBt1pd7mIbNZfHir6xX53ISQGMw7S0BYn+CaLMHF30aY2TV9y+v0GX15XQ3yIiUBkDUEBTH7+Y7ib5bpBmpCEmD5DeAKMMvvfKLwZ9vzish2o0xEgNg4YBw3VHbKAAFHGbDKfafSdysRRm7weFAnGBeEh/qwEuDEFQXPr1rF04wV2sZbqreFv3pBpVIYUdibUYG1I+ojlZVGpyhQtqMfe7JEFxjlXBBoe0qhohoQByIXrrl1eUpoXHUZ7/3Tf1o/+xU/878nQen/RVSJF3yz35ijrzKfsgk1c/1rlCC2LvcgpNOjSnen/e0P9Un/B8xiXqVP0g+NYDWSwvZ+sHmP91FWJtyXPWwOG5SbEcsQGWthXda8HszbifMQcQYaEhYQbw/zKIGAeDDzIMYLZAREJOH3siGksuVh3jUvOYhMC8PD/dxDuEaey/OpS3bfo4GqXf6f2o+CsTut0E9H5E0x3e72JjSBFtTPyzIHDyQsP0qSbtRViCg/ng40GBQSZ0xW50G7GxfipPN0u9NjPXDDgNxbeCghqP774aV6IV2+xF/6nVtsek/dsusHCAr64RuVAKntoJ8bWcG5H1BiDLJOu+bz2UuXyEvOgTGAQQF9GFm5kBXq545fkvNp4Bytjidj2mWhoRnmXfqdNREJMpN5hTmDsQyjHWi/hrr2cJjqrJYchUZ6yYVL8ycfWw/TxqTtyAruYd4iFB2EBWuQ13FSYasc14/vKJRChw2xO83CiV23zTcnDi5+7uFXnzy+eHp0VRtzv+7881Of21yuroWxUhIZ068Pf2uT8NLiybF5bbg9pn0rXrF0evRju26/8PjY3uVZ5Y88IHrRBT6i+/ZIJo/JK+MDxUp3WF4WrC0pj+0Rx/z3ghLvk2p5RNGzui5z4XuV8HjLHrRV35NOZJObh4UakE7+Zy6BXAK5BG5SCeSExU3asHm1cgnkErjxJLBDC3FUhIssqq4wsIpVKMSBAUACftxVp7R/1Bm6b8QJhhuOHwCcUAbCaaCUAQrxN+8MfgPwJg/+Ng8Lzh9TAnBCqQD45hoUGMJ3YI1L3bD6wxoWJRHlz0DTrNINSGPlM1kYiE/DDnoncM5AepRQ7qHMKEFGghhYz2/miQFRgeJkIa4sHz5NSbRncQ6QjL/NTZ9nUZ8sODVYbu6jvkaEZIH17LUGqPFp72a7Nkvk8B0lD9lmQTgjQYxoMXmackgZ2CCWewHU8LQpO8HQg87QK2tOb7ngeBVkDEhmVsSUj+fQZ67FMWhJaKAidTKvFPOeMW8QZEB5jYCyNqIu5r3Dd9qZ3zhH3xQel1xksb7TcbYJcETZIeDI/7ASYZUAdK2dDDgCsEQZNwty2sRCcfDbVbHe32HjIQ8SABZgJLLGAhJA4Qc3yAOLcwBnNu9mrqCPvSwOyIpON/LbnTBodnpjpWKwr9UOD4qUmKmWCy1tZp3o797oUHBmbKTiNprdssiKFXldsLdFR+Bo52p5WlwPAaZE29qY+vivTxcXnj927NvfuSKEq09Wdna94ltqxx4ZFmIFgX25B+Ao1tzM748okTf9/xkl3h3Mpczbtp8PfXGdvBPBdjmg6mbkXzavnupPmXg+c529S8ybjrHNWGCe5zfGOePjISXmFsY7pJ1tOM7vEDt4ngweWGlnD7wY/5MSoVsgiLjviBJWyXg9MTfwPl1RGY282SDbnXlgpZu5C5N1i+rjVbEQfaMBHWXtXSGyLr6gH8fjOBZky5hOptzYva3nxGWxvR2Bt0GrE4rI8+a1BzHyumEIi6yHkrw/3GdmL7jDtZKrfWj68tKnm3op9f9+OZMXtJmSvR95x0CoMZ5ok59WynoCbdRfeAcx1njfI6AwJbA37Fs36UnWFaxLeTdDzGsgaALUqA8Kig/oOy+Uask9lRGn6nrucfX9J8JuMKv9G+6SuQOyfrX2aqiFPb+9eGrscYH8B/TpdBq2tc9lSY11AXNClpRgjNlazwxYtsuceZVrx+TRAPk5JW+KdqEYtbXHxPnR3SuuvCoWSkOdcHzf8l6/GO3RdVMTB5faQTGaaC5XWr1uUClqSSgixum1ik4Uah8OeY2Q5EHSPvPUnkCkxfTIrtU36e8DIieOqpQLyocQk7fp7wntjfFJERZNhZz6Zslq2C/E49rDgj7HfDmjxHyIcYc2+nC91spQ2F5NJuTWN73Bph+EuHqTEu8L1hv5kUsgl0AugVwCt4AEcsLiFmjkvIq5BHIJXH8JCBzNWoZbgQygNcspzgOk2LX87elesyYdrEhfiRHYcCkVBJjheYD1AKSLTmG06sz9CftYtJzigcd1DhAS5QClyTb0NXCeZ5lXgYUxgqQAYMGL4ZQSgDjPQCEGAMKVm7JivQ2ogwKGUmbkjIHs5G0AtG0ubNdkw3mYu7iB9FZ/U+YM8PqQfrDNsrFcNe8E6k3dAGYp++BhIJeZydm7kvMGZqF0AWBZuSzvwbpk68T3i9o2fbDV0T6tvY14MdDbypMlK7KkhoXIsnP8bRbCyJzwLVhKmwUzIaKec4LJwOmel+IY+U7p8LDTOYZVnoH9tk/JBmK6tFObEHbWZibbrKeKhbbi00gs8/yhXiSAGuQFqAcBZh4qhA6g/rQT57kGYIY247vtD2FtIv14nf/JEkE7GV88kzISCs3C4xgwyfP/Vony0H6Ef8FzgfYA9MTTgv6Y3ECAkZEmRqj9nspHmIcv2aDFGV/fhVwFqDLeVm+gemxQ3LVTIh3csZFyIF6iGkfJ/kard0TtLwtyFwC3Kq8LCK6Rdi/aPVIrPa3fpuR90RNQe7JSKiwdOTC+cjOQFmoz+i5jnTFCHwW8G6/NfvgfjXz6T5ZX7vuGPmGx9Nq33Tv22G86Xq8fTWyrgz5tVtyQXYDxvAcA5AHOGIPML5DYfDKuba8hIyi2e8YV/50+K1kw7m0e5/sgGM+cYe9qCBbmfv7mfUd/4Z1J/RgTvEd/QwlA9P9Qsjl5M+torIkhADmwTjaSlvkDWeHBhPyQ5UsmNeU11FFfP6WQT3vkRVTt9aL9YZzs0rlC7MQt1/N6onRHFM4+1BiZdOO4ppfqU0IrJ7zIva1cKl+olopntJdF60bby+JX3/OU/4lPn/K1aiqp7LSP3+2GXrlYiKrVQksNEc4vNQmx9pL3fbniHXH7DM3ggvcNFues4zDMoO8MelRslNuv6uQ7lMwQgfdmXf3/Jfep7Yt+w13BGGdNxL5M/RGKd4V2nOjvX6GQUJVS1elFYTC6dHbooID3RHtTPDg81dijXV7Cdr28UhltOfULQyunn9zjy7ug3NW+FZe6X4X89/TQZI0McNwl/cd8kj2y5JN5wG4lTOYeCAvW3SIIkncNT6+2d995vqeyf0rlmxPhElfHm/sL5R4eVIHqzlxWCArh2MjulWWdP6m6jcsT47TIi9etXhjC++qTqnMscuJOlXWauvY6QSS5fEJyuVfkxPv23nX+tO59E/tZKLRUJPLmyz0v3rd8brhw4lP7jo3tW/705MHFT5aGuu8TgUEfnKX/KT9f1xZPfur2sVJtSV4ujY+EneZrk/6Wahcd2VBZF63TbrjelRcol0AugVwCuQSuiARywuKKiDHPJJdALoFcArhLr6+fs0QEojGA3QBpi5vLb1wLMGIhYwA8OMf8bF4FKBMWs9VAa1vJ67Frjts7JC7YeNHCHAGGDDu1ezvO5FcWncJk0fGHCCWAImGhKADwDBw2zwSzTgWkMbAJIBlrUAAZQntgwU8dAMWpL+WFHDBLdKv7Rl3HrOkNuLc9L7jXNtVGUc9am2WJAJ4L+AbIioL+tUpY9kK0kCcWrFxPeZCdKYGD1muWZxZMNxDXvCo2ilmerZNZ/GfzMqLFSBnUZKurAWbWhyhzlpHaivgaJDz428JbIRPba8BAfMikScevSlZivSbfUnDaz7ecs8doQ5BJ7qWv0GfY2+BKHIPlp+59ZTltB8wT+W5hyfjbNo0E4CTkGH9DpCE/QBsAUupGvWgfAD9AHABE4tJz0F6QA1igAsIa2UYeFhN5fUzp3IaW2Rt4V1Afi8EMYUGMf8aMAZuMGcLMMB4gyP5vJcYHZeV5Vy1efVrvl/rBeHtM6ReVAEK+f4MM36ZzALN473xKMoK0uKEBMHlLuOVCUHZrzpjC+R/udHszinqjOcUda3dDgTie6pL4vV44ttpQPP/Aa7luXJMVes33k+MiLjra3yIS6Nl7mVtq03eZByEq8BRg3Nwh9OwrJz/6S44Ii35zd6bvcbpTdznlsxpOff58/aD/QlKQB2OPPU0A15kX2ZcBkJ+/AUmZbxjXXGcE5HpGl7lHywbd8fJOZZ6/IRCWEhrmhUQ9eC9xYPHLOGd8M6/wLjRPsD/X9w8qsUk9e8JAOECybmSGbe8UPnlHfasSY+rXlJjvmL8eUrJQVUbMX2qFZcvsxiIqYmGzDYH6XZEVHc912iIrhtS8ZW0gnMSeU9TvGh5ORQBuot8rvu8XReatlgrBsMJKDdebHdYrl+P5cqll3vZ6eVV4J84uFxeWWmXVadj33TGNVzeKk1j70uhr0lptdJYV3qpVLgU9eVeFGr/I8Ibwttgi5BNFNG8K3uO81/Dge70SBiIQyf9wWwGteTFBnvPusbBjyy8HgnkHdbukSwgplMqUtUR/vw+dGCpWtHmCenOv7Z7oNt1PNJeLhdby2GuiyL1fYZ7KCodUUdikpcZitVg/P9SrTTbxKvAFwCfa10Fem4oq5San9GmhUTcqF/ML819Z3gZOsdrThtQ9X6GkLsSx29X+EVvVZVvcRnlOizx5hcpxUOUYrY62v6E20ZiSZ8UJPadUqnXnRBZccP1kv65h7QMRyjpqWCvNaXlBfLI20WzsDc6f1v4WyZ67zj8roiLQ/edEUCw888jtp1T3/cr7i5PQi+vz2sViPnnN0pmRr9IY+4X9952ZVb73SZ6j5VrnPnmkVGrjzc6Zp3YfWjk/7B/9m8PHtBm3e/9bPnNM589Irt2nH7l9pLlY3d9pVO4rD3tj5eGJx5fPzsqjpf05GQaI9wj9PbsevqR2zy/OJZBLIJdALoGXnwS2ffG9/KqUlziXQC6BXALXTQKDRAXKgBESFqoIZQWAFSCQBDgBiArAw3kUaBQoQA+AIEgBAFAOs66zPDlHfgac7MTiiGdZ/FiA27ZTua/gRAoJFHe1CadvpAPPBIgAMKGclB8gGPdtygjgQgJI4TpAbsAYLLsAW3DdRimGAOE5vG+MuDHSJUsyoJBbfTi/5v2xZrEKmEYdyQ/wF2UvC3xnwWUD/wGUAIm5jtAaWCBSVsryfFpeiBmuMyLD5Es5jFQwxdaIB55llsDUw8qdvd6IDysX9xrRYZ+cy3qNWAgjk0HW0yAVzbpHSlZu9lv2HN+tT1kZaSvAQ0A1FFSTqazrvOed9gu7ULwdf4LraV/aE/nTV8jrShx9a9c0I8aGeaPwHatkI0kAP62vUBbIJ8YGwCBgzUymbPQHSDHK+YISzwAYpf9CHtB3OU/+jCviOvNJfrQP/cvCZtEegDlZM/L1MbUJWcH4xSOJPsSmkpQbLxYLuwaJwW/EtycMAm1AWY0Q1Ncb/mDsPaTE+GMfA8iLwYPwV1+RyvQZyWr+RgXCCBdz5ny93IuimsDLPQJeJ8X5Don2na5UiiWBs0Xf82sF320KfZIlurdfoMnp2HHPygJXwKdTbrS6tVLRj7Vht5FON0QjbhPnnjJaaDqz2gWwI+Y9YDrsRAqkazODs084u//y3zbOfflP1rSPhXP+y37UOfh7/9iR3Wy2rowfQhnxnuCd9VdKNvfwLEAmxiN9nsPmxJ28q24ImVohNiBUjLmx929/3lAbMMfaPMd8BMjGXjWQvhZa6pf1/c4dVBBPRPbCYQ5jzqJ9IIJ4F/M+Q+40yKUQhG6n0wviKC6qf3vFQAGiEkV8iZJ52XlPaBzoHeW1Ze/dlMX3UOAlETisQkKVBFsuiADodTphUcSGSAvPgyjQZu2X8vwdVPvSLpGnh39+frUUhvGoBuhEGIdjIlgmxLbIQj5ORLokJW0WLkBVoa00vyduU4RNvRdGtF3vBve2oC8xTml/xhRrGN5tJNZjGBRsdTDW6G+sMXg3QeL3632jztGX1vqXdbWtl9i35of7OehMaShxChphldHkI+Vh3z3z1ORQY3F8RPs+VGXScUD7NWi5FHdEChzQfgzd9kpJ/xXqCp20oHMQD1GvHRzX9tNZwoL5b69AfPaQUMi1hPVHIs8ELbfZKyNKtAn2ksI1zSr8UtBaKclzIbs03LR+vIsPKRFGinXRCM7WIgGioamGXyz35pfPD1dVziFtqL2qZ7WL1W5Rm2Xfr7rSj/A6pm8xlzB+maOXVc79IjOGa2PNukgJ5pcJhYlqqrxFhZAa23Pn+adaSxVV3A/1u3YXd16vmpVEPBw5/dTumWntiVGqdfZ6QXw7zxMJk4ztW/EPvvK0c/yT++/qtctf143d+G9+/zV/LHmd18bd08o79UAlfFVSlFAVosr9HIywMoZgti5k/4rrOt9cVo/Lb8olkEsgl0AugcuSQE5YXJbY8ptyCeQSyCVwsQTSkE8GVDO3mvUjwK8RGYANAJyARWgkKKAAmwAdnAPYtM2hUWpIAB6cB5wAmOA+gEMDKQx0xdHCYvJfBAYNeF5YSCYU4DXkKVoIHH8kcpI2ADWWVigxfeUlLS/5AQADTgEAcx8KBs+jThbiibJSNpQc8kfBQLmmTgZUZYkGUzqyYL9Z3/IM7rfwIkboUGKuNy8B+7tflfRAnpAUyO07lAB7sADneYBp5IkckamVwQAm81KwT8vTiAaebdb5G9WF603+5G2x0c0TIwtkZZ+RdfvnvHlakF+WLLHfLB8rH+dpB9N0bX8Q+51+iBINcP9LSrQzfwN4HHXKt3WcxpM9p3q71Y1yk4eF8bJ8Nv3cIOQT11JOKz/jgnrST+gXRi4gW36jPLaZJX+j6PMbbUeIJdqOccV1RqgQ9oBnUB9+o49Sbp6Dh82M0seVzJKc66yOEDeUAVDQQmfRf7Mb9Zrni05fdFg/IH/qglzJG+tpxjR9b1aJevAJEUjYNEg98n+5AbZ97wkl5qTfUfrHgwLR3z+ihJX++5R+X8Bt+0YDxCArzi80ijKFrRLqptHqHPBc96AszsdlOT4ig+xqwfdaYRgNVSvFrkDdTiQMSyDokEJCjSp8VFvXCfXx6S+hznWUZyTA9rq35zYW2vR/IwlpQ/oqfRfQ/MeVPsvi3w3bzshn3lUTYdFv6tU73uz0Rg842t+CPwHJCG/G+GCcMt8yDvEe4j2ybnWvPtC3Yr9VjrTPD9a5q/aBaDDjA0JAET4Oougbt5ENbUT6ciUI159XAqCkDxIuinch88tOPR1iwpsViwGeEvO+646LqJiPu71inLg9fSdUmrp+3NQkFyl8VCkOk55YDT3HFfwfewqhNqINuxXpv8D8dhGDda3bGcLk2OmligiIcREWIimiIyr3Qe21sbvZ7g6JoFgIfAGv2qdD9vPz2rdjtVj0Xmh1krMay03tW4P8jFC71sXf7Hm8X0xHn9F3DAwgFukHvGswCDHPQ8tjcM3Ced5xv630P5RYT/X7y43uAXcNGgH5MgdePO9JgkPioEf3JntFcS01l4eqq4tVBWtyRuRhYBtQH4BoGJpoFpvL5SmRFW5luN3UxtIfKhc6/bXlQGioY7peAH7kiJioBIUo1L4XIwqt1N8zI+oGvbDjnwtK0UJ7tfiKQlXR2EJfnh5mC/NZ0jCPYAuPyTuXtdEnRZrsG9ldr04cWJrVs47Lo+EZkQfjI9OrQVDu1RXiabdWzxh5WHg75hD6GQ9jPXxEibXLnK6bE3nBuQnfjVZU/76Xz4H7T1dbK+VfPvWkRBS5zGGE/tM0kszLO+RekQ/mLa53rLuSRN6Q7vWrYy1XhMek5LRHe4GMawW0Vx4rkC4YNa3pG/L48osVdKRFhYPSZudJto//gc6ztnDyTbevwQjJH5FLIJdALoEbRAI5YXGDNERejFwCuQRuCgmYVbx5J6BAolQA6lhoJUDle5RQ8m2TWgBTlBDOMS9jNYXiY5apALR4LgBSoGwQmgXvC4Ans8znfoB620R6MwskU2oBN9buLYyp3FHoeDXKAbjPc1AUKDPKByAw+aK88DcKkoWxQrmgHig+ALdYlKOEIAuUHxRCygZInAXh9ef6fhB850CJNNCFsvCdezmP1SrlohxYhFnoIAP6jTwAEIYc4NmAz8iEjUwpD+cpK+Cr/Q3xYqG3jFjKkhaUi7+pt5WPeylb1gxu0COCa83yFoDBtE/u4zcL8YBMjGgwy3vAeMJ/zPDw9PlZrw6uo32yJAplzL7TzdPE6sIzkSloI/keVJpVAgDBw6biRKsCpQILZ2QAvsk1LcrmH0aMibgwWZiMjahAXjYO6Lu0IeAm9aWclM9IBKz/AP/pUyi0yBBLZdrTyBcLvwIhQZ/EQpxxQdgLCA7IGLwfkDHy5Hn0BeRGf2Kc0X/pT/QVymQEo4VBsxBk+mn9oF7UiTFKHlzD8w+kz6CsgENc814lgErqR90AFq47uJ2tjH3fJiQPMf4pO8A0/ZW56rs2yOfbdY42A9D+WBoe6oaor6yo2YDXk1V1WWDrkMLb1BTXfpTY/ZViMFQs+gV+W212xgTSUiGbiQAAIABJREFUOmE7LjZa4Vix4PnaiHuxUvI7AkFHtFn3cLnoB6pUSwRHU3kyR+0ULN5I9FfrHGOXPk8/pD/SLykrpAIhZX5FaZD4zJQlcYL6Gad85pNOb3zGicqj8rL49+898AffyRzCHPp+JcYL44e+zbl10vxGI6uulpAvIV9kAzjOwZzBHIRX1h8p8b7650qQnVsdX6gfSdzLOuBHlZjL8eygHTYNMWfjO914u6MxsBi58ahC8ye+6+NtUdTcXRaBV5RdcyAwdVpeFLKidtpE2MfDQn1ePhluWz4XxJHyknZYePcHWZpcv2O53vY73bDa6vSmVacpkY0HlA5pXA8nsQBP15UnlbdHxMVI4AfnFezqtN5Vcbnkt3o9mZoHftTu9Cy05fWryNqTjahgXPE+4X1JSEveh6xf3rxFAY/qN955dszqCyDvXyjRz/A4hUTOrdPX5j3e/azPXzzUwePQ1SbTTr1d9z/uFcqv0R4PQxAMUVPLDXlJyHPBUVil3vj+pcLIHq+msEfsP8E+ELH2cajPHZ36G5ERr5QXD+sXvCoq5ZHWUhDEYyINatXh9oo2tO4Wq0Gxs1psaUPrxfZq+YVi3D2hfSUmCpXwTK9ZWBJhsVlb2zqP9bAdrJ2e0I53z6osh0RM9LSRdmd4V/0jIlbuq002ZkSsaPPwhPUT97OW4n76GzLgHGsjCwfK+5t1Jn1umrrps2+opHBO1dseOP6BhRPjD2nvioq8LPCqIxzW451mcejsc9PtI689/ozumdC1Y3KwcCUPVx4Y2hskOaFy3CZiwzyECNXKu4lyyX3FlYeHsxSFvVXto1MbWDigN32xEl4xELS3FBF+UT/N/8glkEsgl8AtJIGcsLiFGjuvai6BXAJXRwKpd4WFu2GNDTAEkA54bpuKolBg0YUCwGLdAB8L/8SCHfATpYHvgBAAoizOOQAyAIU4z3cUChRaAF/AD/IlZcNDbQQUAjYaocKzpZ0tJU7nrNSLr0CJA1CZUeI7CQAYwoQyYWFNvSx+N8AkZAZKDgoNMiBPlGZkkAXLB7/r54u8LowMQJECZCM/6sfzzAOFa1CiUFQAT3mHAdzzSf7UnzKhuFNGgDnyok6fq9S3FkvLSV6m8JhHCdcasZCVnX235yM/8qKuZjHLNdk6Ak4BIFE+2sc8RfT1s55BHZEzoAJlQn7vUvoHSrQvIY/Iz2RPHuaVwDOzRBD9jXpwfpAkoZ3od0YeISvKKJl6K07l7n1OC9H1fzfLWeqHLHd0ZMYCZeBe6t/fuFcHzzc50G/ox7Qxij0y4pl8h/SCAKCPc3AN9WVsYBlIfowlDvL4OiXGFwAE+dOH6KuQUZAdyAcFl/Fo6x6eT1x5lG0INg76Bso7YCBkYV8OqedS1P2ePp9lxA/KPmUg5j9hNrgHK1jQO6xYOU8eH1JC5rTHy9GzIhVN/wM5UhcIIcYM4MFGYW1oD2Tzs0rvTuudzeeqfRcpsVnefZJQ5EJR3hHVoOCPlxz3oIiJ/e1mZyIu+ApxkxS1GfcuDZrS8FBpqduLimEYVnyPwDfeecXET3pRUllZ7Uwps+d1b1gpBa7IDMLixDeCl0XaP2kbxj7jD5CH8cPmsvTP1yvxntnZkSS/VlyafX1776v67aw9LR7sfuA//mJx/jn6OHMWcmV+ZY6Ic5JiW7Hau4RP5iC8rph0me/wniB0IfMkc9fbtsiN9+uXpe1JuDn2mcH6mAHA/LcpcZHmGWsPh64K0ZX3UOj4oiMStyqL5hH1HJ13AxEXmrTitva9lc2021UAm3GFWEo0fjQZxwVt1M1+Fq72cvGuZ0illUZHpXBqzVY4FSXxQXmP7FV4q2kNAM8PfIGgyaT2nOmKzKi2O1EliqKCSIoC+9SUikHYDSNPY7hFHSSbDclVkTzbNux2F+wgXJuB6LQ/ifcd7y3eocy125FZrBv+ixLjm/EIUfEeJTPcSPLxeVErIWPe+etHV4HQGlpxKQLe7qkj8YE4amgPhniPvCKclbkheRR4zviBpV51rFmQ10ICGSGCoCOPCE8g/B0iLCryJnidPB30OvH72y/omlfVRtsngkovYFft4T31eXkhhNoHYq88DUInCYuFaveAvjcqxfZC3PNacezzDr3U436RK08ofNPHFIppsVTtJrd//uxhPX9cRMGYPllbsW5lXcV6i/Uk6yHbO8eexzhgPcUnYThZe9E3uZe1+FCh0rtn+sj8UYV4Oi0vC94v/XWV6nD42CcOxFOHFt6lsFTPq75fGPWCSXlSjBFqbvLwQiLy4lk5Ox3SfEMZTM+xZ0+ItFgKSuUkKJaUX1cyXOcl8KalzRgTOel2qb0jvz6XQC6BXAIvUwnkhMXLtOHyYucSyCVww0mABb1ZswJ6ogwA5gCis8jGnR8QAmCBRT+Lda4z638D+VGgzIMCBQOgyLwuAAu5FxCKTwOleJaFwbH9BrhnI6CZ6ygreVEuz1n6eOBMvClwopaFdgKoBfgmX8Dh2fQ7oXmISc51KDk838BvPg0kt99MqTDPBV2yqZcF9wJGU2dIF7N84zwaC+VAcQIko+xYpPJMSAOzBKNcfAeo435kD5hm1vJczzVmeUz5qacBfPxmoZuywJJ5K1j5kTHPGNxw2zwLuJeyAmqTP22aJT3Ma4T8KBtlpj2xNKNuRsgApNNnkCPX0R5cS50ps3m58N1IC/M4Ma8W6mpW1MiC/kZeJgv6yZgTrsjDRtWJ65STspAfgJqRDpR1yyP1rLA+b6SdhT8jP8qNIoxMqCf9BBmhFPP769L6co7yA/gzpiy8lf1NX6ANZtI8yJc64WkBWIMSTP1oD+pg1qkAeRAa5EcCdKUslGMtJMGL/c60ZMpv4df0td/mPAPwiLHJJ30RZR5Z4tHRD8+gRF+1fUCcmwQssv4BMPp9Slh4A6bZAWGDDCCdmPOOCqiD0Ole5/r3x4Esq+kXNcW1n2rHyYxOHuj24kq729wXeF4Qal8LAZluodELFeIi0vfY8722PC8mOj3FwnGdVREXHYWRKSikTlceFqFSdn7LiOLKft0m5JNZZtPn6duMCfrlG5Xo899/CaXh3cS4e0Qi+ESwcppx8c/W7ncLp77+v3SP/OqbIIMZFzkIegmC3eBS87qArGY+YlzZXhV8h2CaUWIeArDLevWRHX8zp5OY5/7PtF2YDyFoNwP21gjUxJl3k+SEOo/GhqOQUMltsfq5KLpI4aKW9XdbsaGWFBatKOTQl+eCfBKc8/K8ULgWJxCp580tNjYE+V+aWHZ+t8amiuSWwzielAfUNKNRYZ+m5EkxLaKiLsS4oGiZsVxEPJEWuwWUljSGayIhQ32Gbi+cFxGDvCCde3ig7PzpL/lKxi1tSPvyrqXtbT2AJxPGChDr25EVFATjFsK0sWagPub11PcSvN6b2r9kSV3ZDBh3vKeZwyB02MNrbcNtnVEIp8LwdMttLvWelMdDqVTtBEEpHB3ZVQ+174KnjalDhVyKRFK8EIXe3MJJLWsSV6SDv0tJzgHJqsZMf10qj4y58mirrb0jTuiauST01c7JiPa+WNRKtKX7a37of06vVdi9Ol87KU+E14gEuZzadnXffpElrNEXRVDURF7wHmYOQKfgvcDajjUJcwn9gjUha2X6DOurF5QwYuEc6yg+WTexLv976TUf0LtxlzbjXjj16T3n5AnCOmhtDap9oLT/xsTj77n3uQe+6e+elDfFqF8ID5SqzkGRNCP1uaGySJ0TGoOs+VgjZj2CUqMnt+wFhWWFhnraK7TujjoXOVJwH+11Lcfo5bRFfk8ugVwCuQRyCVwhCeSExRUSZJ5NLoFcAre8BMzDgtW1Ab4s9s16HyUCoBOSACUBMAkCgN/NLbu/wV36Nwt5LJdY1HM9wCsgEooroCmLexQizvc38Uuv434LO8M1G4UqAegGFOaewOme6TpEgeidkwJzhHtQ4igTn+RtJAcKDfUzSyuz1KXutqcEircB9+Rhnhf62j8GNbEsMYBseCYWp+SNIk8yjYXvgAooUihdyM+AOgvpgGxQ/CmrAdMA0ihdZrmIzC2cEp9r7uhrzyFZuCYrr3lOUBfyR+6UEet9IwO4NqtE8X7lN/P+oJyWD+ftWuoLsEQ7026Au1+qBFBFKKEZJZ6bJYQAwiE3NvIGMWLD+lWWNLK+h1ywsjP5tZzKHWPOyqOxE4xxH/JDDtQVOe/0MAJtzXNnrb9SfrPCpg0gG+h7lAslGICGNiBEDWPimBJWxwA1AOH0b8A8LI9RvlGyAUtpXwsV9ZC+G2FHmVGgyYcxxzW2bwRlAUTHQo96MlYYZ3g8AfZQDiNc8BAwxdj6A21G/rQpcoEgoU6EaOEZf6zEvhnk+wklyn3D7eOgMr3Uw8isjyqjH1f6p0p/P80UssKOH0llyjz2PgHuW4ZduYqAms05nlBLGVcr/JOsxAVuLomA0D7CXlEgZ0/gbNmL3YL4B7fbC6sjQyWFpXATxcV3BdSOCxBNtEl3XC0Xu4qJHyijqkiOkXY3rA/XSoyXaw2iWL3oy9l3DeOEdmCeBOxkDAwejJ9+yJL0oO/TX3k3/Gb6fY9inaxUTn/iSa+7ek9cHCIvp7X/gbvnHvzhvzrw1p/KrVw3EOxmp7bo332CW+ODNkD+zHHMOb+rxFzIXM88hdfWVgeA4luVeKcwR80qAUCa1+X6vWlYKMI9Lalfz2qPipb6tjbQ7W+0XdKm8/sVBkrhXpxhBfhzRWK4cq7o6Fy9WAhOVSremWbbmYMGUKbJNQb51+vxjoePBoxPAaBtkZBdfSkV/GCkE/Y8lTdui2DRbgCOxvao9g2PXJ9wVnFHwK6GdDSjQJgrIiQ/5cXOSknBMRXubcfehJfQ9IOXMm5pX1vP8Q6kjfibd9dXKH33JeT/27oWQJo1Au9LQj+ZZ+cNG4LwEup3tS5lvc16FbC+7w3Rk4dFrJk8KCWLI9PhcKG88oy8BrRmcccVBiqpjbfkmJfUtel0XWRAJY7cZ098av9RbbR9++ju+unGYmVG3gSuSAjzKnVETCStlUorKvvDCqGkURatDk83KqWhrp6nkIRdERjqEbpnOl4tTWsfmWXle3Goqp1JYE6BoNoXjk3cpT00Hj382hMXRK4QGpODdQt9jjWWhX1iLU2CBGC9TV+BJKMPskZj3cxcwhzCPfzNXIW8FrQnxefd8QUvPPH8R48cU/1XNQbxCP58XbEq+Rx46qE7H73/LZ9ZEHnzoCa2p1v1crJ0ZmS42yqy3sLoCl2GtaId/fUsfKPyClzPv5spSQ4s2Y23GSMYvbzcvVUz1c6/5hLIJZBLIJfAVhLICYu8f+QSyCWQS+ClS8AUUAPuATNRfNlvgsU/YCjgJwASi30s51EkWKwDTgDoEcKGRThALXMzYDLKAcCpWdyjPFiIKQBZ7kfpIm9TkCycEgqwWd5ngTQDuQywl8o2Iev6UslRYIT02aa0kz9ArIU2wmKPsgKko1RTX1OEUGi2AuwMrOf5PHuNLFmzaudA2bYwRyjbAL4AbSiU1IlE3TlnskxvvciDANkDxqFcGVBje1QYwEb+kC4ohShpAEKUy0gF21OC/AcJFspJvofT38gzS1pYmSwvZEQbG6lkJAO/A7z3Q6komecEoVtQICmThdoy7wnkYx4bEERGDlk5kSlyMhlz3sgjSAjuIS8AdSPVkNUex5P/PWSFzPKsAvo0smtQBplL1r6m3hXIxkJkUR8US57FOSMI+OQ8BA19m/EBcEo/oky0C7+hzPIJmHNcCZmTD22PJTLXAs7wO3LkNwsNRZEAbMmT9kWOjCHKYoAgCjmhziBCqCeeAZSNRJ9HjrTZWae52Ah/5wfoqxaKivsYy9zDWKYfodRDhNDvLNQLm5teaxCbul+LwwhS9rTA+h5Zv3mDB/+Yzv25EuMcIA2y7XoA3YwDNgse0ua8ZXlFTMsyu6ZNtEuu55REYKwKl8VWm824FS7GLcl6fLfCxTTbrVAG226tVi40ZG0uXFTBPvygKbA2qpQKSanobzs+rnCD2FxFn+S77R3EuKJ/E/7ue5T4e7MjS1bQJj+XthPjkXcRc37fk6k7cftKXKj8jL73CQuF7PiZuTf8sEDSn+Ldkx9XVgJ98iJNFn4NMHFWifnrX2zzuG/V76R/p0QbM88RJ74nQqSX3b9AJEOsMEhNjYezUZR0CgW3rn1dFsTRTYuHKCauO6quPiIyrywOb16vhjmFo1eZEoWscVc0flb1O/P8dTsmx6qOiIkgCqNKs+VX5SmhOifTAp/lBJV0nG5UklsUPlBD8gpp6wXXiuUlJJJj2PedisiZHiH/5FES9rr9DYZ5r1ytOTtLVNCWrCH4NCMIwOT/vIUw8dpjfWAHZf1vaWKsMvZ5VzLXMqatH1239rnBH8y7HgMRQPq+pT9khUIcOQsn/Wa7Hs0r7NEr1Xdepf4etOvlYyIXipWRdsefaiQC6Z9QeKPxiQOL3yACzJW3xTBkhYB58by2zOvnt6u5WGlplZCI/CAMlB8Uw2Ht76CxJdelai+Q98GKqLURel4/NNva2iJL/m8lStod4kExq+TDoTBVQ1Or3yFPi4f09zG9IVir471KvzZvbPpH30NOifUKBjjoK5Cetj5mzcXaifKw5qJ/cg/leljEy/juOy4cXL0w1D3zzK7bVX/mKfrycdXBOX906shHfvfzPjzz2hN/K8+K+rnnpndJPveLjEGPeEMq8+xagLK05Bn1bNhpjGnXnCklnbKldH8txx9Xc4xuJef8t1wCuQRyCeQSuA4SyAmL6yD0/JG5BHIJvDwlIMVWWM3F2FQas98qZICtxf0H9ISYAFRl5c2cCxCLosRvRhoAJGMhBwgKyETAZM4ZWQDJQd4AEFjBcpAn10BcoESg/LKQt1BPKDAbKd4oI+a1gFbVlnV91QnrLRlWUkZAYgNubYPQD+gcoUVQhLmf+vEcA6cNFKdcRkxkCYpBkoT8KTMH31GMsNYGpKcM1BdFnmsshBOyoP4oTyhR5rkAyGAhoSw/wGkUM5QngDfqSz6Ay1h2mccI1/EsI0q43yy3uD+rLRlIyCdlQMmzNrXruN/qmpW9WZGZnGgnCwMB0GDkAUoqgLfVEeAREBxF0spDHkbEUDdkthEhhXK3buWX1ot6o6jSB7nHQmLVnaTbdjwVqX2Ufsm9yNc8O7hvu8M8jLjWrEfNko82QhFG0QXYt/5sYTDoA3gqQIZBICAbZAIRwcGYoEy0F9fQD/thD5SQDQo5eVk4NJ4LqWDhqMiLcWhWgxbmirzIB0IJotA8KmhbDuofxc99WFtZPjylwNa7hWggF/Ilf/Jj/CFP2gGvFfoY6WYmK1Lx9OVD2yKvH1QCGKXtBg+A7l9QAvCgLaydNrj0qpxaRzyEYta0Oe+4Qj1NKn79qObvOYG1NQGv4iKSlpBNxfv2gi5Ap0LeiLmQkWes2B9xRfEuPOEwDVmjNyMv7nieX4K00OXMLVcL5NxIIIwX5jaIMiPJmSf4/s+VAIN2cvyWLmIetxAyzD2MT+ZDxhpjMjrw1p+MHzvxb8jfDuanB7Rvx/v12QectH/Hts/T9VxjbfFZ8+RO8tj2ITfXBciWuYn5hDntl5QeUcKL699vU9Wf0O9/ozSrBPn/e0oLIi1aIi3MY7GfhYiHVqHgy5MoaqlR5H3gTKqn+26UHBFxp70fHBEZbujEXltAf6fbCc/1enFdhJ7IjosI7msufQiLerNbazbj8aFqcVTjW14gblnh2laSTugLvx2RF5WrjWtENcYj8qbwAm02rvOLqmtXeGhP7hdlDd6ahJ31rLwidZG8jaQgP/JnXQOw+2VKb1ICCIYg/GalB7d4KO8pEmHCANdpV/Y8YZ8KwGYLXcj6pe/1ckUqcPNmgoxYI3NcNHnhabF6wYtaK9rDJXGG5CFQ83ynKaLiqAiGO+VhMaHPRW3ssrdQDu9VCKTi0pnRdmulXF05P6wlwotkBZkD3gvMX1YopEAkB5tUt7ygfKhQjOREkDh+ELU6qyWRFf3ncfAOxZhjp4fpBrreddr10meU35jCSx0uD3c+KOKCvkb/YN3Iu5p1FX2G76ypzRCJ9wDvZtZV5Mn6yAwweMehc3AN8z/fTytMlnv4NSfw7CguHB9/TAROXfXrG5yIxHlzY6F6/5Pvu5t3CjXD2Ih3Fs9/h5LpO+aRa2vrPRKMAtNppxy5QKF3pQfvKtrqWhsI7LQd8utyCeQSyCWQS+AqSCAnLK6CUPMscwnkErg5JTBIVlBLndN6WprG2mGEhc2tfateJaxW8UoAlP8aJVyiuQZwGJATBQEAlJU510AUsMgH5AWcZWHPwWL/NiWs6FAcAK0gKgCTUEZY+KNYAO7zmwGv6e39D7O+zwCL0t3CC5Gz+thZZ+hufkeJodyAJIBjX5uWifwAaFEaKB9KH4DxYP78zW8GAACAWYgiIwSoK9cApiADlHADus1VnTqhMFEOnoPMzBOBZ5AHv5OMuLCwCChhyNQA1Rl9N+IIpZ/wGlnrLkCcjcIoWV0MeLC6AMwbMMCn3TsoCwsxxXkjPQDMaVc8Kai3kQe0JSQEf5M/QDiABkokoD33G9FBvii1nLNncJ+FNTKPCvLhHH8jOwAw2pF7kDPk2MNO+9htTrRacOqfGLR+t/yy9drsu8kDudN29EHkQvtkPWV4PtcYcMZ3xgIEgI0L7iU/+jOKM8qqWZMzfhgTyIeEbCgnbQ24x++cp76MFeqMEk3/Mus8rsc7AMCHMgK2Mw4ZY4w/+kqY1Ofc6C9+dipZvXC7zCbph8iMcuAtQJ1oR+5jzOGtQr+7FcgKVbN/0OdIyPn7lL5NaUaJuQhZ2p4q/0rfAVCRHXNhP666ZXKVP4089TVXaxN1J9JnS4SD+mgcKIaM9qrwS9pEuK3wTgvEuldEf5FTSaAIMSVfjhnqIb1mq1eTrXZVFunEnelp7u+022FbIaWiWsWqefk12cEeFfRTI8yoE3/Tr1+v9I+UCHdm74qtCsIc80dKf6LEOIDEhKwzz0DOsYF2di6gfZmv8PzjgBj5oNJnhRvKPlgkhb0bs4SvtQeX2nvA1bXWlzYs+y1KaCAT5kDahrmG+YdQdLwzeS+zntjswKqaBBjO3AUw/rz6GXMXoeqiNJRTT54Wofo/G3DLe8jtFVz/Me330FR4GtmKu/MscbTJRUv/zYnIOysPjKa2eumycfcWz7/qPy3X267COCXNdlgOAq+iceitNDtj6myLfuDOiVgpi3Bh6daW90Up0Z4bGuvyqtBE5Lsr2oC7KQ8rTy8GVcdlPF2xDcRTsoL3rlm1Q1QQ+vCrldhvZEYJ0mK7Aw+1dyvxDmR+pe0hC9+rxFjGsKM5MF63y/OW/v3jj/xW8rlf/FbzlGVcsfZYPzoNd/LkE5WzI7udA5XR7ll5Q4i0iCdcP1mS98RUe7U0pbBLkBHJ8pmR4PzzU4QZ+zvtQ/EGbJpexNj7WT4nz4zbk7jcFL09rOvKDQUq0/4OTkGRBOW5odBS3uA9rIdY12eJC9Y3ts7MhlJaLzfPFTlyQGGhmlHkjYzvXx5VuQkrx7qR/sOczVzMWhMdgvwxtqCfsmbi/cI7hYPv3Mc7hXUVaye+c3/fa5V9nuQhclz7WdS0p8e+s89On5FcXinS5o50U23Wr1lPafoq677smvBiAkI7cmsPi9iVC5SIRV26vkygzqz1WJtRl2u1fkjFkX/kEsglkEsgl8D1kEBOWFwPqefPzCWQS+BmlIBZQ7L4ZlEOsYBFOUADlnEs9gGGfkcJBQGrcCyOsbhDUeA+FFuuM+WJfAyQZnGOdwVKy2NKAO4oD4CkAElcayCtWYwBdDcJeQCxkgqdcwCJzP9rBEHj8Zaz/3uHnNEHZvQ31k+AiVyDQkeZAWFR6sxzxOKjozhwZEMeZcF7U0RQsng+11FO2y+C57P5H+XmuSRkA9AMkI+yhJJiipNZYPFpYBpltLqgxPCd8nEfcp9N86cOKDsoSsiOZwAEUZasFSSKIm3A7zzfFEQzm+PvLJDHvVa/LBCn0+veJnw3wI5ryJ9yAqxbOAiUOBRFymyeJZQPjwP6CPdxjXmWWJnJK+utQzm5z2Ji82wO+xv5Ul6uof9QT+WZlJ3eStUpTHOdkRxGQOzUIp7y0cb0FfoyJBP1o4/yPNqEccHv9GPOA+JAkJlVt3kdIQOrK3kA1FFX2g5ZQJzR/7jOyDHa0jyE9LXfX3ke1oQ8GzmhQAPOcg/nKTN9w6wK+ZvxU1OA6V78lz9fdVbOHhLkRR81EN720SB/gFzyoWxsrD1I+HD6VjiQyf9I2wUQDiA1CwJxjrFOO9LHGOvXMjxUnzxVKKi6rLD39kOYKfYEVuKhlxSqZVfG1rH2342KOlcoBn5crPgJG6dGUeiWy4WWANyeAF2/XPIbIi5aIi7mFQ4qGh8xR7Or0sw2zg2sYc4wwpixDPj5vTt88jt1HfMLZDN9ln5POzAW6beQFJuBQPTvn1f6r+mzeH8BdtH/NzxSssLmTeZSxp+F/jMkir7AmOfolyFNO6zSzXPZNnu4JOkeF8zFEKp4x/yl0o8rsX/Mj20jCUJEzSphlc+9f516W/QJh3RPi648hupR7HRE2skLwTkjl6JawfdCKD55Iulf0tS4aWsc9TROrnsc+aamaBV/tdnpnZE31ILIQ1l2J+Je2FybPTf03lFIKBW8v3bRuO0JB/VFYuxTHcf1Vu4V/eACkXSCJKZ/vqT9OFKSwjxoAXUxOrkj0/eZF/Gc3OmBV81/V2LeNM9OiCf6AO9R2i8HbncqzYuvY95h/no0baP1X8VdtRdO7HnFcx8pjtbGu8Gu2+fG5U1Rqoy2TskrQuGgCtWFU2Ox9mTwwnahJZJgTqGO7i5Uu7JrcJ2oG8g7YJ2EGNJ3bYjtEaps7Yh9py1PDHld9D0wBgiO/hVKg56t27ux9TN3h/FVzzcJAAAgAElEQVT2iI9NfHp6ZiGamplnvcM8b+GdWIuhe7BGo0S8B8yDgnHCu5znQ3Sw9iRhVILeYYQ46yXWZ2NeEDe1Gbn2gonvV9rVWKiVFk+PBiIuhlWvGV3Dmoy1IPLGa49nURbzlO6X2g7GbdhuFiI5/SbysMgcs/qO0UNOVlwksfyPXAK5BHIJ3NwSyAmLm7t989rlEsglcG0kYFaQKPAs7gGSADhRCLBmRAHgPJZGKAJYYxtIhCLA38zHKCgooljT9eNn6ACwIs4uIDyKMIorllcAThwfUbL4/jwPyyn+5pkbWf0bIGQgu9SIVuCsfKzrlPYsOpXbbQ8BlGHAfaywsK5CSf56JepImQEb+R0w2ay9zPvAQiwZKMUzAZZRUAAFDMTid86hPFE/FBnyNVKFT+4lf67lPj7N6p+/eT73AaihGFF+5MM93D+jhNcKVvqEXELhogzUn4P8sfinLoBp/E1bUI6spZmREaZyGphuYDl5Za2J7TrKaMA/11g4I/oI12MhCfBuZBCgLuVByQQQpG72DJ5p300W5sVD3rSN1ctCM1kbWEgA2o58uBbCgL73WqdyV81Z/bT2MqkYoEh+Rs7sBITPAqu2P4R5TvAcNE8IBeszKMmQCRAPKL88A6WacgGGQi6h3FIG5ENbcC8Hv5E3sqR/8mzqidzoDxzIDxmQZpQYV/QbymAhVr5A3z9fif6CpwVlAdA9KbPH2eTk4/uTheMVpzzcdatjn1YA6lgBoigH5aGfQSAyzrBW3omM0qK9PD+2AVSp/7IAuw/rk7HzjQO1ZCzSn/8vJcDVP1Oizeh/10J2PEPRyd1VdZaFMEoORlFvQqFjhsRbFNvdqMX+FDKzbouI8AVsrrKPhay2L3S6SU/EhCLLOAr/5K7IEntVoXBWyqWgNzZcpl/Hsv6/0qChEZzMY8xZEHXID/DzjUrm6bCTzvTTaZsAzDHWGHvMl5Q92knfpX4iIB4eeNjn6W+svfltPSxUSlS49UYnUNgt5tqaZFaV7AJZ5g8LQI40lFY1mxe1aXlTo3dVQLPtr5P1crvSMt2JrF4O1xjpjeyZMzFY4N32I0oQWoMH7xDm9Zk00Z8gnvC2IBQlYaL6QL08LfoEMKGV9Ek4qIraTO8YV84IsYHjmgf773Pz0LiuMlM/64qhONdqdV/Qp4a4N63hekT9yxeJMYr7hApf1oAqQFiqsLwzJxTap1Mu+rPsz9HthtTVxtyG9dnCA8refeQLqMy7nYN3EQYHkPK8q77nEgTFePgD2kgJrwzWe7T1I0r81p93lPIxcglCHbiU9QAGDHirsBZgPYLbtOP5hS+Neu7U8rmawoYVbisNdaKxvctFbRjdDQrhvPZk2HP603saIhyKIhxYY9ynPR3iiQNLujd2FI7plEIz+VEv8LWZ9md0jcIP9tci6654OjcvUyIz+hmsha2paWfGGusZ3pXbkl198kObyssLZOnJ99/1zL1f+uzfje1Z2Vuo9L5C1Mi0QqZ9RvZLn0zry1qKtTFGI9aneDeQeN+YZyvlYa1DGSgzBEQ/dKfyerW8Re4d3VMfrY62LzQWq4/UL9TK8io5pH05mDMYH+THu4f+jC7E+4t3w+ABISrSR95Q/YrYknr9MuTAGtHWfBtkkZ/KJZBLIJdALoGbSQI5YXEztWZel1wCuQSutwRYYZvFv4GvgLeQDCzSAaP5ROFEOWLhD2CNpSTAK8AueaD0YpkHIMpCH6AWMNXAaBQJlAyUBkILoERwHXlzABgyvw96A/AbC32UJp4LWSAzsChwqnfo2jVVJ82PZwJsmfX+t+g7ygvKAuXnd/Iyi3jyNkDdwHwULZ6FIm8gOefM2t3CMJklGdcBRBuZAjg8qLXwvKySTr6AEOQBgGNW9VyHMkbIKUA+QBtzgc/mybO4x/LkPtqQtjHwbN0uLq0L5abufdBGCWDCNCsjGEwZMzAD+SBbnoXcOU97UybOmwUy+WXLY/lY2yAjCwHFd+4zUoJnUCYUQ84hGyMoyNf2hqBe5AGwQvscd5qfqWkfi91O5xx50sZG5FCWz9IaedDAYSSVESr0RyPN+G02LQt5049QPJEbbQSYw9+AB9zHPiOEqqJvQ/hZaDDy4X4LN0U+1Jf60CexvmOMUWfKbf2KepuXB/dTLsYlv9M/ICkYQ+SBPOrRh34ldsf2dURWTAh9mEo6+ilJLISELum3G/cRisMsxDl/qx/IFjCEEEX/Qekr0zYysgn5vF0J0P0nlSBCmR8ZN1cLfFsfH41Wt6JY9wpl4SxBTqTeZwoP5ZZ8L+jIFrspAEbkStIolYOKAE+n0wu1qW8cC9w8IaLjjK5dDIIA8oJ2h6y40oQL4xZ5MU8SThALeuZ2+i6AVZasYAxw7eB6njmA9wdzI4QtYYQgjSgzYwyi4lLlDTAO6PorNKIOvDvelbZd/4SRFZJzQfsiDGPFLqZnMmSfgDBe7PSSaYFmwwK/V7RXSFveKrrLPQOYBwmkP8zjoj+PXgUiKC36TfFh/Y4xB+hq75P/Td+/NFPDwX1lXq/fIGq/XwljiCE25O6340MP4GXTFXFhnnodeSdo/l9fG5Bt/12UhpO6roLcOz0ci7Bwp8aq0eJK+4z2oXFFJJZEuLjah2ZK/c+X6xR1mNMQntB4rgiQZhPudqkQzIusaOlaeaB6y3ESGmm2kzrZO5EOzPuc9QJyNmIIsh2vMsYuxhg7Pf5cF84qMX5ZF+IBwDuSscE8yXjOvu93mm9+3YAEFBYqVlgo5Ms6BG+CNcJCh7YmEmvXvS1sO21tKj2uvScWBMS/UCz32hJ+c/Hk2C4RAnvlTaFIaQop5mt3+unV7u475lYE3kcKibSqTacb2tshaS2Xn1s+N3JUJMIpjaJDIipY39OmjLntDuZ1M2basSufnlFSL3EVomrPc3995Nk9d58Px/Ysf2Z4epVNxG/Tiq6lvTPkcbT+CqAs9C3WU6yF0CEoJ3oC6zFbYzHX0NftfU4/ZdwUlF/gDcXalcNpiKgoaGPxp9jPQ2VhbQcxiiHKlygxdhgng+tK5v6GbliNwt4uppx+eK0XJcSY4rkvGlttJ73891wCuQRyCeQSeNlLICcsXvZNmFcgl0AugRtIArYABwwG+ETJxOIR0AkAgMW9AamATyigALLEz3+V0pH0ehblKAucMzAepYC1OwqEWddTdUALiAWUCAP9AC5QPACmBsE0szRHYQIMp8yh03gydPxh2yvBPCIAfikj5AiAGUAkdTGA3rwDqKdZimVJDGTA3zyTeyh3P+wCBe8/92JPB86ZDDcC0yiXKSt2HQoU5SZfA2wA+lCSUECRKWQPpAX3IE8LncV15sEBkGcEC882kgnFyuTN/cjYrLusLn3r7fS6wc9BSzALAYVsbF8KFDVAD5RESBcURCMtzEOD9zV5mQcIsjJywMJdAfxTXvoUdafd7PlWB55PP0T2KOmHlVpO7b5xbbweOMt/S93t2cga+dJ+OzkoD/3awm1ZWC0LY4LCaXtz0GdoF+pNWSk3wA7yQ66QAfQ/2op2hWCg7ZAZ5cJLgvP8DfHC/WyszT0c1IH2JC/KhReFeV3w26wScofkMAIE2U85rZWSd9vnB04Ulr273jAXPftw01k5NyEEAznjQWAeUcixa5a323ggpMW6uT9SEDyUTABC2SMBwmIjS0qAC/rgjynRxmd1D3LdFES/AvLtz2siKZbKxeAZ7Ukx2u51QxEXSblY2F0sCtuMkwsC2HWdO0Rs/MiPhXMm/T4t/OS8PC7OKizUikJHyfI2CkdqpUsF/bfqAIxV+jZzA1bZ9FMsX79JaWaTG+n/2QMCiPcJc8EfK0Fa8L3/LrgMkiKbN2Pzvyv9G6Xblf5J2n6Q89lD8bUSRRJS+QXmCUQuy4NlXC07EiXxblXyNmILeYkgwdDtaK+Qp0RuLMiqdlEI1Tn93tDfZj1+JeW7lexfzr/RLryvIKaQG1bMP6TEu/q1m1SMPvYTSrNKzJ18Mp+2NQ7bpbc+YOsGyAv3RiAnNqoHhNaffeJUUqsW2ZfigvoaG4eX5SJ1SFvNaJ8Np+f5bk2kxMmoJfcL16nKc4rNw+VQFa/KA2hFdEVBnSzWPLAT0tTep8iPdRpjlDUe7zD25plRYt8QvFHxZNnJwTuItRQeTJAUzAG8p3k/8s6jbfsko1I+HnYi0Z1fY8YGvPvXD8UOxNOipl5Si/WWaq9UJvobY2Ns4Tqz8owoCIhf95bgRhHd9epYa1bkRVshowrTR+aX/GJ0TqB9oj0l5hQ26ndXF6qVlXPDUwoRBfHLmnSnBwYSdnxMX/DWHgwZNZjXV6uMX9Bcqjx/7LEDTy3tGTmu/SYWR6br90Shf1b7ZzxbHW19THtPfLQ63vzCtM+xliJf1jYYkNAHWVfR1+mnX5M+hPmBNZwZfrBGXJQMSoVSrzV5aPH06ny1KTmMSVaMDQhUDK1YxzLOWI8OHvJWSZyw2z7fazdvG9hwm2stXGeHPUh2Krj8ulwCuQRyCeQSeHlLICcsXt7tl5c+l0AugRtAAunG2yygUX5YVLOQBzjlHGAAoCwKKMonoBwgMdcC4AISoAgBTBlYZZb7eBigFPE3lmDM2YR+QHFA2eE8YBT5c52RF5yzPAYBc7Oy5x7A6DUPiLDecyqH8dj4gNKDStQDIJd8AJLJE2tBQF9AMAgKFHKzVtfX/vN5noHsppQYMcI15t3AJ7/zDLO2Ms+FLMmStcLKKjkGjpvckS0KEeUi7A+fKF2ANihhLyih+BtxQf2tLJQL2RsBwXfaByUWYM6IAa6zMpjCZPXgN2TEYXtApH+uf9i9WEUbsE65aX/Khixoc57LOfOSsfJkLcsoH39zGLFkpAf9intpT8pi7WKEDcovCiggCWTCpBMtB45Xip2lh7mWRFnoGwAlgxa6g/ViV9OY3efTa827wkg2yALyox3MA4X24TlY3llsZn6zfgnoZuQH9aQfGqiAjLiX+tHGXEedeC59ExCX+vOd6+gDECDcD/EGkQPISnnMiwbyivouO1Gv4u6910tOfUrtJGt7z+ecEU3mBWXkkW7Jjw0kQFsQ2u5HlfC02Oj4Mp1kPgNkBxgxLwCutfnrkoAJAaubNUZs4W66vbhdb3Y7vu+9IJDSq5YLhIEa7oVxWQ/TuErKOj3SbveK8gKYCwr+04rrHwuMWSl4zslWp3deltrL9U4vesur9g0Swpt2hi1CytAHjchmDPA3cy2kBeNmZoc97H26Dgtt3jHIFeKiH+KH+68A4UM2zGGMOzu+WV/+s5IBf26r3SuIsChj5S7ypyzQbJdkd4/+3t03mXUSrGeZLRqgxspSYbnck/Je0RydNBUQRA4ZSSQwOWYj7tzLYk3U24VkU/+irWkfPGF+QQmgEU9NwNGNDsBGxijz+3cr/aESBP8p5WVzdyyvi+SH/pdtn7/JI67+6a967f7oQ0/N9UaGSl11uJFOp1cUsdhqtHrharPXkHfUAfmIaPy6cxrfvmJGaUMv11N/WwqbvWV1SXn4JMuVcqGjPTGy641+4dN9Kfhq6zPWKbwvIIMAjvmbdzDpX6fy3GnF/0oXQhzxXN595oHIe5n2JG/mwOQKjd+dlutWuQ7ZsoZgf4a1ox+SKNIrv619KELWt1VWNknksaZg7XERdsLl8lRYETnRCQrRtEIvDRWr3bp6WUv7XbDWvzC2b7kmbwxX3hYrT33wzkB7PLyfzbf1m4H4PJn1o5FVm+EzvB8IxbeTg3GtvVzcqsiSoaVTY6dUpl2LJ8ZYAxfj2H2mVO0uH3r1qXsLlW45KEVt/U4ZWCMxx7OO5h1k6zrWwlYu5hnTJVg38xtrrOMKjVW9/e+9cOGZh29/pD43zPqTecbWcOYx8lnjjAppLJaCYjn2C4XZsNOcWVtS9g/Wx6wjWTvzTsyPXAK5BHIJ5BK4RSSQExa3SEPn1cwlkEvgqkuAlTXKBGSFEQF8QjSgIACaooCikB5VAtADFEA5+ColSAGABoA7yAus3wGaUGjIA4WKvwFjbZ8DFvEoAygPfEcJYFFvlnicHyQs7G8UCBSONYB6VdhW+yRgLEo3IDJgh4FTZvVuzwcc7m/orQTImw1RlLXo10/9g+cYEGeKCp8obGZJy7PMi8BIgL6intbB8rJncR7lyjQazqNMAvyRJ7IFFOcaFC+UPAOZuceARiMRKJ+FlyKvdyrRbiicWUs65GZ1oUzkw33kAwmQlZX9bkQD5ARy64cdUqK9aX9IIPLhPKAj7WuhswAxjDDJgrdGYnCO7yhxtD39jz6CzA3ssH5A2Sgj19L/UEYBNgkFNec0n9rtaL9DCp3eb+XeULlMr8t+cK+RNvRzDmRDO5NoB7MKpBwQBxATyJN2o98BAtGOkCnmeWLWrJSHOpIX+fAJ6cB1pshiVQ6YRPgBiBC+A+DOpNfSL3gm5AX38UlifNacsHM+adcL8aO/5caffq96+FJR+1lEIi3OysMiC07vGKhWvrfcgSW/gD48Uv6rEvtV/LbSRqFRvlfnGRN4F/2tEh4sEE3MRcyTlxKmZTs59+cTeUdEAtVXpidqz4S9aEihnbqyuh5V5Js9pcDv6aK5ldWOJzJD+/E6c77nO67vdAWgPyveYkHW2Q3d3xXJ8VL6gI1J8mCMM+cznwIw099/RIn+vd3BHAIhxDigHz+cyoyxyBi8JMJnu4elef60Pt+eXosl/68rAfo5z8xecCAqJKuyvFh2VcrB3UEhmBFJNNRo9kbDKJyQ90RFGyN310KUu5HA5bsl9xGBU7FuqhQL3qK8X54Q6REJRLb3ww6KdstfkiXvIf8gZSEDscj+t0q8ywYPI6N/VT8YAM+7j3sYl/QpxiBz5ZXuS1eswVabcuEZqXRFdK2qH51pd3pj7U5Yara0c6/epepTceC7UU/9sBgk7UAbb/d6yTld+5lSuXBSLhaLXc0LuvaiMa05zIBZ3j0W7982u+adgRcs8xWh2t5yCRWCqOAdZ7LlPczz+Zuxm4cZvARhvoRLaW/mXfo23i1fTl4QFmG3o+VAsxoUSvKUKDFObO3Ceog5mjHRX/sJpMejIhFRMS7ygn7CWoe1POvyp0UEjLh+8mp5YDzxOV/+1Oy556Z+4/lHZ94jIuGL9fvXpvnhIcXeT5thM8yxPHdbAxJdY+Fb0R9Ya5a1l8Z30a9EYAyVR9oHRycbDW2WPSaPkOmVueFWZbj94cpoe0Fl5b1NH6cs9HFbI6NrICs7TPdgrUpivvlTkQ69oKhdxlvF50SKzKTlZR1ma8vN1pOifhB9OBz1ujNxqGXhi4QFskYPop2QTz4+Mg2Rf80lkEsgl8DNLIGcsLiZWzevWy6BXALXTAKpl8Ua+L+2mAZYNUs8lBes3vmbUDYoAwBUKCtYNGKhxIKfePooroCtpgyRD6CDrE/75ARgroXzoX6AECgn5IlCxX0XkRSULSMIrsMzAsUYQHdtT4DWC1WnfZy/uZYyQFgYcYCCRDIyBqAZcBFAg2dRXwCzQXKBx1pZeN9kwQAjI7jXwHV7J9k9pthky58lGFCebBM+5AIwDciHTKzslCEbusmIAT6pu4U/Qv6AElxLHuyfgJyQtXk6kJf9zf2Uz0B9KyP32rPNC8LkAjBJuCYjimh72oNnmjKMaz4hJniOhdIZlKs9y+SFHOhf5AV4MqMEqUSeg7JEfuQLUQJBgHJ9wQnGpZh6JSdaNRKKa2hvymokBPXf9Ei9LJCpWQlaCDRC/tDfzZMCsoLnUxb6LvXgNwgmnmnkBjIGyEbhps9Rb66HzKOcWLdSNoBtLALJ48H0GuQHEUI/x/KP78jD4ilzjnHFdSTCH5xKWivz8Yd/3Ysff9eIjHBlA76QJCvnx5yoSz70r5cCUuv2W+dgM2cBfgA2tNG3Kf280hs2kAD9gcS4BbwBPKUffUgJoha5E6rGCLgNhbidBXK6qXA/brg22cULoK5o48+JnDhUqxSrAtpL4qTKhaJ/3g/c80XFux+W1bYIjlAm29q3wruw2ggbAOlK8bPH5i8XwKW/M+7o//R35q4vUoJE/KX0t606CtcBJP+cEu8FQvUZacn4uJp9lDr/spIRFgBiWNcCkCcCjt1KKfC0iTabbE8qfNaEom4VO92wBGinkD2jTi9KdH5Y8h5q9xTl3fU6YTmYEAF0WzmJpp3EOyZZn+5P0J2wLi+LzlXYJ2Qr+d4MvzFWIP0Ye4xB5tQ3pv3MwjcO1vP70hN4Pv1/SrzjIdB5bwGuZ8HKG0pGeFkoNFRX+1nMy3OqKWKCcTopokJjzV0eGylX5X0RLC21fIUla2n/ipFSwV1QDLiz8qxacQM/XK63Qwt9lRIV5vnEu4d3kHnnMX6R4TcovSkVBCT4To5fTNuDuY6weYwb1lvzzJc7ySC/5spJIN3HgrZl7c1cjIveuMLTsfGzE7ZbTlIbZV2R9e5lPc/7iXPMh22FQdJCwZkTQN/z1wgL+g55sa6AiGDtMawlxReVap3XHrz/9EMiOZ5/+oN3TotIYK3FOhRDla36AOso5v6dHLxP8bBjHcjaaH0tqjK2y7VOPDy1eme3WQi0H4dXGW31hiabC3uHzv6t7yeEvaJfskeR1Zu1HGsx1k3UGeKEfFl3mtc4dX6l6vPxuaOTq42lCjoB5WANyRyylWcEv4XirBudZv1Qr7Uq75aLOAnmsFkl9Kf+Ozw/cgnkEsglkEvg1pBATljcGu2c1zKXQC6BayMBA5ZROlAsAIvNu8AW633FRQlPBhRgFuGQEtwLqIuFMWE9UHYgBLCgRaFikU4eKAwoRABFWDQBUGO9hLIAoABgZWAteQ4qQCgQgBcoP1yLoiTf9+aKbI8XpCW0ZS8GYM59BpibFRrXcj/lhTxB+X6zEgAHz+e51DlLmGRBPSMgKCdgCvVH8bEwQcgle5hnAeey5IURC2a9DwiNQoO1I/nZnhY8G+Uye3AP5UQRM7KCvK2u3I9ihmLEcwxYz+6JQH5GVPCd/MzqjbwgP7JhsLjG6vJKfQdEMu8S7jNgib5BefkdmQBkGtlicszKlzwNxIVcoS/QpiiXg94R1jf5JG8U6TU5xtFpJ1ypO50+RkgyTxP6CH/T5js9rO/TR1Dq6dPIDnKAurJhMM9FyaVf04ex5sWbBWCAtqSP85224G80V9rUvIdQhDlHOZE1bcSzaDfalfsZN1jkce0aKbcWZ5zfyJfnIWfAXoAK+k8zefzdcfSn/8FxR/e2ICyS5oJInC7PRqYbKsrbAeW675Y9UtLC+tu/lCBeowTgvdlB2+B1wUF/oZ8w35EH7Ul7c2wKWij000Z5Z606I0Vz8s/MrTgCNy/IE6AoIJ1xpDZ3FULDWamWCr4+A4GelOeCQM65+mq4KgNQQsd0p6u15DveeNeOCIs0pEz2+fTtr+s/z3EeVfoSpV/ZYSfBo4HQPcy/9GnGB2Oew8bvDrO67Msg7/qhUtIcIN4fk9xjbWiu3VZ9tRsbNTuuCAc22N4rsPh2BeWZFBFREpjckfeKvDAK7DfgajsBJwj8fWqLcrMdPt9shXGxGIx7XtysVgqMvfy4PAnQH8wT8jf1nbUFczlE779QYg7c7HibfmAvBvoo8/dJ9WO8dzYlxK73PMgG3Cof87822Y7PsC9KtVIcUV+bkOfFWKcdlrzA85qN7opMOObpW93I0X40cbvbi8KvffKHPUJf6eCdy/uUccq7Cqt73ssPKvEOYT4aPCDtNjt+Rz/gYcY6icmJMfunSliy816h3DuaS7Z4Rv7T5UuAuR/iF8Jg3astiXpOr9OUl0XLC0oMgYsO2rBv/OEH8bnJw4ve2J4VLZ0Tw1V4PzFHsoZ7UMn2hiCjJS0tVnfdNl849tjBpeZiRfuvuPzOtXZkQ36Sl60vzdPgkM59VqEGysj8zPuS6+jHHK56WmHl/PBSrxuMamPssF0vezpbUMirV41M144PTa12VQ/usXcsBiHI6NVKv6f0LqXvUGJ9yBzC+4DEBtv7lN+ZE0/s68h7BN0ALxNIDdZXjKGNjJq4ta8HyLviQrexPKxNt9NL12tEXcxzOB8rAw2d/5lLIJdALoGbWQI5YXEzt25et1wCuQSuhwSywDBKAkoNgDSfALTMuwbEAuICKADKAQagKAOuAsytEQlrgAH3ZYFjnmHWf3YNiolZQPJ7NmXlANj1g0pmNUbePEuKkG6JV+ccbxSljfJCqgCMcVBuysonihX5v0cJANLA8ew7BcDKFHGzRKN8lPMDSgDVgCefr4QyhkwA7M2iy+7h2XbOZEudyZ/nYalIOQG9UZqsbFlCwRQcU9r6oEb6TCsn9yIHyki58H7gOWaZz6eFczIiyFzT+eQc+Rr5YX9b+Y044hkkCANkC1hOu88qfYGSWcbymxE55G8Kq8nAiAvkRh6U1WJgW//IkhbZ+1B6n1ACfJEpW3PU6Z5vOxfebaGb6BNGJCEX+syOjtTLgjqYdwTfIS3Ij34O4IXsjViDNKAuyA4l3UJ6UQbKySfKuZE6kBMmf6zvLTQDCi3XQ1qQP8+CtCBvFGUUZgAiZMknbcnzsIy1EFmx90Xf6bp//Rtu8swHyQOZ0x9aAuO2sg7UJfmxmQRS0sJCoNGnf00JQNTG42a3fr9+IP07JcY3oA7gCXMXn8yNNjfgzcGRaMPgzwI0MiSGjfeuNtUWTq4IFFEyL9ByebhWOilC4mC54FeVgVcXsClcvauwRgsC3CNhnQ2B6styuejOLzU3tITNkBNWLvoz49LISJ7PuPtuJcY7x04sq6n//6P0biXGKWOe+tOP+/Ps1bbQlpeDI28Hysszscb/9bT81MeTdXr0joePxvKsWBvPkp32CajJGWWv9t5OtJ9FV/sHKCRJ3Kg3Fa9HLizaC6RIwC026RZxUelF0aTuHy+Xg6FC4I0IeGae8PO9LFJJb/GxBWFA/1hS38SjDpCR9sGThzYk5Kz3Vf0AACAASURBVAtzJfPq4AGxgbcTx+8qMYdC5DPHMq/fUAd7naifxGfm6s7uyaHlTi/0ul0ZYOg9qr0pzinGW2GkWFDMsWBF3j093/cVJiqpv+LoO7qHZt/p71v5FF4TrB949xLeyUJOvjWV06XU9zt1MXMUnlOMF/oxXivIkO/Mgxa681Lyza+9whJIvSzoJ6xJ8XohvJcWGZqtFBOQjRXYS0Frm+yTWZMI2I/nxg8sndt124VCaagTyosMQyIOI6PwQgDUZ33CO5CxQx97tbwy9t75RUc//Kn33PuHUdfnfYg3BAf9hfWGGd7w3rODtaIZubD23ewdyjqHeRmyADLNjIjE3blB2PVr9bmhqggLR54ex1cv1BLtrzG85+5zh1VN1r9GmFBmyss7jD7L/AGBx4uAfgyJQFmXle+pdr3kX5idOKyNvs9HPR9vSZ7L/LIduYKMm4rZdiHstF+ZCQVl9Wa+gSQyg4WMSPKvuQRyCeQSyCVwM0sgJyxu5tbN65ZLIJfA9ZKAgcMABSzWAZYAVvm0PQlQRlAGLEwNwDDKB7+b9wOgF4ApyhSKCtdYuCmLG8vftojneQZkb2a1Rz78Rr7kz7Moo/LR1rLdc3c5wSjgMM/Eot3c25ElQJk9D8vAf6KEssK57HO51g4D7uxv6oD1IuAb76CfUsLa+OuVAE3MKgylKUv+8N2s6i1PrrGwTgAv/I2MUW7MqozvGyl1WQIA5QtQmzrQTsgGkB0FiTaydrOQRgawUyfyNstO/uY75TRvEzZIx1LV/NuRv3kMQLSQpxEhyBKwxKzJUBDJfyuvFZ5n4ZsASADpURRRZrMatpUROVI2wBnKETnds4cdtxc7XpHn8zvtgAxIlj9129GRkhZcy3OMnECuHPQb2p1nUD6uob6cR7k2Ig3F3ggX5INnBCSP9Qtkw738bW1NWelf/GYKNpaT9GHyhgjkN9qTZH2K/mTtGBf/1QfZf6Ef+1wputpA8JpYbu4j3dOCsURItLcrYWn8LWkb0O8ACDc7fkI//IES/RzyjPZifBLywkK4MYdxvqu2Iz+bl9byfOgB52cfXPe8cAHXITEEXNaVVgTSBNqXIiiXgkaj3RvRRtyRgHM8BTrVssxQFTum4HsLvecebfury8m3vPXbIUhsfBkYRB+ir9HXbbxjVc04Z059vRJ9fUbJyApKNzhHZuXAHMS91JvxzdyJHOnP9NEtw2RlM7qC3xk3f5KW6Zv0+QNKfyGw+M+1h4UIoNgXGVQVuTOqvSo8IWReIXAlw0Q/xZFIirbirYzpc1ghewjNtaAMxR65k2wWIov4M9r0XN4sbkE3rLa74Xl5wdxwAPkVlOc1yUpjsJeGaCP8zawScyP7ZwHQbkRYZMv1rfqDEEi/r/SvlZif6fdr75AbxEMg3aA9grigfBrTDYUp6xXV2eRF5baWFtxqkETdTqNXd8Z7n/Po2937z/zJWCFq8b64RwlwmfUAMoGwAXDe6cE7BRIIT0fmJd5lzFGE0+L9BQHCO/WiWDc7zTy/7qpKgPcFaycMh+5WGtIc5cS9rkN4omJlyHEDWzKulyMQYdHxg+iMF8SfllcCczPzP2s43gWsSW39Q59i7cGY4bOjb/XxfUuFofHm3PK5YYgsIyx4H5jBUtbrggdbyFPeAbZu3ej9wRxNn6Y8Nkbpk31PaJELs1r9vDLsFORBUlDIs6RRKIelVr18Z228dV4kxsNK9+ta+r95H9O/GSO8a9FbeJfxrmMtuaz8FN0v6a3O1yoiKzBksvcjcwtjgHWf5UVdsod47fCZxuI5Pw43tA15vy4mFOiyCKbPMkgYzCz/O5dALoFcArkEbh4J5ITFzdOWeU1yCeQSuLEkYFbgfLLQN8CY1biBwSgugE4s+g0o53qu4XruM2ICIBaQgINzpgwYMcF9lrhms0U9QB/gsHkioOwA+vacpQ/XnamvHlWIoAn5tps3BPnwPN4XlMHAOZQrwvugiNu+DfZMq2sWMOc3rDNR2v+nQO1H+oVMEpT6z1PCYo0DOdi7yRQxA+4pt1nYkx9KG+Uk3i7KE3mYL/mxtI4WviFbNp6DjM3938JGmSwJE8T15IUXDGGc0FaNOEiLuv6RLae1AeeoC6G97NnZMFEot5y3sFNY5iFf7uM7v5kcjLgx2duDra+gQGLRR/0BWoi5TV7INtsvjEThPEpsVxtJu9q7JHaax3pO82lkSz2tPpQNmdNnLulISQueTTmQtXlYWIgr6ki/Mg8f8ufZ/G7jAoWcPFCIaWeUevqqlR8LP4DbbNisLOFBnzCPDvKC+CA/6mdeMVkgtC8rrCl1vHj+v11kWXlJcsgvvkgC1l+xZCVECoAp8xBjdCvCgkz+QZrT308/8YyB/AA4Z4wyngBYaKwTad58Mr/S1+MfeuiB8OnpNyWzE6/zjv+ze/3dDz3gf3LfN0arxalkqHvBXZy8P3JG9iy7vt/rj4uRO9ygNtwZX3gWr4Go0U26Dzz6dq+48Lwj4Jf+DCCUnWfpUxAR9DPGI+PpDUr0Webu//US+8M7dP2HlBgjs2metlHvZoT0JT7isi9n7GbD7f2o/n4v8hABFGv8h/KikFOF44noKSdJWNH5xHfdlue7u4WYTXme3gXadFv7iCRhGM4Xh8ujnpcMSaCHlMWCTp8ST0STuiIsLrug+Y0vSiDj7cS8zHsDEhfSgn7Mu2qrg/fltythyEBYN/qlvW95r6+TeBCU11PuqbeFQ/i22qO/Gg2vHA06wZAfLMwGtaXnSqXuUpx0WvFw5xzvFkKafU0qA/o0ITG3CvG0UdUIt8Vm9La2Y/wjH8ZJn1zPie/r2SO2fnbqZcHc+kEl5u3vYB3A5tu9dtOJBKJ7LxIWTEqsaTR+3Ge0/8OFTqP4jIiLk7WJ5mt1nnUMaybWGfQB1i2861hPMcbMYKjhF+Ldh1598uNPf+iOp+X1cLuIBPb60RLco/9ACrBuwagoexgxvlWleA+yLmIdw+Q5aLxCvz+qKlJXrZlcRcDyuosnxkeqI+1Wdbw5JMIC4o31lK3neefRn5kzqCf5G3E5qzI/nsTufhEWmtR9jHSyByTOXytBAg7Wh+vmeq3m3/Sa9be+uM/2+u3/U9/+UgmZW5iqreqe/5ZLIJdALoFcAjeRBHIN4CZqzLwquQRyCdxwEjCl3dz/zTLfgFMIiX7sVx0oN6YIARIDstk5s2Dkb/LkuvVjYFPt7YRgIDDgA4oUn2ug3spHQ2f16YZTvees443xHLMutNBWKGKUBUUFxeWw0puULJb5RiCFgeyAI4SkwIJxn5RB8gQoAeD7QiX+RhaAgOZ5YvIy8sZCDfG3bcxMaCPuw5qNc5QNEgUZ4t6PgohSZmSBydQsk83akboZCcI5LNyOKKEkUW7KaQRHlpSw7/p53RsBeZp3zfvSeiJ3ykEeg6GzAEmID2zEBHkNHuY9w/ms8km5AeVRAgkBgOwgk16MWfwiSG+KJ4ATJMxnnLhVdaKG7zQ+ZcSCebFkw2v148Bc6pH2S8VnTswrhzJR974lfCojZDXoRWKeFVxDuwEkWNtbTHYzdyRvG18U0Ug97uUak5vdb+3VH1MAq9ykMurrRZvTX2p18+t3LgHzhMGaFZKNsfvjSlhvAmiwF812B4AiCaCRA8CQsfVXSvQxxhMEKcQlbUxYjSfumP+ge2D5MRnEdova67T6qtN/JGylfMyLo0n3zDtrkRdEruuNxIpU1C6Onzh3+C2ni0PDvf1P/nbNay8Oe0JVlA/9F1KQOYK+SbkhXsxKlmcDgpJsrH/bdhVKf6f/Mp4Zo5AVhD3DstTCw5kX1A6zu2qXMW4JT8X8z0FoP08bkXd3TdbaU2O1ZVm1L8o7YlUht1Y834k0aYnMSMKCSAp5TvRWw6gnw/dQoHJF+wlU+kbwEr42FHAUzScUSdHQ5tw9hfZR1qVBsvaqVexmzzglEyKRbrwr6Fu8myHHACfxmiQM21bHD+lHEu+2H1b6Svqp8oNEJE/CTzFOCFN2zYiLjMcT47PgvH3E1kmMU0hR83SEXOG9whjmGtY5OxmfeDuZFTzyof9D0jFGIWFZE7Gmo+79cXot679Nm+U/by8BJhq82DCCIO2HsIjkZRFrTwW8LURmr4o/PalpivXDkDaYHlk+O+Jr34YvGZpsHJsZP0FYKNZLrJ/Mm5Y16qwSBj7mLcq7oqJrvd13zM0EpfDJM0/tZh043W0VTq1eGPqY8r49Cv0JjaDtyPytavZH+vEfKmW9jBkfrLNZ1y6oDF8jz4iqXorzitx33C9GioQV08/t/WweGrybqBfrfsYNdSH19RXlQfnp98iQcYAhAfuC/P/svQe0ZdlZ37lPuPHlepWr1VUd1N1SK4EsgQK0EEEkE4wHsJcYWICHYTywhoFhZjBmmTD2GC9jGw+DFwabaCEwGGkshGQJdSNQo9CoJXWsTlXVlevVy++mk+b/u3W+0qnXr7ordr16d59Vu+59556zw/+cnb7/F9gfGNEAri8gLPI0/UhvdfEWMUQiNl4wZDCmkAd5+sMj4BHwCHgERgwBT1iM2AP3zfUIeASuHwLrfNxaQcPVtwSitnlm8V8VOJsmtwmrTaBumuDcXr33gnyvoDUIBA8pselgE8DGibK6LuumLpZS19InGm4WLmF4sBnhOrSEmTMQArOB4DttMbdBJnTeSEDBOYQGuESBTEDIxd9o2SNkBw/+Jk/yYeNjbrDAh3s4h8YZGx8Ek3xaAFBM+M8JKc6dg2gwN064U0EQU7Xa4FryAld7HtTRNlrcw28II9G2ZANK+02Qrq/nySSzRuB+00Bj04YAA4EORAffqVOVcEHDjYN6cGyEG3WoEg9GYlWv53cELmwCq/UEP/CozvPUlTqAJcKVWdd7qu76x+bd6T9CiENdzBUB3zl3SIl35ooPrC3Km+W/fhjcmLaaNcl6IqbqZofbbKNr+JiVi21eOU9bq7/bdxPuVi1jjPC7AG9PVlzx473SG03LFDdfWEIgHKFf0y9wM/Szl5kxRCjv+3crYW1hB0LU31WCBHkqzNMD7WQhLFxImbN5EHdqWY9+inBpNcxSXLjIT0bnTfX+4tj4o7/eDIuU8QdhJ0QEJALv3s8pMe7Qt6kzpMWVHmiQUu6TShAsjDkQIH+qRNlDQm4zCD8rcSx4fgi5v6/Elrbf88r9s184dno5m55odSba9dX+ID0hcuJZuXvaJ5dQMwp2PiUCIq3F8SAMIAnDIYEpf1HNNM1WGzXFOc94D4oJWVnIJVSRKdZFlRS+Uoz9fesQKN8n3ESZlRrj5QeVcI3D+gBriqqAfj2GzOO8B5COCP8PKSHUZM2AK8Qzyptnx5iPhcFVkRdljJpqHUyhwRQqmLtoA3MX9YGkIDHXoeGN7336GSTD25T+rRL9a0MfNOsbq7//TAmtc8rFzdvvKGHdybjF2GPuCD1RsQF4N8Ep3k9zPfnX+v4d560sumuSpWvWiGNF6Ak+FzfHmvoc0xvdWZsf2y/LMMXeKbbJwuBQoLhIupc1MiQ5azbePfoTa9P7lehTvJesxxD03zF763x7Zu/SqtjzXGmit1afXjw+9d6jj+x9a3+1/i7pU1wpfGY5xP3UyVxqsib+apEVJ1R+Mb59bRg0XOTJ6eZEb5fOz6rMvj7py9SdPkTftrmOPoeVNHsD2rmHfITH87rP3N/SblNmon+gPPQCv1pUTBYsE3IFpXZu2EyIFebdRe8O6kpfA3+fR8Aj4BG4eRHwhMXN++x8zT0CHoGbCIF1AtENl+WlK5qqf2M2Pkh1rklLi48MtarQEsR1igUdRvjGJoTN1JR79mePulf+EsJ1NuJs/C2wrZl/QzKYqTqCNdt4VdtkFa5aDLDBIQ+EibQLASMbHcq2OBnmk5e6sdFB0MFGCYEC36kjwnk2ThYcG0Ek97GpMpdHlHNACe1RTNfJw8gOIxhMa8xiXrDJoo5ghCUEbqpoB3nihsbcaFUJBNP6rbYX4QV/m3Y3RAIxJRD+I4TkN+ZeM9U3YX71IVfzreJqZJZZ2nAdbaNO5Adm5rrKLEqq9xspAY4cT7nu8/e6M3+CoAUSg/PgBL7gQr5srr/AuxN8zXDDe1VHhbwgH3vXX1SQVfaLy+kE68mIq6qzv/m6ImCkpxG0vHsEBP6vSvTd+5TefQk1sMCk9N3qgRXGDyghwFTnUzH6F+jV08Cqr2FSBOEPBef55OGYwbtGfzgksoLxCoFs9SAGAHXjYNypHlh1MS6uPyBmsCSpHpAd+LxH0Mq4TNvpvw+W3y346nAe2CDPG32KMRHXJWYR8613Hdj+iGIGiHvIu2vdwQpWFnIBtabviyIixqPANSX3K5r1aEWBzIsszVoiNToiJVYlrFro9hP9mc0V3WK53RLRKaJ/eS3NpybMuO1GN3nrlS8iYdgHRQgw5iOwxUqJAzcs36b0wy/Sat5p1gsQdhDHvP/MM8xF5GNxn44rf+Zpc9/HvFWd+6oWNOvXEsxDVes8I/75ZD3AGoI5kWtMAYP+zljw1UoInxGeMg8Ti+OfV9pj48aLNHH4E+Qhlii8iLiio49C7Bhh3itjhARXS8y8VEX879cHAYThb3z7u3l3WfvyPkGcD4/+2rKE6okb376nXeT512lcOitLizslnD+b9ONHFfvB1duDA/qb94/+hEsoC+DOOwZBzjrWXBsy1nPNUBFIU1EuF0yRkpgRlzYne29vT3X/amr38qc+94F7fy0dxMxhvN9mJXs5IKB4Y8ootMvWwFrzBopfVizVW4NEVh7TnaVWKrdWy5oBm5oSI4UUYq3KO844z5rdyDn6NWtw8KLvHkl68d8snpjaI2sT1s4bWVJsSFZofTcIwvC1smRpfFGv63zzfl/fPlRi6t1BXc5T99d6BDwCHoEtgoAnLLbIg/TN8Ah4BG5+BF4GLW/GfHy+swFhE8UGAn+0COfYxHTc2iOrbuHPH3Az7xxTHAs2HWz02VQhHGADxoYJYQNCNtOSB3wTOK7XdDd3VggqyIdNDpsdNBQhCSgXQYe5SjKhBucR6HEPAgmzvKBs8oBYMEsBhBamhWtBBqkrrqYQQGIhQL1NmM+1ZiFCu9DgwqUJeaKRTX7UiXLYVOKeBeEE+dHuKmFggnQTvlggXPKC3EHYSdvBqmqhUd28GbFj2NmnERSUQf5Gctj1ZjkAdibUqZIdXG/ap9xj/oj5/nE5St7nwsZJN/9hiArKMpKIdwLMzB3W+0u89PHyHyVhtxkFti8/GDdxiRLkXewYPlsJNHnHTTv1kL4j/EE4SMBtxgAEkPT5n75MGNZpiVd51KKm4M4SuYSS2wyrcW+FG2CM2ugwsmKj3zYiKxBOmaYp99AmxhTcWGHVZWQp1hUIjRkzbTzZzO89Y/G/U8IlEAeCqvETZ1aWx9v1vkiG0+PthmJouzEF0e612nK3JaRlOcHYW5egSrEt3JL695osKeQ6TjgUxZoLg57iVyRJmvX0G1ZZWRlM+TIfu7/8MhHgXTNrA+YNiDnmzz9SwhphI0s7yAo7mIesbxB0F0sG3hGEncyxH1VCcGpuHyEAmK+YH00pgTrYusKsNs2lE2sB5nfmWK6HMPtaJQSp/58SdUG54PeUWEf8pBKWFJdCeFaaccHX79VfCGUZQxA6497HrEqpZ1XBxHmy4mIw3jTneV95d1i78X5uyzMto8QoRIphkWWJqzfHUUIxt0YzsqoIJeg/feLgzkcb4/1ses/yTgXj5n0xV6TMXeaiEoKPd8bcHNmaejgmKp1Rj+iISo8bY4N3yWrhgfHZzrNLJyeOiQxhXXq5chvWdbSJ9Sb5Q4LTB8t1a9GpNcQaT/ZW4nralBuqff1OPWlN9JIwLrCIZp/A9ZoXh+tie+dpA1aHkDvHtfr+ZNqPp+XOSnCFzGEQ8MxnlE2fpo9ueMjtVk+xK9byhEtfcFDOgTI/mxMvlpU/7xHwCHgEPAJbEIHLnfi2IAS+SR4Bj4BHYDQQkIb8gjTl2TwhkGbzzaaMDQ2aSwgC2MxMu94zNXkbl7AwgqxAYxINWuYLc9WEwIGNCwJw7jUtLNtQmAYXwK7XjEeIbsGT2QiZ5YPdS54IIriPOrHRYgOE0IPfuB8BBsnaYFpnnLPNmbkaQkOa+prQn0+rn2l7ImR8QAlyAr/UaLNxHQISysZHNYIPNnxVawrat5484Her7xv1HUENbq8skLbVg3ut3tW6XSBNrZTHxq1q3WHtoy3Uq0oYkZ+RFZw3t1fUizbzzIRL+ox75h/xN5tr8gNvfjtHXp0TqvKuzPLuUGF/eAReBgR4B3nfTIOfIhknDiihLYprlp9Qol+jQc2B4J/+yxiw/kDgyFhWOURTSEIelN0Za4svHhsZ81wVb8CYi9CX/kSbsB4hQ4RWjGtGUDB2XSAA3aAtN/xUxS0UbfhkpUIIi8e/6b67lz7wwJPJ/r3Tq3EUzuV58XQtjpqCWgFlXSvt5mF3kOxuNeNEGbS6PUW2kDpvQ/6gFM8ibEXBoswsjiZJrjmm0K+yzfDHy40AmPOu2lzw4/oOgYcf/h9Teqn9I3MJvvM5cLHIfPJPlLBMQGsaK0/mKBQB6HD0DeZ3BLhcT982ogLhJ8oTCHvfrrRfCUUA1hHMqxAp/6MS6xOOH1Gi/Cs5sCrhnYbEp3zqy7qIcg4pIXg26xBTkriScvw9mxCB0sqC94rjPMkMaZEMui5XfB3X0GP/4nxxbv0lV0jzz8+MDTr1tdd9w2PPyjoCSyX6iimQIPjnvWWtxrjPHGcEhJEXlGnzFP3idXIzFbcmu59dOjWxrDK4/nIPSET6FOs8U5ihLzKf8i4v1prJ2eZEvyXSYlLkxR0iW87IFdRpJdbOkIOHynpTPu0gUWf6LOvzCc2kr+6vNf761NM7iLmBW0awo99SDuW98CiK52Vs15FlRauzOBfm+Qv4CPYYlI+18oJ3B3W5j95f7xHwCHgEtgYCL7Xg3Bqt9K3wCHgEPAIeAUMArTE2+59TQusJwQFCQDYebDIa7tQfrrjt37Lb7X43msAE/GPjYNr3JoxnA89myATsFl+hKtCvavtTPkIINmxsYNiwURc2h2irsbFhg8M1aDGy2WOOMg1MhBForLHJ4jqECWYxYIJ86sLGjMOsINgAcp7dkFlVmLCf62gDgk40Q2kDwgjOsSHjXr7jVgahBRghCDHLhrKo89YdQ1/dZXnUE5w/XZ6rYmGESdXiwkgL+61KXFTbw3d+416eBfixkTSSwsgjqyPXWHtwS2NunrruyC/W3MrfgCMbWgsYynMxYRLvCPnwnPzhEXg5ETCGwNy80R95f+nfCHM+osSYgDADsgJCAOLt55WMxLD68v6uIyzsp3PFVMOtQ16U1haX0l584hPbonowjiBgNe1yiNX/UNaTc/QxCrY+NxR8vogFyqXU40ZdA7aQLiZMwzXQMZEWBaTFrXumlmUtcaTdrOVRFCrAq1vOXD6mUSVUQO3VgQJq69xMq1k/pSDbc/VGlCn49pOyrHhWlhgnOt0kUSDvq2KLbhQwW6Bcc5sI4Qehz1zBXIKLlh9UOqDEPEdg3fWu2KrNZ361gzUHsTHsgBRhTWBWgnberAntb7PCvBisRlbw+5WQFVg7/a9lXVA0oHzWP7SduZ/xh7l0s7pnuxgu/vzlI2CWpZ/RrViNnfNHp1Fo0F1VHItIqT4X1RoDjVO8a1hkfK0sLfr9tfpvJb1ar5jsvVECf7PQY01bPViDseYyGcz637m2LYuK98liQcL8VkNlH9I5LIhYH65ff75UC6vWfcyftkaWlVuwV66c5pVCzaaNsJYFIi3mVAJrfuZT5jf6L2tgiHfGBPoBczEBvSERxTcH82vz7UDxN95cbyV14XB/GXfDXLOtr+OaghWtKJh5d23+1N1pnywvOCj/Xyuh8EPb6Y/+8Ah4BDwCHoERRMATFiP40H2TPQIegZFGgA0AQgI24WhQIYRH4PakEgJ2BIBLbvEvpkVYsFHDD/XfUUKoYNqF7C64j78RYpgAHWBNMF8F2c5xnQWmZuPDpoTNEBqV5EeCzKAeVcsBBHzm353yEI6YpUTVzVOVLLE62XX8bVYHVh+zcCB/8mUj90NKaMeBEUQKLjHYuHEN9WWDatYMtNHID8uLeyFc2JCipYm7FDaMttFcL3xb/3eV2LDfquSFETFgz/MZ+ubXgfDTyAr+Nn/HXAOm3Mfz5hO8f9k98zMEIQWTQ0oIkrCmuFsJkoX2/oYSViYIXP3hEbiuCLyEy6hCLqN4jxFc8g7/thJCSnM5R9+kv2F5wZjyXUoIeHh3CQ5Kv15PLFTaY11tI7Ligi7KOHRYCWEm9UEbG4IEQT0apwTltTgwCLxwMUdfos8h2LLDtLNvSmF8xcqCtv1vSrjh4UCQ/XElxqfiyIml3p7t42fl8ilv1MOlKHTzURRpbCz0HIO83aqfbTZzWVvUammSHR/0s9NhMzjc7SWne4O0JwuN9Kff/aabEqPKs74pvr5I/2NusxgXzE+897+sZPGrsMD8v66wkeZaZ/3t6/en1yqICe8laxDmPdxIMTYw9zP/IWDGDZbFG4CsOC9J9e6ervAJ33y38W6wBnqPEuvLNymFcl0kt1Cxi+stERY11nd2fE355dMiK775yGf3PXnPO54+IssFYqegCINyT/Vg/qq6G7S1Y/UaLBUO6MRkVM/mJfzHvRqWwKzhrqnsJunVXzN/dOZ4a7Jf1NtJL8+CTHGHprSChEjBDSpkP/Mu68NPKdFn6fu4fWMtzhz8ZdP7lr66t9aoDTq1tbNHtnV6Kw0si2mrWWpZPBsFMM/PDDorj6yeOXZfliQwHusgGrpLpP89p+Qtmdaj4//2CHgEPAIjhMA1nfRGCDffVI+AR8AjcLMiYBYKbDIQrOOnFqEa8wECNYR8K27+gQddns5oZ8bGBAEdQns2KmxQ2HgguECIgKAQI+QrnwAAIABJREFUofZ6osKE7Cbc55PNPwIu7jfCAiEjwnU2Q2hqsrlBm5E8h4KS8ne0u4zQoK5mfcG5qmDfyrP6VDXSzIpBt5wnPKiH5Ud5tJHPQ0rE+8D8HUEkbieMeOB307S0/I1IgEAwDWo2vtwDTva7lc1n9bu5fKL+3G++hs0NFeftGtphrrIgWcwKpYqDXWvED5+QUbT1CffI3/8LfRK3A21SNqY8e37jXQB7hI48B/A3v+ZWZ//pEbhRCFjfo3+QjJDk/eY9hXjlHUYzlD5rsWgYp7AcwhKA/ohlAGMOBCMWApAOInMLBJYQGxB3jEUQvEcrZUEM4s+bPmLCz0/o+0eVsPRAwAJhwXVYgjHmmcBlq2pnI0yzA3cg/0TpydLKwp2YW+0f2Dd9Vg9qIMGb4lgUS5L9zSV5OitCApxOiqyoy63IfD9Jzypo97yCb3cGSdb/4W++9wWSrEpZ/uvLi4C9xwgScZMIYUj/o38gSP1Wpao1xdXUDguli8WQuZJ86ccoHzCvoS3OvIZQGgtF5j+IC9YlrEUYExg3tmp/vRL8Ruke3mnWQqz9sCAIJVFXyK/UYQmAlUWtNZZHcd2sYQ2bPRrp70r6tT2K4/BncRF8TlYWX9CPzC28c0bOMf+QmBssJtp6fNvqWe/QyRPt6e7U8qnJp9JBRP+zd9LWsqakA1FOv2TuYY1ufYd5j3MXPURQnJB1xGfnDm2bJo6QrC3WFIfjWQUAh2jhXnMPB1lBX6e/EMCeNoHBs7qvpsDdszsOnH187tDsZxQPYzII6sovsHnQ1v3DeuRZ0l5bOPX6NOnvAtt1B+vmf1NidEiffv35Yg/Q/+YR8Ah4BLY4Ap6w2OIP2DfPI+AR8AisQwAhdF8xCfqKZ4EAG81gNgRob6EFDGlw1nUP3u2O/bv73Sv+Z4gKNMzYWLFZYlMEiWGCdHPHZMVwTdVFExsaEzKy8WEDZH/zG0I9hO9sDi3gNoJCymUzhlASEsDy5R7mLjZ7bMyqxEHV1ZNprRlRYASK/W3uLvibNrGhQgDDRpJ8TXMMIScbNDZRRqJQLyMEaHfVAoLf2Cxa/hAKFmPCyBHuqR62cbW8aB9lGk7mAgCcTIBHmWbdwn12ng2ikRhWL36jfdSfZ/xBd+o9uDpAMMuzh1RB2IqwiZgl1Jd3A6KGvAZ6V5zeGX94BG4YAus0wKvk3PDdlwWGHfQXBDUW1Je/Dyk9oGTjD/czttD30CA1qyrc42FFgXYs/YF+T99hXECISX/AHYYRsIx15MvfVXdP1GVYxxHQzGZOqR5o3OO2qyitI4pf+N1PD165f3ZRbp66SZo3QkmzRFYoGHcQSJu3I7dRrl6PgjTLOgvLnd7Cci/Rvd4NyDpgN8mf9DcLfG0a1P9U5yD4UXhgDfEWJYg9s6iEILiYNcVGzbpUsgKFh/UuoJjLWE/8uRKWWPRzXExSV0hKhMjMpYwP9Hero7losxgVmwRuX42XGQHGbdagkFgI5s+7O+t3VpxcQcmNXRhGY7W+vph7Jap4C26Qlk9NrMgl0pxcK0nfJ39KpMXr9BvrrfWHkQ0bNk9ulpbzNHxEsTEiESDEVaMezGusD1n7sZ5kzWwxXnjnIRJZ01vcCuatjSw4qmXuUTlvXTg+1Y7i3O191cnd4hBY+1E/+jn96VYlLCro26YkQN+JNcvtyNNoXifrtVYyG9XSxbiR7hmb7TyQdGv7ZHHxTuHCeh5LisUiyxb6q8vLeZK8fgOygsv+QIl+yrqc5+At7DZ8Q/xJj4BHwCMwGgh4wmI0nrNvpUfAI+ARGCIgoXMh4TMbHQ580CK0/iYlBHdoGLLhYaOw0x38kUCEBRqIFgwWARKbItsEsZHgHBsirjFtMc4jDEA4yP3cg2CPOYdPhORmVYFggrIRDiIYZHNE/RBwUI4F4bRNI8J1hBQI9K18hA9m6WBtq2q/rbessODT3MfBptM2g3znXkz52ZDRPvNfjcCfw6w47DtlUncjZ/gbIQh/m2sm2+QZqWKbVfLiWu7nWsvD3DvZdWYxYps3O09+XGubUttAUwfahyAWDNnocg4hDkF/v69sB9roPCMsWCgbcorA438MQcG7wjtzrtn+8AhsXgQqhIZpgjMm2dEVocG4Zv2w2hAEmhx2n7lQO6xz9EmLo0EfXd8Ph4SE8g6qn5sXpetSM/DBfRxCNQ6zRMs++/yyw31USVwMY/y89+PP9hVUO0jSbDkMg3yi2cjnlzrBytogqNeiHLLiutTyBmcq0ubFalCdDza8Thje0BZs4DLKCHWe6/PqAxB9uEH7MyUEnPQn5hbm0v1KaGS/XQmtdQ6soZjHLyWY8Md03VeV92EFRZ6U/6NKWEORx0NKECYIcQ8pMfdhaUU9+Js1CWMAh2mrMyeux97PdyVIo/ih4M75G9/+buYO3k8scs67ElTMBddbXZCFxXApWCUrzkOVJtGUSIZme6o3HcYZa2As/aoHay76wkXdnImseL673Dz0yH+7Z3d3qfkWCfyrMdtY/5pVM/MTFoKMuSjcvFOJtazVjTUdxAuunRhXSfQ58oCMGLqrUv4zaT9280en3cSOlYmJnSu78izsKAC3xbaDbKRM+hZKLyi0cNwmy7htum6n4m1kImtmFHz7nvHZNQJ4t0Xc3H72yEx90FEYDvWqIk37vdXFo/21FcaBjQ7IROpIebhmM0Wci1zuT3sEPAIeAY/AVkfgRdn9rd543z6PgEfAIzDqCEgg/SvCAA1jNj5oZvGJ6TcbmWfcbT/9WXf7z3+bvrPxQdAAwWDkgJlqm9WDaV2yySEfNh7VTR3njGQwLWjyMNIDTTE2c2joIsRns8cmzPLhNzQl0boy/9nca+SEWSLwWI0Y4F6zcOA85SO8h7SwYNOcN9dJfOcY+mBXQmhJG6jHek3OqmCDstnMsXEEB/7mPrOKoJ5GQpA/bQV3E4ZyjnpyVF0/8be1xfKwOlYtKAxb2kvbqIe5zUJIw+abDeDj7qMBGuH4+GfTjCbdm8sycStA2WdEUvxDK8R/egQ8Ah6BjRCAkNDBWEeco/9cXoPbEIR0QyIIwoJjA4F9lYytjmkbCoxvtMD+er8Bwocx3Mj1Fwjqbob2i7SwuRgBq83hzDMISZm/WVfgIoe5iPmR+ecrlbBkRPAK+YDA9f8pr0GjmzmYd+KAEoJkXFlCUDC3kifzMnOjWUs8p++QFba2MFKCz1Gxerrer+uWzl+EBe8xlr3ERPqR9Y1tz+xwrclZFzfH+jISW09cDKZ2rfzha7/+sazRHpySlQXrr7+thAtODgjxaiDsavbLIg/+4PQz258+/ez2t0nY/w1E8tE51m/EWVmvaMp7TxwlLAIh61AOwj0b63SzdKa/YOEwtHKoHNV6QDaitOLkgsrtufvUokiHx2ZvXRiXayj2BfRlxnMscKlLoDpNyDJjWzqIm52F1vjK3FhRFCH9elLuq8ayJKyJ9EiWT48fXzzeFFlYe1eRpy2F2c5lqTLeX110WXKBtyf6JrGQcK+IUg3rfFNAciKS1lXf/+kR8Ah4BDwCo4CAt7AYhafs2+gR8Ah4BC6OANr0/5MSmxmsK9hIQRRgVbDHPfcLZ0VYsIF4t5JpGyM0MA0vBORoXB1QMosCBPYIEWyzYcJ/hBgcJkhHOMN1bIAgD8gLQQTCBurB9eZLmg0TZAUbNCM9qkGwObeenCB/7qMe5MPG0QRBnGNzhXCfTR5l8d2sQCyYN5qibOw4TLvaXDutt3ZAMkce5nbGCAoTlFA/cxXF5hDBHteDJeWjVWYYVskJI2KM/LB6UCez9qgSQWCH8IY2gysCHHyCIxxCsw7nTli08IypK5tQ2gi+ECm8E/7wCHgEPAKXggBjj2muc/0tcvE0E4WBWa4M89hA4G7j50hotF+ChYVZydnejLnCXB5eynO44dfICsPm1zWRF8xtvBfM5wh1mf8OKeFSDe1ySAr+Zo5mrkJo+n4l5kEw4O9fVUJZACID60t711gzwJaZyzazAmVutDn2AuxeJKj4DcfNV2BzIVBaWbCG+vdKrKEgZM8TE3Jp5OTLztXS9HhjbOKkvvOO4laVo7622Po6WUg82BgbQB7wLrP+soN19EakBf3juCwdzhx7bPfsyumJhr7HuJnSAWmw0UHeb1PC/RrkHX0Jwo++QRmsK0n8vZ6wYJ3IGpi14JCs4FC93cmndk5PLq3sEXnRFXFhijSsH39Z6TWq02Q2iMZFTCwtn5k4M1ir310fS8bk/mkmrme31FqDorPQfjwIksPtqdPBwrHdy0XmjqSD7pf01pYUC6Q3jAmy7mCfcb8SMaFYp54nKzZuuj/rEfAIeAQ8AqOAgCcsRuEp+zZ6BDwCHoGLI8AGAc0v3EJBAHCw+WIjg0XFO93Hau91X5Wwu2DTg2DgQHkdcwgJTTQECbYJQ1DBdSQ2feZyiduqln0Iy9m8oTmGdiXJXEaxSUSowd8IvixeAwJ98sMaAIKA8s1VExur9dYIbAI5h+AE4oRryY/2ISRBOMJmjXoZoUI92SxRFiQB91COubKqunni2upBnY1gADNz88T94IPLDDaUaJo+XpZBfWjvV1Qyqlpj2GmzqODvKo58N/KBelNPiB++o3nH5o/ynnAPfyNtxW0AzxrBERtqsOFv2otbjfsr9fBfRwSBUlt+fWurVkv8Zm6TXoCKadKPCFy+mRciQMyK4TF8QYrilg88cPAogbc9UJeFgBHQzDtmecj8ZeTFZWV2Iy+ukBe5yAtTNKBKEPXMi7hoYs7FbdSDSsxbzEXMocxF5sbQ/PSzrjAsyMcEmkaSVIn8G9l0X/bWQID38ZDSP1Pi3btPCWshWQb0XW95ATdHt9WarRMhkXiCLy7JiizcsbbQnlHwaiyLIARYI7MWJU/WrvTzalwL/MUdlyuojtwoTYqoeFIuli7FVZohjeIPCie2jmXtTTlY8bLupK+QX9Wyg37Heo/+htXT0EWq6uC6Sy03NtNpKxh3Q6TFYbl8Ih8wYJ+g64rpLInWeqvNs2FY3DK5e2VWliD1zmKr1RzvpyI5FuN6kifdYlLxLLY1x5sHzzynCEVJ4rJBX2VkShcYkbF+ZT1u1lGerLAn6z89Ah4Bj8CII+AJixF/AXzzPQIegdFGQK5/OnILxc4B37FsqhDgIyggUCDa9g2Xp2Mu6/2Ni5pocQ03bDrYGLH5YpOD8B/tLQgDhBBs0hA8IOjnHAQDVhhGbKx3BcKGiU0d5bKJIl8E62hmYv3AXGUWD5RNflg+QHhU5zET9nCNuabgHJs3NkRs1iibehlJQf3IA4GKaYEiTDH3HFxv5EE1T8qoEgj8zWFtM1LDCBTaxvWmPYrp+3uV/lFZL643yw3L28ozTVHLe71rKH63jSi/IRDiWjajECFg+DmXdWru7AfBweJy8IzZhIIF5ve8AznvhDXGf44OAlXCQeQF74+5frO4KtUYLUNgdI8XSI/OK/KClvLOlEQX4/b9Su8oGS5IaMjZLRmP4koe+Uu4dCIwuY3vzAMWJ4qiOF/T74zzjN3nXRtV67GZXUaV8V2q1aUNrBWqhKjNpxD41bmV72uXELzej0VX8mL6ezZEQFYWmVxDsRaCjH2PEutXW/8O3RklvVWX57N3iq0wpRnyWhWRMb58euLLdt0x96wCUZ9V4G0UQ4yERCGI9SBxIFC6oV/3ZLWwnPRqhQJsL8jN0qM69/WX8WjIg/WwrRlRikHhCLKPfkb9WJNbDDjKZZ3OGpBx+mNKEDJDK5I8C9zCsalPyh1UMbVn+YhcW70hCAvWrvepZ55QkO0nZIlxW3eluUdWFnL9FGRyD1VMbl8No0Z6OEuLhbTXD3srRTPtp9u6S2e+ub9avCJP1UUhdgho8cUD6xPcVv2REmvWCyzzLgMDf6lHwCPgEfAIbEEEPGGxBR+qb5JHwCPgEbhMBHDD8D1K+L1F45HNDwSCBY5+nXv+lz7sDvwUwpIDSmy22NggdGAThuYWgnAT7huRwW9sitiAbBSHoWolgIsH8sQ9Efli3o42F/eh3VVVx0K4b3EyaKqVZxqWVVcjXEd+ECoI56mL+fNl80a9qy4kLBaECUzWu1yy3809ls2jVQGLWWdQZ/MjTNvY/N6u9D4lLE8IHAopQ72J21F1+cQ5w4w2mmCHc5RpJIbVh7zJk/NsVqnDlygdVjrnCuvkb0NkYMVBu9l8Q1RAJPHMwQXSgnfBHyOMgATQRlQYcce7y3vFe8IYYORbrms5n3viYoRfmHNN5704ZCgomPbYtql29IEHniR2xVDAXgbeHlmgKvE+DIMLpHb0odJtFHhZwHjGarPag/zhvM2nF7V22owgX8Ql0/o2VDHxBMRmfJAjVKeStGA+ZJ3GWrFyFC7tdVxv6WwtnNl5OKrVIQjOW/wqWHa9s9SamahlCxL8sz5jLcwcytqLPgzJi1VxIquGg6ee2vGQgl7fuXRqcqCYECizoGxyqYcRFXY960WUej6nhCsnXKphact4wjhi1lusFSFQIC0gSX7MMhB58i1nnpt9QmTFw7teefrTkztW36FVaCJipZ704l2yAJnRZ6O30uwPOvXFsenOvu5qY+XMF3Y/Mb5tbizPlm4ZrOW3d5eDPf3V1EVxIN2nF5AVD6u831HC3RuxOMDFW1dc6lP313kEPAIegRFAwBMWI/CQfRM9Ah4Bj8CLISCN+s/KyuL7dA2aTmyoEFyjgYVwBKHlIXfsV3e6/f9HQ457uYaNEAebIqwwLCaFBcPGtBtSAIEDmyN+5x6+D83Oy9/4RODJZsuuf4u+s3nCagNBqWmurd+Q2cbLhPeUySaMTSECVbTN+DSrCjaMaIhxUG82g1yPKb1tRM0qxNw4GWFgZERV45xzVbKi2hYjKbje7uVa2gOB8MayLhAIt5V1QCi1XkBjpIXlQxnU2eJcmLCHc+a/mO9shM0qhTacksrcqnvih8H+kBLPgk0h+KB9Rz4814h3gUL8MXoIYFVxdrETrXUHURSFCkEQKNhn0YzCcFYCaPpupJ7T1nneL8YG+py5ufDCxdF7ZaotZqw676dd7lGWpica0fxSh3HNC6HOIWVWS1XcjHi2oOQ2ptO/GOfpYxyM6ygQMLcwtpuLKC/cG+1+51t//RGw9dVvqCgUPs7HgsCtUW9lYSaIomxsZtdiEIbbMSAQQbHamuylcpvUWJ1vH1EQbvotlq4cjImsBVl3/okIgAMS+h959jP7J2S1sL/Igu/RucshK8hzI2tfzqPM8y4liAnWnriJYs1pijy0DeUk1stGYpxfa6v+96zMjf/jva86iUIRa+WujCOOLp6c+tjJgzvfptgVr5R1RRFGxUrSjXsuzGrZIH9NniYzsq545cqZ0K2eFcvRE1khq43yYExjDfGAEuMcZAWWFcSsucBPlN3gA24bEv7TI+AR8AiMHgKesBi9Z+5b7BHwCHgENkLgj3Xyu5XQeMK3LpspBCRsru5xg7kjbvGjn3QzX/um8mY2SOa6go0OGw8sGEjES0Db34T0RlxYUOyqz2nbxXANWmxsZLA2wB+vxbAwIU6VALA2sMmhHMgGNoVVbVS7HsE81gTUFwLDhD3cxz1VV1D8tl6wVCUsrFw+jVCw71WXHlWXOmbBQX3YiKLxhnstSBSwQuMOogjyh9/X51u1GDFyyOpE2w4pmaWIkRngwTPh2Zx2p9+D9hqb7QNKbE7ZNHIP1isQROTLO+CPEUJAGt1GwrmDh+eiZi1u9fppe7xdN0JwUt6523VRGGhXxlE4lYcuL0kL3tOhQFpkB+9a4S0tRujlubCpFq/HzvY1QJk12NA9Xmk9sCGxtZndGV3NEy1dq5GFuRg0F4RgY1YUw/lQ8T6qLtbAC6yYT8GWw8iLagyl6vx5NVX193oEPAIXR4C1K9YK9yt9Z/WyPB24weri9rjePNwYn24FoetM7Fj9hAiL19dbchvVj1ECObAua1sfPiJrigef/Pgd473l5v+g2Bf3Xegt6ZIfSdVauXoT62gsKDgYZ1Da4RMiw2K2YfULmYJbJtyCsv4eHpAvcV2+nopgl9JArq0I1XF7XEufmt69vF1WIUsrZ9udMEy3DXqT4msGje5Kuu/009G+uBa6rqjqbABZgZup89VizYBVBXiitEMst6GrUhETXvHhkh+5v9Aj4BHwCIwGAus1Vkej1b6VHgGPgEfAI3ABAtKsR9sJwTXzAlsLc/+CBv5Ol/f2uUO/+DqXddlcIDhB8ILgG00thJt8Ijxn44FABUsHNkqQASTu4RMBDH51EcIgsGeDwuaJ7wju8X2OdcdrlNDo4qi6jTBhPpsuyjMXGRAXlGmBv6vEg1lbUEfyMuGRESdmycGnuVhig2q+wm2urG4KrR52jX2uJzfsb3P3BA6fLzHgHBpvlGWBxcm3qi3H39VzfDcBFlhC8Pya0t+UeYIBGoAQEee0dHvHj7pHvwc88aPMbzxT8uAZm/uqz5TvAHj7Y3QQ4N1uNevx9Nx8Z/viSn+bLCy2rXaTXf0ke1UYuDdI0PDqtW5661onuX2tm0QiNJppmpOMgKSfD4m0ioB2dBAc8ZYSx0KJceQjFSju3LdzkjmC84znfL+YUG0rI0ibaTvjMtaClhAc8p2+Y7GYLug/pQstI/sZry0xrlfnJy/k28pvkG/bDUWgFKLT91ACQakDa4Pzh6wQZUHQdWtzJ/b3Vhc+lQ26H5blxRERFp9vTXXnZ/YuoeRz3vpM31l3Er/iiEiACVkqdBZPTL1JsSvecIVkxYvhY2QF17xaCeuK6hqSNaCt31kzmnXwME/qM+jWnSw/5pT+m041Fcvilm23LP79bbfMj4VxZz7td8bWFlaay6cKxb1IxlfnlvZ1Fvpu+bSCdy9q+bkadAfdQEG2z1cTd1d/rsSeAxxwVZV4suKGvua+cI+AR8AjsGkR8BYWm/bR+Ip5BDwCHoGXHYGPq0QE2wi/36xkbpYQrkRu/iOvcmsPz7vJt7B5Q8COgN8EMlQWgTjEAUQCWlRoT7EZOnf/ufOQE0NtbCU2U+ZaBuEN95Inc5MFkTaBvYFhwnwEYdQDawXM3c31k1kqkJ/F42CjCflBexAOGWlheRoBYG6ecG0FmYAw1+ph5Rp5wL2mJVu1BLE8q646jPAAAzaFBFMEBwRZWFgYabCeEOG+c654ziXKo67gA+nwlNKfKqERZ268qDeYkCfP4zE3/6doz/E8eWYWt8Pia/CsuZZn748RQaC0rOD9o79tk9pknufFjkGStpuNcCZJsluLvJiWlKGRpPq/yJ+vx+Fqp1fk7WZtZ9hS3wiC5bSf9+q1aKp0GWV92frTiKDpm1kicLgclxiPf2Z8rPF7+mTMZfxnvBupANxlLBjGasgK5p8hYa5jSv2NeYB5iTGeOEII7Ybzo+7LRAANxXsV0sK/ZB4Bj8ANQgBhugJwM5Z9tBzj/rY+f8SqU0ganwy6buXk4cZgrHF2373Z4vYDSxNyDbVHFgkoieDiFKtjI/dnRAY80ltptBaOT6V5FrJ+M/eKD+o71rCHlBgnGD+u1cEYhLUxRAExN8z9KetlLC0Yp21tqok/UHDx8Gzaj+N+p75TBAxrxSUthutRLW02x5c6SbcYzwbpzkF3dRZrE+J65GmmRbaWs+eoVLPk4PtfKaFUZGtz2r2hG6hr1WCfj0fAI+AR8Ajc3Ah4wuLmfn6+9h4Bj4BH4JohIA37g4plgVsmLB3YRBxSukMJQQobmhX39E813Os/PCcnvWy82I4gnDRrA4Th3FclEdCuRSjDeTY75MN1bIrIt2rRgeAfQTw+dbmG/M2tkwnYaa8RC2wgsTKAGIHsMIsO5jaEsUYymGUHZAWHlWlEApsnrD5wyURbCITIRtFwMPN9y89M6s3lFRswyqBMi3thxIaVwb1sFmk35bBpJFi5ubHid4RWXGNun/iN68HFCBDwZuOLlt8hJTadCAohJDgP3uBC+fOuf/Sv3cEf+yp9x/LF4ntQ12eUXqVE/Y7z7PXpjxFAoOIGinc1l/B0T5bnsYiJ7fq8I47DMQkqxs92+5P1WuzarTgROzEuQmNJv++qpeEgzWInB93Lg0G2OjPV2q3YNsS24P3F4scTFlfwHpUuk7izalF1Xnv+JnCbxFgCWcExpiAojDNmdYcwbjgPjELw7ZKssLEdsoK4QQ31IbBhnrhNxEVXfU9jdTGmT+ZM5hHm3zXdn3j3alfQifwtHoHrhEAZgBsBO4QCa8nzhMWwSDEQeZa9td/p3n3m2fQ/7n118ey0VrJBJJeq59ai3Ef8MtZ9ne5S68NPP3hbf/nUxB2ab1lvMh8zNtxXNgEC4XocrC+pU/WgXBJrR9bCwxgacgEl65HabJ4HLbWgq5gWHwzD3KWD4nVhlDzTnBg8LYuS+/I8nIWoyNLE5VpIXOT433UeK24UG55TYq1fVey5Hm31eXoEPAIeAY/ATY6AJyxu8gfoq+8R8Ah4BK4xAu9Rfj+sdEQJQTgbFzZpbHAecgv373edxyM3dm/fhRECKROmQzAgMB8KY5QQVEEgIBg/oISwnN8Qypggh+stfgS/MydRHtpfb1Bik2cEgJEMZoXArgghO9cjpOd8NT6FCf1s92QkRpVQ0C3DA2Ea2q4QF1gtmNYr7aDORsoYYUH9zWUWVgu0ifvNmoRNmGmumUUExANlk/c+JQsMzgbR3Fqxaa1aY1h55F8lYcgfvCA3ICPuV2IjyGYYTM/5Kc7TQ+7k777FZau0AazYCOOCit95tmy6qT/P3B8jgECFrODdaSi4dl2C010SmIb1WthO0mJ2tTPYnmbZ+CDJJ5Mkz7M0d3Ec9Zqt8IAEF53ltd5TnV5yQvEsdmd5cabZTJfHmrVAIdvpR0O3Nl7Yemkvk55H1arKrKh4NkYCpxLwE88geLEYEJS2yQgNxi7GLcY5I54tXsoouDCy4Njj6l871OADkmfh2vj3AAAgAElEQVSOS6i5Xd/DoCim9XejCIrlKAgQ3mk+KdbUD5kLTOOYOcMfHgGPwCZBoCQtUJJhjfpbSt+7vmpFVsyefjr8occ+UvvJN377oN2cKG6RlUVNIzpjIX39qFxBnTl7ZNvn1xbad8q6AmsNLG3PB/PeoLmQCJRrgbuvByKsK5nDLSbcQPXc0VttrCydHD84uXMplqurXS4qYo1TY0nfTT/9ifx7kl5/Z5amilXRx3yMejGGsa63A9dPjGmsrf+6/J2/R2EeuB7PyefpEfAIeARGCgFPWIzU4/aN9Qh4BDwCL46ANO0Py8oCQTZC7rcqQQiw+UBDHx+4Y+7Uezrutp9nc4MrC7TFELAhwEcgxaYMIT15EKsBLX7+RvjC75xnU0RCcI6g33yd853fydOCuCK4MwLA3EPxSX5fqoRQjIDSBBfEyoINHZreRoBQbyMz9PU8aWBkAJsrykcznLpDOlBPtGKpgxEc/G4BC6187uM66sJ8yjXcDwnBfWbKTx1pAziBGZtTuw9sOU+7zZqEetrGEULB8hr6+lWiTdQbsog6Qi6hwTsUQitBSsRucPKEe+7/Bg82wuTPfZRtz5R6jfHMKdAfI4MA7wnvX1u+nppy5yTrCLcjzQq9Q8UOxaaYzOJwm+JaNLOsyJMiT4u0yONBrZ/kaSNw4b7mRNyT0OJ0ux4nIjRO9wbpfLMR16IwpI/ME4TbkxYv/j6JgDB/4YwnjB/0/6o7vKEFma6jj1eFO5tV0IN1gB206XWz0+0/P7vYMZd2jF2bte7XrPNXrCuYC/bKqEJEX3G7+thtgfqaRvNELmRS9TcFsy1mgziSS7ZCRHNwMAyHpAXvwKLyWVAf8tZK1+zJ+Iw8AleHgNxCkQFrOYTvf6jEWuqbqrkis096wcSRh+O/J09R43d/Zbrcmiq6Ua04G8XuMQXl3iWLBCkBpRO4hBIpwHoXV6zrD8qx4NhYJldJgMttCPmYxa65aLI1MHmxxmR8hlAZxh0SObGglXM96yennvtUsLh2tvXMnW8ZnEx6Ll+dD2bUvrcsnujPpANlfWHwDasnyjO/qIQ7LNbGYMa61VtVXO7T89d7BDwCHoERRsATFiP88H3TPQIeAY/ARRD4cZ3/10oIyAmCjTCcDQ+bpq5bfjBwvefmXOv23bKyQKDOeQQrCMZ/X4nYCVgnsGHhO5YWpj1MkQizENxzn1kUmBAVITounthMIfBHKG9ayHYteZjLJz4RypP4zjXU2TZg5GuuoxDaUw8LAE4ZbK5oG9/ZSJl2GIJ9rBbYTPKdwzSE+W4Bh6kbRAdWHrhD4TzfyYuE2TvacZRrdbX4GFUCpixi2FZLnCMv6sQ95g4KwSBYY6kBCYHbLnDjWUBe3C2rivvdo3/vjMuWIIw42FhbnZ/VdzQEEVrzrP0xWgiY6x7636qEqLxPilnh9ssHhN7hYrLfT1siM2K9iLErwjxV7MxOP03EX+SuyCLdM6GYFs8mUZbV4iiWVUa2a/u4ZLKFEwHCe2h9arSQvcTWlpYujAlBLQ5bSZoHwm0ycMH0UAM/cH2lVeBMs3y91v1mFfgM/ZsrWaDX7YpvYuOqEc+XiNBNfdmQlNFzC2WFNDa0sCiKeu6CySLNG4UrVtSLVsVYiJtw00EWDOc4PX/NDzJ1Cl1dP/BurJbxLLY8yXNTP21f+VFEgDGZeAzIUbAi/tEqCMjv89R95dEvxG7uUOQmduR/LKLikdW5YLDzjrxQgO24vzbIsyQ5HUSxKdhshKMp8zAeXA1hYevlqjvUKmHB+abMKZm7NQhF27OkN5cO+hrPg0FvpXf3U5/IJw9/tomSw70E0NYYJqsKXf3CSOFY87J/ABtcl36qXA/0ZKHi41WMYm/xbfYIeAQ8AleBgCcsrgI8f6tHwCPgEdiKCEjjfiArCzZj36mE8AlLCeI5nNs89Y41XHq277rSHW3dGYq0MA1aTNYRsLPpwSc3BAHkABpd5kYJyNi0MP8gbLff2DBxLZ/mbokNFcJ+6mAxLGyThQAMQQ+/mwUH2yfKxrUSv6HZhVDfBGjcaxYV5jKKe/gOOWKkC22AhIA4uVsJyw3y4X7qYTEizO1JNeC3uX0ycoB8zVrC6lzdtFXbo0uHJAfnqAtkB/dSf4gIMARjyAcLnk1dICsgNM65xsrTj7jn/9Vb3eJfEpCbc+aOik/ahDUKm98/4FlTqD9GBgF7740Ua4qDkLg8mpKINFLnk4A1QGCK2EIhN91Agbgnwzgc5FILFyERJplrNdN8EDfCvf1BdlqC1sVGPZqWJv3hndvG9I5KNOOPiyJQuoEaWlJIoK/4BW5nvR4VwnynhEHbhLNcbzh9uJ7iQKw1avFp/bGapBl9n3GJMQ5XUZtNkG1jq7X91IkzK4x11LtKPG/1t4O+FWZZDvM0rTQmd2lwfbKsGI7r47Ji0vN2sQLTRooLI+4vbOlhNrKimMszd7IWB8wbzJ+Mz5uVoNrqz9G3zyPwYgiw9vwLpUNKrA+/o3oxcnzFoHZr8/IFNR/9Hf32Jp1bWJkLT2mFNx3Vg1um9hStWuS+boNCGOOZR1nnXZCt/rA1JuP/sXJsZW1u69yL1ZlxqUp6MBaZYo3cVBXtdNBr5YoeXmuNPSayYvtgbSVIemt1OYa8XYG0b+/R4vP6QxtxFe4xXUAMOOrFJ0pLrGE9WeH7kkfAI+AR8AhcEQKesLgi2PxNHgGPgEdgyyPwx2rhlygRAJvAzgjL2XhkLmrVXP/4dhdPtRzKv0UjdVFkm5+v0DUElUZrDCEVWtwI1dlMmZsnNlpYLSBQ36/E32bBQXn8hhCeA4E7v1fdJZmgztxlYM1h1hNYWrCho3wCW1MXyqYuCNQsmLcRBQj6IQYOKGFJwqYO6wM0w16nxEaQvI1kMPdS5vrKYlSwwbSg1uayCeLELCOw1LA511zBlE0cflh9rK1mcYKwj82ftemQvn+lEniBHcQQmNG27Yr6GLmVh97gnvkZ6vPOsj1sSimbZ8GzJD8sXHjG/hgtBMydGf0ikiB8OQ75KHoSqKI0WcQxQbZdX+fG9HLLmCIoZEQhf08BfbIpM4q8Xo8HSjMSZIwrAnd3Yqze7HQTQgobqbfZhOmb4imXZAX9H7Jih2KIzEhwfZvoiRURRPIPHtwpV0G1MNaYGbiBSIxVPbCpsHBnwjBelhB8NQxDSKSMmBabjLRgjGYcMpcj3W+67273gQeeZOwaErGbrL7X650YEhaMt+pYu9V/9onoo3O0ZXUxKYKipXNtWdOc1fMVOejCIpBrvsLVdf3tujZVR8z0nM1NIXOAPzwCHoHNhQDjGhZljysRUJo15gXuoahuxQABa+NXYJ3AkWf5p9T3tVYUTV1I8aYoOjKvgvggFsSiBhHmhFfpj0V9Mq6ynrW1MmNMR9c9rDFkWtfs0Q9dfWfsLWPLFbJ0CCiTteRG8p6a7kuUt7w+5k9l6WCxv7L4VhEU+93i3MEs6d8lExDVzryivuSU/j6V85wSa+eHlVhXs/Y3JZzN9fR8bTwCHgGPgEfgpkDAExY3xWPylfQIeAQ8Ai8vAtK878rK4j+r1G9XQtCNlcG9Sqlb/ULius8cdXl3v4u3jbso1oYksoDXCDW/oMTm7YASuxw2TKblj/CfuYfzCN4/pmRxJohJgXuaoUBPCVKAzdfQdUqJQHXXZLEdzMICYgLhDvlRZ4iHQ0r3lefZzJnGKvmSl8XSwE0S93MN5ALtQEMM10tm4WHX0x7TJuYcm1buoVzaRn1xt2Qkg8WXKJuwYVusXUbMUE+00yiH8nkWxBR5S6Vs8KGOxA2g3Q/LVVfgHvl26o4VBa4KqD/1AY9Hldj0YmXxX3jGViH/OVIIfJF81HsuAXlbZATvLsKLoaRVmt5jcmdTFJlLsqBICnl+KsJoujfIRGC4ibVusdsF+YJ8R+yohcHeKIrmZ6drk/LV39PbRn8M5c4m93EsXvBeDS1bWs1aQ8KiKQmub5OFyoG4FnYVwFz+zIv9sqqIRFjgDmpNf2/T85mV261DuvGIyKGWnsvqeLuezS91UpEW2SYiAWgbBCpjH8drlQiyau75XlLitUV6ITgQmFaEnvypCQ9iVYgO3C7RZBDL9VO9Fm+Ta6h5PVtpLxfRYJDWRVCIhsrHW41YQstgVffMKY8F9aPh3On70hZ5O3wzthICNrZhzUu8Botj9t+9VCPzNPmHi8efc+3p7WmtOVZE9eY2jZTSAUh6jPsiCk7H0gMo8izO0mQlqtX7YRg1dYGIbFlpuCJSJJxbkn7nFNfm6eBoY3xG3pwiAnyLEMmeZ/wQCXKrPMxN6JM14AUHhWkeynsr82/tLs9PKT/dB0lR3P4SYZOIk3aPEnEpsMbmeL8S62iUIdgvjETMopd6zv53j4BHwCPgEbg6BDxhcXX4+bs9Ah4Bj8CWRUAC7b8WaUE8CASQCPIRcJ8Tfi98XHr935O5dF5e1uUSKh0/6uImwnCE61+uhAsjNnMYkaM1hsa/EQ9oXiFkZ2ODdQS/IUznb37D5RHlHVBCyEWqBt42wZcRIcxlCPaRtSKspxz+flAJiw+sJLgGAoA6mgsn6mckBO00X/Fch5UHbrC4noO8qSf5IEBCc4x7P6GEFhv1RVAHEUJdzS0O56inubTi076XWQ8/yMuIFja9ED4WnJz6gA1/ky8YH1bCgoO2sBFdct3nl9yhX1DNThjhQpD0c3FHziWsTrCseJxnWy3cfx8pBOgPvJO8R7PS6F6SsPSUbClWJCxP5KuG+BXtNC1qjVo0p7d5SUKNSb2gcagvulYObZzU/CVhb8aNei3cLsHImTgO27gxUp70o1ERTl/2izM5Vq9ryKzLWmJceE2Cm1wCvUICbbkPcntyCbSlfTsnmZMsW0Jp3ec1dfo7xBTJ+CVclSZ+0mhEnR3bxjpn5tdsDLvselyHGxgX/5PSz5V5f7U+f13JLCxyrEI2OkS6XIfq3LAsi4FC0Yv7A49lERJrYiJmZE3Tq9XDJT336X4iAlDu1brdJCV2iTqL3KqFa+pejPsNkVcKbu9m4jhgPrE+dcMa5Av2CHgEnFMMho1gGFo9KCA3gxtrZda2rD1/6aUwywY911teECGRbqs1NFwwaHRW22gFZMngS1uTswS3IajEIBv0XS7NALlsaoW1eqpAGAudxbnbBp3lO0VYnNRF+0Q6HAvj2vs0fx/L0/4bRYLsak1uC+J6qx83223N08N1qTiKoemHLCraIjxcb2VBJIWWrTonssTi0l2s+oxHtPV+JdbHtBnrCtaU/OatKl7qwfvfPQIeAY+AR+CSEfCExSVD5S/0CHgEPAIjicBn1WoE9wi80dh/vVLTNXZ1XTxWd9lK4pK8J2/ccsXUZDOEcIrg0xAVmIbjVso2MQhKyQchDMJ5rkNwygYPwfvnlNj8kIc0vIbXkQ9Cd76bbbo9CMrjfoQ8EBXmkgRBLMJ9yAI+EaBCYkCEGHmAFqyRHMyFECVcj5AJsoK8zN8vBIRtwigboT/3oF2GWyZcMpE3h7kDMT/D1I2D8k2IyzXVtth3c2sFOYHrJurH/fgF/l4lcLBA5QfK3yE30Gp7SMHQv8Od+C02kkbQ2P20C2xpI/jyTP0xmgjwrvEO0P/oWwcgGaTpnYdF3u1nRaJ4CisSbCC5mJKQtZNI6zLJ8m1hGsgzVJg2G7H6giJe5MWYXuRoYaU7d3alt7Rtorkw1q4v1mst+pzzGuEbv2ANsUCyrAjFRtTkHqhWq4U1ed1Q7IpsRkRGOyqKFqKjUBYuIodcOw7kQiialvDaKSzCScmyDo+PNQiIXhehYW7xNsPbzPiG5q0djDuh3EJlehdGKQ5DIXdfqUgKLO8Oy9/Lk/q+rJlhbxiEuyVMTDq9JCd2CSYVcq0WN2tRS89a9hgyasqLeppnUzLRwB3iuEgq+qnFntkMz9nXwSPgEViHgMiMrkiLz+g060/WcD+t9Halr78YWCIH3KC35iAN4BJkRaEQZDJ01LiPg0aRE07kBEQCa2XpBsWYYCjuVPYaxZs4myeJCANN1bgjVV6695Wu3/0JK09BtIf5yTLDNadmnYgLXZaJFMETFVeJ/e7KmC/LzuVyzn/VCywxyvyYa7CiYB/A+vgDSqwxme9Zo/Ldu3/yPcMj4BHwCHgErikCnrC4pnD6zDwCHgGPwNZCQJr4j8rKAoH8DyohnEfb/yG39IlZN/320NV2irRIJ1wtqLvBUuTiiTPaHeGqiA0b1yP8R4BupAObG8zFzaKA6xCmYw0ASQFhwDUPKZkrJu5HYAPZYNYL5jrJBDmUgzAWIQ/Xs6miTL7jZgrygU0fhAnEAOc5R3nkBWkydNeihLUE5ZTehof1gTgwaw8sRtic4Y6JuBXngl1/0RLESAudGuZvJAl/89vQZQ5/lId9NwuPO8p6Uj7abriBIg/qzEEMCup0zopFsmZ36Ge/0T37cwgLaQebR9xQcUBm8B18afev80wrZfuvI4SANNnRcuf9411CECoF8GKXBBYSlIci4oL9CrWdSnaS6mWvZVnWStJc1gByAFVzvXqgUKGFa4rAOCthS6PTH0RZWuT1Zhy3m7V8ZrLFuww5Z31nhNC9tKaKcAglhJ7o9tNbwkC+x4tgOsuzMeGdKfryknCVFm02rWegeAdFVyTRouRIAbEtNMR06o3amOTc24X34vRkK/2NDz0x+IF33bMZCAHGR6y+7DBC2MmtEQTWpQF0k1+lduZqb6oYFWt6Tst5VqyKpOhq9qiv9ZKxTGyE+lwUS426VosSsU483naSpImsLRS/YmjNJB8xQVOzRTVI7k2OjK++R2DLI8B6DyUS1pmMf48oESvsjUrEV8Ptqa3NzoFxzqrBFegI9BkmdDD76hiIbHA9jSTDv84tMc/xDMP/zfr3oqASf2JomSECpLt4RoQInghZMp6zsBD5gSXHOYuLix9YEbPm/BdKz5X15wYUksxaeLh2FWnjLStfDEn/m0fAI+AR8AhcNgKesLhsyPwNHgGPgEdgtBCQgPsjIi2IX4GQE4H4bW7tsRU3ON1zY3fX0cR2/RNnXTy902VxW0G4xxTXAsElGqamgQV5wGaOPLCmgBTAaoFPYjPgA9jiYLARQ7qF4N7cURlRUY1lYd/5RIBP/hyYpls8CcgWCBQ2i1a+xa9gc2UCIcvLiAnyMQKDOps1B8QBm1Hqg7UJBA6/kxfXI6ylHOZXu4e8zMLCiJeqxqxt8szSgtgbxJngPD7hcbFlQbOpLyQJLgfaLl0YuLWDdff8v4KMgbDADcsHKXD4+7l2U2esQh7kWZa/+Y/RRcDckvEe8/7uJeinRCFYTCQDkRTqdWPSAFc07nxCgvJI8o6eJCp9iTp6/STHtQRBuTsK/twfa9X6E+3afFa4rD/IXKMeeS3Li79bhaxWYpFAEzKzkKbskFSticDIBoNgIk3zpixcsKwYugcKa6HGU9dIFENE143V5BJKn6mIjUxa+jXFshjs2TGRSUBeICjfBK80JKodjOMW72cTVO1lrYLMJQrZToTjtVrQjqJgVn2sXY/dIFGgbYLaJ0m2KNdQ8kuPHY1oqyAUYREGojMIuN7RPTYvMPYzV/rDI+AR2PwI0G9Zc6IYosDXwzXmnyh9mdJ7y89v1iduSDk+r7SjDJz9wtZBZgzPXhkXMCQoZJoHOZH2MY48VwQkiVlZrCtU/l6H61XW+v9WiaDirDkZg7ibv8+7+dN31rvFRdxlvbA9/oxHwCPgEfAIeAQuAwFPWFwGWP5Sj4BHwCMwqghI0P1vRFpAQEAiEMh5j1v8aNO175l0jZ2BIvXVXL4q2/O6XMUgXNdmKKpZ3AQTtpslgbk1wo0SQnVICQTuJuCH5GCTx+YIAgEhHdeZhYORC+a/3YgCIyJwYYV1BgfXcC+bKiwMOMjHLDTskVrepjFW/d20l00QaxrktAu3J0Y+mBsohHRVYqVqTWGxOKpt4VraSIwJyA82htSf2BhvUAIvygKnBSXIjL0uky+BpQcjd+gXj7tkhQ2yubx6nb6zwUTTD404rFie0TP8TWus/xxdBEorCwg+SD0EKrxvk5Jr3FYEbiXKFag+JO52Ech6Yi0SO4EfCfneP9kbpC0FiHaNWrwiecchCd3nksQtSXi+ImIj7fYGg1v3TOMC6MqkK1v8sbxy/2wgQbV8aykeiKTUg0EmY5WiLY1XxigFVM3HXaYfJNAW59uVZj4kRkMePZIYpiMOW3oajb5uSpOk1k/C1nirzji7WVxDYXVmB1rFo7rPUCiSgHlsXs/7uKwmbpdLr7oi4nZlddFQmhY3ETfr8XwcBT0pPOvxBgv6nnSSYqC+l9ZqIgo1sw5Fh94l1BYfGXzzthgCzH+s9UimKPMpfWdt+KdKEAEErTalme8u24/CibkXvbaQDIkPIymGa3nmf9avv1bWA6tkW4tSL9bLf6aERTQHawbmGZJ3UXdtn47PzSPgEfAIeAQugsCobiT8C+ER8Ah4BDwCl48Am5d/poRLpDk396GDrrYrcTv/7pirbROxMJG4zjNyun6rbM1bKy6axU0Tm53blNioWXwKhPJGJCDMR9jOxok4FOayybTAEfpghcEGCcGqkRL8beQCLTHrBNtQmXAfYT/Cfwtijfinau1glhGWH2WYD182aFxrQQhtk8bciQUIm1HqRlm0z4S0RlBw3siNan1tM2ukCH9bYFUwQOsdN1D8Dh6Uxye/WeDto677VN+d/F0RRw9g6cFmE4LD3EohOGSjDPbg/SuA5A+PQIkA7xzvB/0GYkve84vT4iaW5YpoVVEWJCfPOxKqZrUoWpOgY7/88ovCEKWRF/00zQYSlB9PinxequJLLlBciyLoHjw8l37rm9X//bEhAncd2F4cO7XclzsoOf0o5PEj72dy2JFmQ4JRGq1Bs58OAzZntVqcZDK8EHGxJoF3T8xGoJgXvV7fLYy3a4p2Xs+nJ5otkUeMMUaQ3mjkq66pGHc2g6uqG4FJJnJJ8V/yvp7zvJ7OYXFMM7JYEpGhThcEO0VQ1AKRVSI02opFEujvcX6KIndSLtgUVUZupBTIQpX3/elGPEFfpkfgMhG4iJUBc2xP8S2Yb20daG5TWT9iBfzb5VwMmWFr4a8tf/sLfaLQc58SrpneWX5y/uvKPFn3oajDgYvV1yrZOvT39Z015ZvL+2ytzDnimmGZy3fWl7YuP6zvKLoMLfqU1ltQ+DGpBNt/eAQ8Ah4Bj8D1RcATFtcXX5+7R8Aj4BHYMghIQ/+krCx+VQ36cSU2WR23+vCMm3oLrqHk9X6p4eL2muvPN1xjx10uOStCYxaf5uZCic0Qgn02aWyQcBmCsI25yIJmV312s7kzssKsLWzDx4bpnO7pucOE/5SBGyRcJh0o8+YeNMowca/eY8SBneNv6mcH9ULgBjnB5o260RauszgUVi82mZYP58zqwzZ2/G0bSPvO37Z5RMMaywnKwEICYgIhJnVAoEz+tAEi4qDrHbrTPfPTE27u/dQPF1IE6cZUH/KCWCCcA1/q/as8O2uU//QIYGUBCmU8C4QSOIj4gv6flva3XvBgWieUikYmP9oSmtcVE1iydXdGv+Nof01RQmv6PUkkdJfQtbeU9zLl6wUZL/J6YXnyXz9zVCEr8gU9gE5Uj8ejPBy4IFuQYLuGwFpugWp6Dm0XyEUXnjwKd1RuPYo4jpqK1z2lmAi3y9fQYGqyNWjVpbYvLX0V2ZVbqA2F2y9z7Ahc+6G5y9jFYXF3RqrT8ZyJYyEXXmsi/VbUP56kL/X72S481YugWFEniwggM/QIFQSdTDZNkeLuyvRmJQrcaXEYi/rO+G7zyUhh6BvrEdhKCIjMyEVaWJPo15AWKKowXkIasPZk/YeCDVYWrNn4DfKAdTSxJD6phBIKa03WjPeXYywuP1kr2rqTNTAWHJz/dFkOn8TPIKYba03Wk6wtSdSDudvWo3wOiQolf3gEPAIeAY+AR+CGIeAJixsGvS/YI+AR8AjcfAhI8P0pkRa/qZq/S2nSrT6+yyUiKJYfrrn27bGi+cnnuiScvSNrrrV/n0uR70fPuLi+V1+Gftg5oYQ1AJ9s3BBqsTFjk8QNCLtIbJgQ3DNX8RubOfPTbsK5qlUD3yEXcIPERs02gBAVFlPCYmEY+EYa8GnJXDtxjW0ssdDAWoQNI5pqXAuJYDE5qsJCs9owC4sqyVItz9rCZpFNqVmT0HYCIpO/uXphQ/uo3EDtcp3Hxt3q53ORFVwDrlyHVQgbVPLkPJtSPj/EM7PG+k+PwAYI0OfoZ33pc++Sa6ixtMgkMHVP50VwpwTmTTmEWpb1RUca/ieIDhoWwZKIirlBmp1J03R1MAgH/STdLG6JNvVDrtXCtNGIV4T1gtxoDQb9TJ6BiuWgiJ3wnZSm/WSSFPVeP20SoFsDxrT8BfWatVh/hEWt5jqyvjhdj8KeBpoeBJIE4LQ52ASuuBjL8Mn+tvIhHNCnuRTZ1M/lOlSOsZh57YSeKy7UAmLf5nnQUBjdlSTPt4uvCGoiNMRHBcSAyWPXEzF1TBZMi5AYer70zeGz3YiQepnJqOsAkc/SIzA6CKyzwDDFF5s3ByI0IDFwDUosILOaY3BHwYc1IIo9kMKshVk/s8ZlnDFLCFvDouiDwgrnGZO59qHyes4x3w/zV51G1QpudF4831KPgEfAI3ATI+AJi5v44fmqewQ8Ah6BG4GABOAfFGmBoP6rXJEcc4ufmHfTX9l03ef3u/qOmqspxEU6J7HaswPXuksuZPpTLti1TbqjFggb0/gnlRCws5lCUwwiA03hQ0pok3EeSwM2ZOc3V/puZEDVlZMFuWbjxrUIebAyYMNmRAnX85u5lDJNsiqEbBzNXRXXcrCpYwNJGdSNjSPXQSpAYnCwibSA4eaehU2g+fqturVaHxiXepE/hAPECnWnLDae5h6Ka55w6Urd9Z5puw//hyAAACAASURBVPmPFu7pnzRCAxxxvUVsCwJq40qKzSq/f4xnVdbRf3gEXoBAaWmRy9JiqFEpje+BNLuxrHBZFmSKnaA/g1yS1rZ+U6Btd1LncrmMWpSAdSnPspMiMk6LrOh664pLe8GkSZ+KYEj6g3RNhMVJCa13SgM/DuPwZFBEjD/jYVQs6/dEAbibcRRnGoWSQUqciywZb9bWIrEaaZEnGmF68gjFPRb75tIqcf2uYrx+ayV7xl8EZaN60J8UpyIiSP129aXniUEix2qhrC9iEX512S0NArFVsrwQr5GfjKK4H0YKuu6KFTxFlXPBqOLn2+0RGBkESkJj/RqR9rMmtIO1Jevjix4iPvidNeF5RRrlXei8kRTecmJk3irfUI+AR8AjcHMj4AmLm/v5+dp7BDwCHoEbgoAE4e8TaYHw/jvd2Q/c67Z//a2usW/K5b3ELX4sd63bmy6M6yIrOrK2mHRRW5snyeSjGi6NsAhAkIUVBMJ2tMogMzBNx6URwnoEcGaSjsCfvy2IN+QGZvP8zm+micZ3fjugRJwNSAcEaGbFwXWUxTkjJuxecKy6i2KDyP1s/PAffEgJzTRM6s0ahLZQDnlQBmVbDA3zBUy+kBkcbBJJ5hqK9ljMDsrju7lQGbrpUYLMeMSlq6dd/7lXuZPvqbnDv4j23bcpQUzgt5j6QM58uxJ1flTpD/SMcCHgD4/ASyJQBuLmOsVzztGIJ37FkggKvWty+zTIxogArDcdUiOSRjhxFTpKshLIIdb8cYkIrKz1i3otHpKR8uj0rIaDPY74BUGwJldQIi3zcZEQifwENWr1EJdBxA2Rd6iiX4vimmIj6FoXKKZIItOMTPfZWIUbohfU4mXWwme8/JdKP1FWBOLYLOkuEaEtddmQcGjUo1UFrX9S1kpLena3iLhoa3CvaZJIijDvxHHckqsveKiT6mXLIrQWdI0FueWz2ATWM1vqwfjGeAS2KgKQE2XbLiAmKue3atN9uzwCHgGPgEdgiyFQFdRssab55ngEPAIeAY/A9UZApMU3qIz9St/h7vrlW0VUyPd6reGiRuGSucw19sYuaKUSdOYu3r3smrsRyGPlgAukO5Tw04t7KBPQI2xH+P8GhDRKWB0gheM7lhdcjyUG90IEQAxAQkAWMKdxLecR8iDI4zwHRALnIQXM5RMEB+ckNBxaZFgQbYRuRm5wL3XD5y95YlUBUWBWE9QHAgafwzItGbqeMl/CZupfJUJMe84CaUP68B3CgTZaftSdeuFn+JQ7+2exO/WfZt2J30GYDA7UgfqCJaSGkTx/pO+HvWUFj80fV4qALC6GweklFG/IAqAh4qImgWtNsnPJUYOBtMMHshRIkjSjP6UWE+NKyxu1+973qSO15ZXejOiH26RV/1qRPndEilcgy5UpEUazsmiZ6PWSutihloTX9O2e4les1Ru1w3LP9ejEWPPgxHjjmM4tRlHI+MR4wXjwAs3Zl4uwKMkSxs2/pWRu6H5H3/+BUv/lqsdmeZdKF04Wo2loBSiCD4L5LvUhCPcJ9ameAnEfVqcak3eocQW8P67nzbWQ0MxDzG3MAaknLDbLk/X18Ah4BDwCHgGPgEfAI+AReDkQMC3Pl6MsX4ZHwCPgEfAIbD0ECG6NkOov3cEffcglp4+7vNt12cqiyArRFL2mC/LQ9Y5FLj3TcoNlC7iNSyUEMx9XsrgSkA3Eh0DgdVDpCxWhDUQBwlGENyak537KhpSw4KQQEGZBwafFweAetJrJA6E/5SIMelgJooFrTROYsiBWjOygzgQ6xBqE45FKXkZu8Ju5ZjEzfPKsBvE2/8KUY9YTxNzgO3WjrriGgrQg4av4hDv+myvuse9fFVlB26gLBBEkxbHyk+vA5S+VKJtn4g+PwBUjIAKC/pQMkqybpvmKBKu4lzgjgesc3xVfYUVkBf3HkxVXgPK3vvnWZLWbzK+u9Z9Th/1Ms157WtnMdfvJsV4/OSImaE4WFcvC+kS7ER8db9U7jVq8IIuMx5uNukiKYFlWGAORFfR3xh0jSa+gNtf8FqzO7LAx75oXstkzLAmGYT8qx2XFIAkWlR6XlQWuoY7IWuaI3EWdFEG1yjPV4+R65gebtyDGvfuWzf6wff08Ah4Bj4BHwCPgEfAIeASuOQKesLjmkPoMPQIeAY/A6CAgTX4E5+9RwnKg4x77B59w/WMrrnNEAvRixUUzfXmUabr6zszlibx1HxNpceoOl6cI8hH2v0MJ10pYTRBU8GNKHygFNrv0SQBXiAO0iCkDl0wQG5xDEMQ5XEmZi0PyRcDDJ8J/iAqSuYc6XX7HeuEPynuZC41k4HtVQARBAJlAedTn1UoElEVDlr9fqYSFhQVB1NfzLqqGcQE4UZ4zUoVz/IZVBRiQN2XSLoiKYaBWYdR0x3/tDe7g/3KXG5zgOqw8KBOcICnID4EWiTqS53vKZ1IWe/Uf8r0+tMbkUyksE98tca76t11Xvd6uIZ8L0tXX0OdwnRDgneQdgxi094z3kL+HGv3esuLKkd821cq3z7SXFGT5pIwoPjcz0Tw01qot1Gq1k81m7fPT482js9Pt+Znp9lPNRvy4Ylw8XY/j42Nj8ZHxdmNRVAXPgj5v8XJuqGC7tKCgDrj6swMypUraXjlgN+GdJWlhbgAZR3lmzJnPKWFdNycCIxdRMdCnArEHzA2Qg1wDCU2/28in/U2Ihq+yR8Aj4BHwCHgEPAIeAY+AR+DSEfAuoS4dK3+lR8Aj4BHYMgggdLbGSEhy1QIRuYZCsP9TSjUXT7/K7fuB1E1/xS4Xjr9SwaJTN/7qcbf25PMuSCPXvDOUV+/UxXtrrj5uVgmnhvd+MXgsgnusDxCM4m4JUgALAwQ4XEf9ISqwjjB3T8xpnIecMHdJ55upLxZDAoEQxAXEALE0IDsgDSA4qgfXkzeCI/LlOsqnPtwLwUAdOW8BuA3X6vxqAb7XCxQhaagnVh9oq3MQn+KMG5y+w81/aM49+t9/Tn/jrgocIGtM+Ed8CkiSO5WeUqLN/1RkBXldk6MkKozMMSuYqvDRCBgjeap+k88He1RlOG/vmJ23a9evQ+wZ0Ybhb3o/b6gg9pqA6TPxCGyAwG986IlovF2viYCYikK3T/Et9vXSfKxZi7qyrrhVmvfb9ftZ9YFev5es1GrRE1OTzcUmEZvjkPGHcYO+lUg4Tn+8oUfpFooxkTHTjnv05clRcwlljS9dQzGWkcxFFGM38whEM2O3ETt8Z24xl4Y8Wx+/4oa+1b5wj4BHwCPgEfAIeAQ8Ah6BG4GAD7p9I1D3ZXoEPAIegRuEQIWoYPwfCtd1bqjxfzXERSko/8ciLt7l0sXCHf6XUy6Z3+5mvmbg6rvaLl2T4KXouSyZdf0jkattl6soCd+TbQMXTp90UWxxJyATTKsbqwqEPGiiIiiHFEHgg6AOgmDoZ18JbVSzuOB6c8VkgvKhD3glIzKM4OA6yrVYGCZUNwE8f5M/wiWLGYFlBec5R3wNcxtlcTGGkG7weO2caUQbUUMsD87hAity2ernFavije7M++tu7gOU8SYl6sPv1NOCj9+l7xAenL9f+H9ogzKv6FT5jhhRQR3ACexI5nLLrFYow9pkZAMCN74brpA8tt6wZ0I7TIjHOfI2V1l85+B3hVA4D+dQeLe+UXpvr6id/iaPwI1G4AfedU/23o8/W6RZNr/aSfv9QaYxr2hL5b4v91vLgSsm+v1srtGIgnar1pflxZlWo1ZII3/YN5QYy0ibjdTDXZ25hmIcGNmjYmXhRF7Y+GdWSjxHvhshbtZ3dp0nK0b2zfEN9wh4BDwCHgGPgEfAIzDaCHjCYrSfv2+9R8AjMCIIVITQCEYQvpM40NBFaJLpGgRgV0tcfEikBa6OXuOO/8enXG3nNtfcn7vmrWdd68Aul/fHXfe5OVffHbrBosqrrbqop0Ck27suaprQH4E31g4IrhHI8506YoXBvAVpAGGBJi8WBY8pUSYEhwXENiKB9iIEQsBOHuSNMA1rBQTp5P+qyu8m/TZf4uRplheWF79RfpUQsftMaF+1MNClpcusEmv9jWYtsTTMtdMZ13lizJ394De5Z372/S5beot+g5Ag1gduoGjX3yh9qRK4UC+ImkeuFVlReUeoL+VyQCLQVhJkkpFBaAdTJ+oAjkZw8Ax5Lpw3V1lgbi6F+B2iB0yHAZvLfGiPxRHhu/lurwYsN1/wVYsN6rjZhLUldP7DI/DSCHzXV9w+HHcViHtttdM/XrignmVJLKZuudWIFfA8HwRBJEuMRi63QV2RFUOLCkubMBgz9fuI0veWrX+NPrEUu2pLvpdGc3NfoWeVl1YojFmMfzZP8GlE7XAO2YTPdXOD62vnEfAIeAQ8Ah4Bj4BHwCOwpRDwhMWWepy+MR4Bj4BH4EURQOhsgnwE+BwITRAeI0waWiFgcXE11hbK4/eVvkXpVe7wP4/d3u9/jYumsB445fqKxRDUx119W92lHZUn2Uw0EbmwW7janoaL25LXhWjfmy/vL9d35irOIQDH2gKSBWE+JAXC7zvKttAm2oOQm7YgRK8GMTXXTwjQIC0IlI12K/lZwG2ERZTFvUaAmKCNT/IwTX9zT7VeYF51C2UkDGWYVQHXU7+/Uuq4Il9yc+/b5Q7/i8gtPch1r1DiOeHuyixIwMNieYDBM0qPK72/bPu1+jCswRWigfIhTLYp7VEifgZkC22hnpzDvRZ1I0Fq8DvkA/eBP667wJnr7dni5goB3bNKlEU+XGeWGTxH/gY/CCrqZe6uyMvil2CBUXVJ5S0wBI4/bj4ECMT9C7/76ezWPVP9Rj2O0iwPGo2amxpvFJnMLZZWe8WeHRP0p/Nu0zapUJtxEdd2dhDnZ+SPkqgAhypxU3Wjx2/nx6/K9UPsRtWl1si/OC8TAP0fHBZka5eqa8bhD41ff5kq4ovxCHgEPAIeAY+AR8AjUCLgCQv/KngEPAIegS2CQMV1TrVFpqFuPrMR/iL4ReBrAnCuRyseYRjn46shLaTxn8vK4sNlfnvd8f/wOXfit9ruwP8567Z9bdsV6RkXNne6wZHU1eUaKjmRuKwjQf0TZ2WN0XKN22uKcbHoohquRNDUN+sJq98BnTO3TNYWcwVFWyywKVYAZvkAWcO14MCmHLdS5PFJpb9V3kM54MXv+GDnuwnJuR6hPXlTLzb05LU+5gJ/I7DjXnOlRB58J0/KhAhRcPKjD7uVh3a7R783dOkS+XIPAn2rB3E8iE9hsT0gljgHIfCI0kfBWp/X6qDdlMG7wLth7STQOBYX/G4ECtfwtwX8JnA6vuohgzj/50rEByEf1hrc92VKO5TAnOciy5rh86XtfDcLGnveZpkBsURdCOZrxBLXkgd581l1paI/ryku5OcPj8B1RaAUUA+tLZRM297KrPo921CovYkE2ozTuLqrHoxr9PORPTZ4Pt4ybGTfhs3TcBEVVQUL1kn0X+ZTI0c3T2V9TTwCHgGPgEfAI+ARGCkEPGExUo/bN9Yj4BEYIQTWB/lE6M1mFCG7xXBgDkBAjcY6gmV+x00RQmgsLXpXamkhQXqnJC0Qzr/ZFVnLPfcL2+UOKnFT993j8qW+C5qBSxaOuv7JW4YuorpPBiIqVlzeG5PVRUukRte1bsOSAkHXc0qvVaLO5j4Iwb3FsjD3QubyinZBEGClwMYbIaBZTvAavL7EYb8+KQN3SxAcCMsRFiJIJw+0/xEs8YkLpKobD/LhN4ToZnVB+WCMcP2zSm9Vov7UxVwdPeAe/saDcv8E5tSJ+uHvnfaQF26qsEag7uSFNYi5r6L8Tyl9Qhhz7pocpZUCpABtBmPqQpuMPHha37GKAAcSdTqgZKQChAP3QmxwnveId+7NZTI3XuDzGaUnyzZBAlEewcMpH/dc4IGGNvdjZcFhAYUpw2KccL0FHrb1jAl8zcc/93rBYAmi/9i8CLwE4XAzvcP0QSyx7DiqLyYU3bwPwNfMIzAiCIiksPUh6wvmYPonc7a5KLP5lLWiPzwCHgGPgEfAI+AR8AjcEAQ8YXFDYPeFegQ8Ah6B64oAm06LKWCBqc3qgIIRMpt7I4TPbFRxM4TAntgOCOu5hs0qZMYVHaVA/WMiLrAG+DGlljv5eyfdgpTv93z/Njf15Xe5sDXr4vGGixqha7yicIO5Wbd2sO4mvrQQeXHSLX/mgBu/d9k1b7/ThfW63EW9V/m8W8lcEEFYQDBYfAXqagG4EbYj4IdoQOBnWsomzDYhGpt2BOaHlHC1hAsTtPpN0xAhPPlQFgQDRAHfq0GjwRN3TgjZEbbjJok88eWeujxbc0W35TpP73WnfucNIisgMLA4gARAKA/BgeCAfCEv+MTlE20xEoayf0W48qyu9WFulSBVwI2yaA/EBIl6vE7ptrJgLBy4lusgkmgL14M17bhXCVKCd+tRJZ7RlygZKcQzxMWXWXXQfvJ+pxJYo6GNtQY4gCfEBOepG0QOzwlBKO/WgTJ/3lvyg2zhGQ0D21psFn13IuA2reC3dMlBNdcf1fgo9ttG54ZNVLI2Vt174NJj07Z9o0b7czc1AowZdjCnMC7QL6/bUQphbb6jHMZiDsYCG6vNIovzZpXFOM/v3Gvxccwy0cho0zZff915F13eZc51e7Q+42uEQGlNwbxAwtoRV4zM7bz3KAMw15oby2tpvXmNWuCz8Qh4BDwCHgGPgEdglBCompiPUrt9Wz0CHgGPwJZDoOISylz3IGxB2I4mOuf4xJUPQmYEShYHAmE/Qh2sDdjEIixGoD5093OlVhZVgEVaEM/gK5TQuIcMKNzEvbe5HX+36ep7ZyVJHrh4eocsLk659l0NuYiShUU7lhipcEsf77jJL++75h0K0N1cc429CMYhFZjDzAIAwTakDBtvvrPZRjjOtbYhN9LCApzSPn6DnEH4jrslcCIfSAxcGiHgAkNzP8R13GPxKxDEcw/Cccr8f5XAj6DZb1T6gusf3+86T5528x8VOTS41R3/rcNucJr7eD4ICCCNIC6I50BZ9lwQ4lMu9cKq4uMiKyAKrvmhd4d28n7QNggTDsoFM3CEPEDwaHFA/lTfafM7lMDrbUpYYfBu0QYEeRALPAvIG347UObHeQgNyoJ0wPqC4OOUh6UGz4y4JBAQkB9YZPCOgovdBx7gBXEBzufcbJ0jQXg2kEDkwzPh+ZqFBkHlN6XgfgPCgvfKLKPMHZpODQ/aAM68R7yrPAveJzClzbw3CKAQyoKrHfbe8bu9s9U8+b6hoMoLZCso+q8vioDcW/EePqgEmfmQ0jfKgoRx4IqPDfqHEfOWJ6QIYxXjGGMS4wp9COs8+ghjE+//ASXmOurFuMF13Mu4RJ9gvDBLLvof45ARMMyfNo/QHr5DpPKZqY/kJXEyJID5+4ob7G/0CFwGAi9CeJOLrV94zzl4v7Hi5G+LJcU1KAZwMN/Yemp4wo//l/Ew/KUeAY+AR8Aj4BHwCFwTBLyFxTWB0WfiEfAIeAQ2FQKM7aYxjxAToTGCFzahfCIURkiDpj6/WfDpqjYpgk7zO37VQhcE7aWLKKwGvkvpVrfy6JIbLP6FG3vt14uECFz7jgUXxArGPT8rgb4EQFlX8Szq+r0p91Cxy0Vi9J7LXLo85er76jpXKM4FsRMQUEGwsOGmjeaHGcG1bdDtAQ0FS0om3OUahFm0EYsI8gAjBOnm7gkBFufYwCOw4pPrwMjKZNP/ASVcTc26LHmNyxcjucA6oMsmRFpELplP3cn3HHPZIvXlGUFUQA5AQlB/hHyU85gSxA7lQ35gVfK8MDRhgv685gftBxPqZq6rOEf9IFNoH3W8Swl8wQoiAa1pC45NLBC+k7C44P0BW4SWEGEI2DmwpOCdg5Dh/IEyX8pFkAIeEFwcXEOZ/z97dwJlWXaVB/q+IYacM2tSTZJSEkiAJJCEhAEJkAAxiElgN6Mx2BiWod3QxsbLdttN22YtPDTgqW0M2AgbMAIzGowFQpQAMYMEEiA0QJaEqlSVWVlZOcT0pt7fq7eLV1ERGZGZEZEvMvdZsdeb7rv3nP8MN97/n723fkQw8vIgZsDe9z4vDI7/a3K8Y5GOyETXN9aJQs6NWGxPhL09Fy62QShpQuZQ0ffanInNjRd9wDK0m3BjjjFu3hZGmBBSC0Hr+y+Z4AQbgg+RjwhH+HEeuBCKjG9YwRF2Pk8SNkOdqdtMCj0qVmXmEDC+fj/M3DfXL4aI4Z40vpdsFP5qk/mRG6s8Tt+HzAdrC5Ehw+1Zq8wXa7B5wLPrDWHEY+tqeolZz8wHa5TjFSEBPXdOOXYIo9YZa9mvhOX1PJpnrw4jYjjXW8LGcyPakKKMte5MvHbsdKL0aQ+oyaUffyhC+Elw1IudQyA3GZiH5qD/eaz15qj/AV8U5j7u3uv/DUJ/5u7auVrUmQqBQqAQKAQKgUKgELhCBEqwuELA6vBCoBAoBGYNgQkBm7tN/SBFuiCekY/p8u99O0UVP1IzKTTyczocELISuZP3Bwm4kbs7IVog3P8ghItvj8dPD/vsZvUDdzTD5d9tlg4/p3nsLe9uhuGBsHD3oHnaFx1q+uciLNQhnhfdZhRNefhHLzZHX3Jbc+n3LzSX3nap6d75cHP0BUFMLc5FPoz7m043SSntg4Ef3tqfJHC2SXvHycXDELXIJo8ZTsRrRBQiF8nlfaGN1B9BDIsk1/3Ad54zoa/0muX33tN0Dj6/6Z1+uBkOjzer7+s1o958hLZajFBYD4ZYoY65Ax4Z5ny+z1MAoUDQQZzpq58Ne0MIFdlv8XJ3iv6NfoaJNhs7PBu8TvEgdyvDCUF4KiwThPO8QHioPzGCCJGYGZfIQeeFKSHCuRXfy0IgIgQRQlKs8Jn+Y4rk31k+JZ7AMsMe6Y8MUaXvEfgpuCA1T4VJYK5N6tQyb2bA2yLnbY5R2CNKM0wNgSHDcznmr4VJbo5k0vYMeWasI1qRtT8RZgf5p4bxOjEfjN3XhBlrvxeW3kffH89hnrle4OR6xlyGQnONQZCvsEN2mR9PES+KcA1UqiQCxqqQcIr14FiIFFcSEiqF41yz00PKeXPdMW7NF0Km8Uwc+ewwwoW14tPCzCUiJ+8+HlnWBOuMMf2yqe76gqnnr4rn5k+WL596vtFT4ukvTOryk/FoLro+Md1cnF7nrVFwUIds0xanr48LgStGYHyPm5hNFu4XBGv/77mXW9uNQ2PU+z4nwBmf/gfMdf6KL1xfKAQKgUKgECgECoFCYKcQKMFip5Cs8xQChUAhcP0QyB+mCFyWhA5C0w/T3B2KfCdiIN+Rxn6U2mXth6vQSn7MZkgMBLPv93dCrJiGBgEfogUix/lvDc8Dpi5I60PhRfFYiBfIUWRtLwSMkB/uvLvp3naxGa2uRLioY82RF/Wb1bfd1gwvvDc8MD4sclvcEQE5DjXtY6ebbiTrfhwHZJYf4fCBCVIrvU8yXjniFXlEOMjdr4mnYx2XXhuEBMcjqDzCKESJB3+5WTn1ceH5cbAZXorzjN7fzN8VicUvXmwGF6OOy2ebMz8bYsa7EPR23CY5jchST+dD7iG6vKd/2E/sZGLtON9WRd8bL8z4sPseoQEHAgEiEFYZSsj7iHA4ZH4P/eY7dlcjBI05ycd93xizi3OjAgMEpJIeANPCxfrvECWmi5BVxovzEEiMJXXJsBbPi+d2PxNbYG68DUK0GO30+N6kfd6e3i2er2ECa58hSZNcUk+iAUw+JwzmPpsmUp0jPYjg/MmTa3/VVB14YbDpgtTN8o2TJ4QNIo/rOOebw3i36C9zKPMBENYy2Xtiay5cs6C5ro71cp8iEJ4Uam7u8XAgEhAqXxHv/6hxcpnk4u4H1sYUkoV3S48i50gx1NwgRHzG5D1rz2blf5/6wDmyWF83K+vn2FY9ob4EeMU6Y/00h+Qvsg7xeLL2a5/Xikf3XvNm2otpq2vV54XAdhAw1nhRmEMECvcZ90fihP8xiHjuoe6V1vd3Tcape7f/B2s93w7KdUwhUAgUAoVAIVAI7CoC+eN5Vy9SJy8ECoFCoBDYPQSCc/Xj1HqOoPfjFOloV6sfnYh6hLKCsPcjFmmeIYiQ5D5HqPhR6zkyxQ9Z31/bbUI3xAu7+5BECG7192NaPU6GIc2RVn54I36QQ0ghZKrnyO2jzdGPOdTc+SX3Ngees9QsPPOx5sDJs+Gd8bSm3UG4Iqr9OBceKEUcxFgKFM6jrYQJGOZzxCwCPD1O0jNiuRn040f/aK5ZeffpiFp+d9N7JPJuXIjj5zvNfFS1/1gncnC0mtM/udacfcNbm0t/hMVDuCGhnY/4cSoMuYXc1x+/FXZ/iBSI4z0vk3GkPvoADuoMX3gbN0IMGSfw+vkwWL52ciyCjidE7tBMbwvvC3GlvYhFY2y6yIUBZ32vfxReJvqCCLG+GK/OZzzkeJ4+hheFMc/zBQmP8Fcn5b4wuTS8RtqkV8auhYeaxLPP3eLpEWIcER9OhsFU+BnjLBO583YQEswcTg+S6TbykND+KyVWp89xpc/tYv+lsF8PI1Agv2CJkEZy6Zex50XF7b9SaG+s4yeChXFLKPvpMOvJ14R9T4gVT/LMmcr3YE1JgtX4T1EMqf8VYZ8Yxmthp8a8+baXm7Z4qpkj/y3MPck69fbJe+YRktiatylRXB5MN9Y82enWTOaS0/pfhwju/yj3EP9LCYv2dyfXzBCO98Vr49L/G+7n5gRvPI9PKjX2drq36nyFQCFQCBQChUAhsB0E9vKf9e3Up44pBAqBQqAQ2ASBqaTa00ek8IykTcGCh8Hju/8fJ4GRzhlux49ZxHLu5Hcuu7MRQX6sOi7j2TuPUEE77mXxpAY8TtC/LYSLzLUhrI0d3rnTVr0QvELhaNc7w9JDBMEz15z/zfdEOKYDzS2vXmmOfczRZuWZ3WbxmavNwjMuNN1bHg3hwg/3FAvg4TXsXNN1gxJm1wAAIABJREFUkMm5az93vGaoLOIGLM5FmKejkUvjTLP8J2ebueOxy7d/NMI8rTWj/lwzf8dK0zvfCXHiTPPIGy40o2G3Of3jQUaNkPcI3sfP8binAlFIG+2eF8qnF0KFcCLXrUzCQiHV0ruFwEJggJPxYsc0MsP7MEMgEiRyR7Hv+T68EHL6jeig3emBQSyDhwILpJ3zGKee62fx57MYj9M7qNMDyFhHcK4v6qMvEZz6005s9VcvxKnQLeLVe8+4RxRuGOJog3Nv+60p8ghO8DGnPJ4MM9dcUwx9u76FqyFYSSSemF/Ou8T82OsisTnLYiww8fsJQ8YHgUvoKFhLQFw5L/a6l2bgejwoJqIFMtScU1JUz1wP016B5kZ6FllfzFtzXogn68/XbrNZxiARczvlan//EMrdV9fnRtrqmjmf/6+pA9X3O8OItoRg6x+BZhyCbasT1uc3JwKXyfViTJtH/jcy79zbjKuvDyMCZjFHjDVerjw78/8sXkdPEStuTpSr1YVAIVAIFAKFQCEwCwhc7T/ss1D3qkMhUAgUAjc7AkifzEWBDEVycO9HDjE7yB2DIEbS25mOVOTRgHBBDOVxiOQMl4RIQSL5rvf25EdsEPavD9HC9XhEILrfEZYJtNUFmYPQTS+S3I2KvH5ReDn8UfPQDx0Ne6w5/MJhc+/X396M3rLYHP6oo0339nbTOfC+sHYzfyeimgeJH/Fw8CMfFgj0FH6SUOs1a2ffFd4az21Gj3WblQ+eaUbnDzTdW082F956seksHmjaB6LOo0ebi394OBKBD8PTot+ce8u5Zu1BuKmr9hAlkAeuqw8yhvm3xPM3Rdv3BOO41lYFpuriUV8gP4wjJAeyMb0AcuzxZLCTE+HOMtkuMeHzw4xJu/Dhy2uAxwwPASFUEH88NJJkRFCuL8YnUoWXh+K8BLdpUWP6O4QPhJ95oNjNrM7pWYTEMdZTsDAviHLta/UkmhIpnNs40vfGVnqtEKpeFUakOBVGxHJM5g4xLqbzdKh/5kqZbuMsPOcVwr4wzLryj8KQYAhmgsXDgYf5tFbCxSx0157Xwdrh3pSFgPifw4YxLszpvP+kqGUOEKKNH2HKvugqarxdsWKjUwtb535g7pqXynovDB5+7j87VdT3H4YJ4Wa9+KGwfxNmzXCvI85n+L0S/3YK9RvvPOYTkd7/eeaP+7D7Ha9F/19sVKzRvB6NM8f7H+UpibbLs+LGGyzVokKgECgECoFCYD8hUILFfuqtqmshUAgUAn+OwHS8bwQ8AsgPT0Q4shlBjOTwQxQB47kd0emRgYxBhiBRkaZ2w/qR6zwenQOBuushoaY7dULc/1wIF78d758M0zb1QeJkomVfcf9ChL84zA9tO/oRPH60j5qLb+807/zqEAe6tza3fPJ7mls/7emRT+LuZuHeTrN471qz9J53NXd8fq9pH3la5KB4KHJkPDdyTqyFMBEkWye8H9oLzdoDK/FwvOk/+pzIT7EaCcGX4nW3WXrnQrP4Ie2m1UWGt5vhoBWeF8vN2iOnm/NvmWvO/LRwJhm7He7IBH3whgmmRAuEwaloL8J8ZsrEy8LYEOYnc22oa+ZGEa7J2DN2CAknwwgARC79hDAhiBGciAeOgxORgreD94gcWQgLmYR7Ggehhz42DJGXYkV+brwKn8XjhhiwvhjDxjXLwgvgl8OIJJ8UZp6oh3aq45aE4PqdrUnmTISK6QTgBDRkEM8J/W7sPjcMsY+kJEoQcjJkhzoSMTJE1XSeDzkj1A/5ZHd3JkZF8MKbKHBq8n1j6UfCtF98f94Prw4zV8zvzw3TP8bn+hwg6nC1RXvkJ0COIcCE4YIrwfHBwIc3UcZF39Sb5WYnxyZeCfog1+gn9cf6cEpX21l7+D3zIMvdc+cf6MZYMO7NWeNdmBpznyeW0GiSwmdYuMtVc73X1fSxPxsv0lvOGuy+YOxby8w3c0FuCa/z/ncqnrs3mq/WLnUyTn8wzFpDpDCG9ctnhplnvKQyRxKPJ9+72kKAVeTbcA+3dvyvMHVPT0jzZ1ZE7attZ33vGhDYwLMiN1Wk9557jbFvDP3zMP8bbVSszfeF+Z454L6yVMLyNXROfbUQKAQKgUKgECgEdgWBDX8U7cqV6qSFQCFQCBQC14TAVEio3N3uB2eKE4h6P1S9zkSLyEzEi52jiBq7/D23kx35IdGiUBWOR6L7sYsYQZzmjrtdDQe1XUBCwECSI0aR2Ihq5DeBQv2RsMgpuSA+bdIGhFSSpNp8tml1nhPeFYtNu/to0zkeeLQvNJ2D0dbhiRAq2s2tn3JLc/GPLzQLJ5aa27/4uc3qn43CS2KtufD2VjN/W7tZfPqFpvfoXHPg3vC6ONeP7x5oFu7oNud+eal54D//ULN2Rr0QcUIrIMkQcwhnO4cR8H8YAsW+SGY5yWeBaIcjglDbkI2IO+QiktE4ORn28jBeDIg+ZJv3jT1ht5wDuY6ER/45HqGeuRkIUy8Nu5qif6dJ0cudw7G/Mrnum+LRjmrzxaP6bZl8ex1hlOHCzBnCAVLT+cwj7TEfeZgQKBCcSR4ZD4haWG62acTYEfvfMchV89QOdcIc/AktCFMJVBFOBCNjDuawz5AgPB70izlCvEnhj3Bi7uRrdf2sMG1CZlkfeE9cqahBRHKODB1FPCFwIcS0I/HZkHgtwWKcrDpJyBTQcp5MrxsbimuXSWbtvHtWQnjJNhh3/2/Ylzaj0Z+c+N3XfcZdP/0Nxh1PK+MN0U+I2yhPy1b1JUwYt+aVefL9Ya8Ls17lOiQ3hLkCL+PaXLUOmaMeM0xT3u+8Z8ynaG+euMeeDDNmU2xzHvccx2orby9rnTo5x1eGEWgJhNZDdbrSuRRfGQus5r4QdtYu7bEGbNj/N/v8AdiNXNbdf4w745Dx3HSvsUkgPRAvFzaQuHzfZFzZdGBdrhB+N/LgqbYVAoVAIVAIFAL7FIHysNinHVfVLgQKgUIgEED0IFKQGAhkP14RpIhMOzMRN54jZO18djxixU68TJKL7PR9n9l57XvOicS5GiJpVzpmQvS/I4QLpA2yliFViRhIXIQegSB3jyNJkbQIbe17RjMaDJrVDyDMAqf7EUjaiZBC6p5uHn2jH+6Pizvn33YmEngfbQ69cK45/LxRs/L+fuSmWGxGvYvhkbHYrH1wuXn0Te9oemfgnXHXfR9RpS7ILrt2EWYSaSP9902ZymeR8a2NITgRtzzPBNuIemIAkt2OYJ8hyuH/yWGZsBtJ+HNhBAwEC9zsxE+xAtln9/KVlO2IFchMhKFjXe+Xwk6FGffGh3qo/1KINOr+lNjxgcV0nZKMNX6MN98xhpD05iCCHuFpnMILPr5DrPGal41kxHA114SZgRcPDJj+lzC5LOBpPJmnMBMuJslK442nBQFSfTPmfdYNOas4znvER/WCQeZjIXT43Gv1Qo46FhmqHur1qslnxvCXhwnfdbmSO9HzmP9t8kQ77B43Pqw/2u092O0LAW+Ldu/Ux/DPUEr6Icdurs2uk300mlWPi0m9Rr/33gfWhnOHWo3502o9+/B732iOGGvG+l+ZPL9S7IjShDnCnznmvmYMvz6MMEyEMM4IodYc97Es6XEIQ+fIsHE+z9CIMGde51pgXivGavaJe63rMmJcrpPmgMTa900etZkA6H3znipl/ZsOlzVVxSc95fFxKszaYS5ap6yrOXe39Arb7MT1/r5FIDerGH+8kU6G8e75vDBC4GbF/0X/cTIOzZ3fCfO/ipB95bmzb4dDVbwQKAQKgUKgELixESjB4sbu32pdIVAI3FgIJCGpVbmzOxMaI34RGAiRTHCMeETgZKgZxCryMT0wHOc1IgQpgsx/YgdnELUIxZkqE+LfrkAmdBTS+FPDhMAR8iN30mbeAq+RRdqmjRnmyGsFAQVLJHMShoPm0V+8FBbtb8f5h0lUIVldz7WJPs6FQIKTayPPJFB9Y9Qzzz9T+F1JZfR/kPiZ00LuCeMndwoba5nvA6mO1COQZWJzZBt8kCOIFTuF3xxmB/IrwzInBnLxxycYGqu8N3ayTBODSBv1tOuZCED08n9QegEYC9q7GRHoWO1H/BsHCCJimTnn3M5LFDkZRnRwrO+YfzwgFIS9QjD51jCeQYqx6ft2U3sv5ywyCb6Z80TdjFPXS/J6fILL7LDWLiSnef6kMgnR4xow0Hbn1Feu88NhdpJ7TjBBACOb87o8a6aLPt0oj4C25Q54Qow5+fNhcHPODGO3vno32+skI7UbYZ6vjSPjWD+kZ89qeDLo15kULuSpePDtPzI891FfcnbUjbw+Ue/W2hKvOJ4VPIy2U3g/8VgjdJpnxopQSc5jvSayGTuER+KFtYcYBpcnhJ280BV6IEwLl+tj+5sv5t+TSrRZH7m+Oaxe5rj1BjlMuHhbmLnNYMIb8GvC0tNj/Sm9hteXhJkz6SXpGubROMn9Rl+q9/Y3ApcJ/+Te4x5ifMnzwsNI2MzLiRVEvu8I83/Oj4UR6tyPjOESjPf3UKnaFwKFQCFQCBQCNzQC/qGvUggUAoVAITDDCExCQU2TV4gLxCDhAYnus1eG2dXvhygiEaGTZKmdp4iuDB3jfcSwH7CIDwQMsoch35Gbq0FY75sdnCFc+CFvJ+vXTfDwGumbIXFSwNC+3JGu/doKQwS2ggRCsCLjHYuEgqVjk1yFGcIA+Y4EhtO/D3t7CBVPIYUn5923DzH+jC94MM9h6zkcebl4bYwh64lDxhnxAj4EHaS3MYfER3jbLexzIg/BjACEdDQOXzn5DF5eI1Rc62qLvtWfiD1iEgIU+YdUVL/vCzsVZuyPxYrp5NuTBMHmjvGjDertHOr22ZP3jDPjyBgiZBEenFNYjhQMjSOCTXrjwEKYMNdNocT1MyTbU5LtXiHhGqe6sjJFkk0Lo07iNawYcky/mydC3phzvLi28r6YrgwvE+GjELeIZgIJEvZyYtHlBJkra+h1OnoqR8X6GuT/4saZMbS41ou8OGOxsHWw3W51w4b94XAunhg/g8FwdDZepCg6DlU0Kx4XMY7Mk6ODg7c++/4v/6lvXbnzhQTl5p4f/5rm2NtDAxtroFsWIiYx05prbTFPhFazniBazUdCnnmijMWbiW148t2eP+svOslt4+2cT9ZJ4pM6p9DyBfH8H4eZV9spPJ/+aZj7/K9N8AHocK/bt53K1jHbR2ADkSK/bF3I/0GIde6xxro8FV5frtho8G1h5g3Pnv8R5p47zttUeSu23z91ZCFQCBQChUAhUAjsPQLlYbH3mNcVC4FCoBC4UgT8YE3i3M7u3N2eBGqGbkJ2IhMRi44XCsYxGRpJeB473v2IVXyGzLW7Osn43MF7pXW83sdrtx/lfpwTFxDFYjr7cW+HoRwM4jtnEnKEtfcytr9dsIqY6gggP+oRZYQdBLdQUUmeIaQRR5IKEy8IGwi19TtxrzcmO3J9wlWUDEOCfEO2Id6QhHYNE8+0P4lF2OkDu4qNNVgbjwhGBIvPhWxBesP2ZJhxaPf09K79y/2PYpeovtuquAZi3PHGudfqc1+YsaH/9OuTxLkJ2ajO6oBM1F71N4eY7yDZ4UJ8MC/Nuy8M8z1ihM+092fCkKxIetdPkcx4MXamPZkuS9rHsZct3/L9v5VrQetDn3nr6N33PzL6h3/5ZU+0bZJfoEFue74Jyb2e+NXnhB9191zfEpHgqC3a+rqwTw87GbZVaC/HMX2fnhcprsL4ZgxRYsws9PvDWwbD4dGlld6o1xtcarfbB7pz7U633TrWikQ7vfbwoW631Y+3BssrvWZurtMZDUe9eFxKj4vNBshu57iYeBjk2PiEVn/1zlZ/+QkPp/6hWCZGl9XACZdIeOu0Ndt6Ys7k2BsT82FOQiTMk40fZ42wnyKDx/ULfAhM6p0CFe8L3iMejXkC59/drP8m71uzeKhYb6x/wsJZex+O82eYxw1PMWv4bNHO+vjxTSbmj3uj0JfEfp4U7j1/KYxwvlXhJWd8WavNJfe71RIqtoKtPi8ECoFCoBAoBAqBWUCgBItZ6IWqQyFQCBQCgcBUUu1pPPxoZRm2CHmKtPE6BQe7Te1iFyMb4YN8RyYLF+Az5AZi0funJq+RxpnnAlniGkkG7RvPigQqPBvUWUgm1oTHBXzkRUB+TYsXfrzDRogR30H28FQRHkhBsHuP+PGmMCQa0kAYhmmRAmnQjevOXNisxGQnHyeiRYYMghuyHfFm7GT+FO8hRDLsVnrvGH8wdbz+yTBmPjc+UzAwno1RfQFXgpJ+JJCs34H8K/GeHAlJ0E83N/vUe8Ql5jqEhcwFwVNCDG+F4EJQyJ3P3ktinghhbqnHyTAeFMYU8YMIQsjyHvLIjnBhauxkReJrF6JIaBt1MuZcJ+PkP2mebUUohhgxqe5THuDGhgvz3fH/dccOLzSra/25E0cPDH/yN9+3cuzwYhMkeOuRc0vDW48fHNrtv16suMz1k3BNISOx4tGV3lvaBE8k6r8N+8ow4g2ClpAKp/UFbgjabwr7N2G/OjkfHDO/xba2428GzCy9v5lgoC9CfOgGl99dXu01vcHw2IWLq8farabTbrWb1X7/kYMLc3d3O+2DnW7nUHhWLHQ7g9ORGuKxGKWPtVutpfDIGM2HaGEMhO3K+r3JDvBp7xBzSvg39XhRiBVHD7/3Tf3lex+PVjM4EB/LZ/FU0ULeFvNbv78lLEOUEZef8DRaNz53pY17MF6mxUBzQ54jHmnuUTxIrJ1fGWbN2ax89eSDL47Hnwj7/8KQ2jyVrJWuccPMmz3ok1m8hPuN/0v0o3CfPHFOhaVwkaEFN6u7+6x7XYaASlGMJ85+nTuz2E9Vp0KgECgECoFCoBDYRQRKsNhFcOvUhUAhUAhcIwLIoBQshJNA6gi7g3y169SOTQQhcgPR4XMJGO26RJZ6jRRBFvrxa0czshEJi2z1w9WuaT+KM9HomFDZV+GgRqMUW5K81h6Ep9dnoy2IIAQzIQNOHxpCA6L1TfEaUfRYJsWO17A9Fq+R6Y5Hmr87Xm8UK/ymECvgoEzGBG+LJCkz1EmGwYItMcKjz+CDfEzSkXBh3CJjjEFkXcZjJyoQ0SSgNqaNXyGXjEdj1Xd831h+dZh+sztZ7pL1BXm3viBw0rOIhwTxAMF6cnJNc2NM8k28K/x/hBRyTQIFUwfn0S7EbAo4xhlCiLj1S5NzIluFbckQT3DIEFewuWLSKDwlNmhW04SQkblEloLkXoiOOjwcjeaDxA7Cu9V97MLK2ZXVwVrs3O9duLS6dv8D50YPnr5wxddfd/H8foovMEiCGT769s1hQkZZe8Tih+VGBR7fEGb3uH7gaZMJlXPX+LXWd5NLz8bb/eHo4HA4PHFxqXdnRIJ6+nA4uv3iau+uQcSBWusPVpfme/ccPDA3CIeK1XandSHEiRMhZvzJqBk+ePjAglwzC9G3yyFGadBmnjM73Vj9Zq4LY2XO2fkvL4M19Itaw0Fz4P10u8dL76hpnUvH+K1MVn1fPHcfMl/MIY85V3a6zrN2PmuI+5N7ufWJuAmPLwsjSGxVbFJwfK5tRHX3+MpPsBVys/n5tFcF7073xE8OE37vcrlOsjUpVFC3/e9nPSWIjf9/KbFiNju9alUIFAKFQCFQCBQCGyNQgkWNjEKgECgEZhOBJIOQpMLRIP2YdRspjBxEVGbuCcQRkpBIgSC2yxt7dSoMaSqOODEDIezczoMkSQbpifAa+1Cs0IOwyB/7KSSMCWieK5mXYCI8ECvGJYWJqdd2qLL8/Ilj872b/XFqfIzHTOCbSW5TnPB+ihee+zxFDGMRuWb8GddIFd9DUBu3hARjl4CBfDFGEd/CeyFFnYf4ZGzzZiA6fHhYkuEIO2KIR0nnnceYNzcQg65PfCCUnJx8z/VzZ/J0mBnjyfwiniDTiRJYV9cyLowvxKBzOac2GXs8D55IJL0BSXTN5Psk9FOKmdr7tE67Peh02upzdHmlf6jbbR8L4vvA8NLoT89fXH20Pxieu7i0lvNdPa+oHlt4gAxD6LEuMfXSP/eFWaf0v76SPPgVYZsVpJxiF/HrwwivxCoi1w0Zbk1YrlMfeHT+SLhQrPT6RyIM1NOa1uiW6Kujy8trdw6HTYhQrbnoz/A6GvUXF+Z77UHMl9HwxMEDi4e67W7kuGgeHo5a5xc63bwfrAkPtYs5LfLe5F7DG0roN6IFweITw8y7cWmv/XlKn/6xeynh0bzxRzzYzCvCsPnMzH92QyaSvsz8GYt+MX/MXesdzz4hsV4Xxuvkb4X9zcR03SMB919N3rOWCrWG5DYWMt/HFc3zTa5Tb+8AAlvkqfC/nnmU/cVD9lVhPNC2KsbNt0/mj34X+pNQ4Z43DrG3lQffVheozwuBQqAQKAQKgUKgENhrBEqw2GvE63qFQCFQCGyNQO5cR87arepR0kW7uj0ifBE7SAmkrh+ldloiZ3lg+LEqzA0yCdHqOLvznEeIGue/M8w9wGfONU5EvQ/FCuSoNsBFgRfiByGLCBonZQ1SfRhtuxlj409g2b2HwHUC8eP6xWR85c77HMteZxipJGTsntd3CPcU0Twaz0QAxEsm7ha/27i2A1moLwKGHCJCQ/3VMLuR9bVkva6FKSXw8ZIw5gkIxoQxb04YL4SMFD+Mm3FcfAJDEEvGSsabRwY53nsIdOIEASTzemgH8UXdl+P7exWOZRwGSruiC47GGJ+PkEHvneu0OkF0n4jXc73hYC4SNJ+ILM2PRoioJILHWIfo0ZvObxHvXVOZEmaQr7ATouZUWIaD+ul4LnSWUFCXK0hvRhTyHWGCfiPOaUzogw0J2N0m5DL/x6Sfs/5P9PXV5ogIz4jh+Ysr0WWtxd5a/97ow3tiwbot5tVtc3Ots9F3y+Ex04poUfOjpteZ67Sb4WC4OByuHj640H16iBvzBxa772932pfi+VqEjsok7jtNVOf9CKlKkHK/IYQjVd1f5Gt5UuleOh2ixaVmOH+oWbnjI5rh4vEHO0tneNDYAS7/DTHKvM7k2Ttd5y2G2t59fJmQbirR+pd/vnlg+Zvue5l7vPFu/TP+iXju/9bBzYpjfyGM0GfuwfdHwnis7NWatHeA7rMrbSBWpHic3rHuMX8hTC4T/9f9jTD/w21VzCf3RGJ/zidj57I5TbY6aX1eCBQChUAhUAgUAoXA9UagBIvr3QN1/UKgECgEnoyAH7HpKYDMRaQic5CtnjOEn53lfuja7Y0stRvPDr2MfSwUgM8Rh76bOQAc68csMtdOWM/Hu8H3oViRgos2wSUJWWR1JkqGHRwuBYGrnf30tqiBt7MITIQLJ50mHYWQ8p5xvZ400y/EJSS055lLJRNTEyyMdd9FXjuWYIAo1b/GurEt7kx6NNidjLhLbyQeEYg+RI7vOc7n5pZk3JnkeSNCj1BhXJmPdqu6njqoV87JscARr5eEktrDkBvqlP/DRVtavVa7dWi+2z4QoYVO9vrDZ0c8qIvhYXE6CO92rz+ALZI5w3SNw6gFiTrYSdEizjkuExzGYbACF+SbdUaOCv1DtCBIfF0ev8mjcGzM8dpq1znspxMub3GK7X8sl8RlSgpvuT5ba1KcuyaSPfqqFcm2u6v9Qac1DO+iteELR83oUCTTPhEeM7es9odrkfb+cISA6q+uDUb9zmAU3jRPu7TSW16a7y4dPbTQP3xwrhUeNRdDrLhqYvoyu7+12dh3z2HmHnHCnH1NmHvPhqWzfLY58Vvf3SydfIUcFuf6h25/fQgWyFW5atLDb20P5832B8QOHzkd0i3mXZLVGc7Q+M41sPmXr/yt4cef+u6V551+Y/+2S39ChOA14V7vmH8W9pGbVM969UkTk1OGkITQ/oNJUu7KYbDD/XoNpzOnjAP3I16FvI2si9+4zXNaV/91mDWRKEV8d3/juVSbM7YJYh1WCBQChUAhUAgUArOLQAkWs9s3VbNCoBC4+RBIUkzLkWDIjBQmMk6+YxA9CFghOOxeRsQiKvyA9SPY554jVX87DHmboXROxfPcpYx8Rf7ljtz9hrg2IZ7V3/2M1whcYEeMQfBon3Ymtnb5527e/dbefVnfdR4Y020wDvULEj0JPJ/rP5bx3e08FeLJe/oX8Z6hn4x7RE3mLME6i4PP08i4QAY53rWEd+K9QXxwnM/MFQSPMfEE8TwhUFeD5Mu6Zb6KrNtTQmzsNuk6RXLCKAUg7Ucgs9tX1vrWi48IAvz4aqQ/CMHiw2LXvTb6PBOiZxgrWCxPPC2umuhWmcsVHicTspQ4RLggPMhf8FNhyFeh6jYqhEd9J+GsHflIW94twuToyx2t8xYeEqOJh4X+39TLYyss1n/+M2/+4+bo4YVYu1oHR8PhYuSnCH1ptBgx7NYi1NNKuzWaixBKCyFcdBbmQ4KKNkd/RhKZ1tOiIqPecDjf64XfRW+41ukMb+s3rYvx/jAScw+ivqNrCAuV66W5Z23lsUf4453ktdwxnx+WeYM2bHpr2A+h4sSDa7d+6PFWb+nM8j0v+d2F039EfDQmx6H7dnveXGmf7OHx6bECB+M8c1O5hze/evKrl8KsYWfC48JcdR+Xr+o7wgh58E+PC2ua+990sVOf2aX/nWE8WYrM3sMO3uRSKXrqT95K+vsTwnjEyM+0nSLEHk+a5WGrc3HQmnvHB48+/+Gnn/sdgtSOrovbqUwdUwgUAoVAIVAIFAKFwG4gUILFbqBa5ywECoFC4OoRQGJkiAAko7j9SCEEK7Oz1Q9S6zcygzDhfWSH0BHi+SODEJfIfKFz7DL3He8JkWM3HuLCe2Oidj94HUx26ieyMOJZwRDP2pY//jNuc8bPn0543I3zlJdForiHj1MeGNNXTZEgPTHWf4a0Tu8J8yBDRhGe9Ls54HPzAQFkR7HnxgAikKeRz31GwBIqxXl4ahgXeX7nGYsA68YZz6Os0zXtpN8RLnzqAAAgAElEQVQK6suEjEny2PUzF0iOf/P3cLvd6nXbrfOxA//FcfAzBsPmVu2IP+IEcl+eAUSx9qbgqUrjdSSuPdoNT4ts8yTMlpcZKky9fy1MfH7ZxIUWkrBZv5nLyjiD9KR86+TxP8TjG8IkN7fu7WW+gyfG6lS9rvlpJERvdTqt+fCOuSP6qxN6xHLkqLit3e1EV7Z68dmBdifCfo2ai73BaKnfHxwLQWNxcaHb7odisdLrLS6vddeict1Rqz+KdBidECwyXNiVjtlxuLAJ9sShk2HuQ/rHPDLuPN/Uq2IKkJ8fLB777pW7PuqvR0ioVzTdhbnzH/Ha+4+/7QfMycHNKlRMhMf0DrQmpWAB75zXxrV72zi8XXhcrE5ECwI80c99Pz29vjmerxcrpsflV8QL+XcIHQshHqYYfDOLRdc8b6/iBNMiICHQpooPDSME/t9hhNgXXva8rY4QeYvDztwvrnSP/Njy/K0XHj30zLUP3PLS5d+8/bVj8fBbXvmE4P+kU017+FxF3esrhUAhUAgUAoVAIVAI7DkCJVjsOeR1wUKgECgEnozAVMgcPzgzvBGxgaAgLjEvCkQs0tGPXMQR0QFpJ6wNYs8u5Y8JQy4hcp3rVFj+SEZ0eM9OWTv6kEaZEfVKSa3r3YUZMss9jKm/3eNEG7u4kTOEmekd9AjuTMZ9vetf198AgQ0EjTEZHfMjFYP0cjBuEfHpTeMw+SiMbQWRjdRLMQs5bmwQLcSG9z5i0HiYTj49y/NgmizPpNaI/fGcjvBBd/RHzS3D0fBDQryIEEotbb0Q2Gk7IjTJf0KN9psP5kwS1LDdy/a7FuGE54R8IP8zzI5x4oUd4XaGb1SscdZDdUfwme/Gwq7X/Rq8FTZpStMQif75698aEZ+aiPjUiphQ7bOt1ujssBkd6EiaPhg9LXJTXOz3Bt3zayt3d+e6l9rt9krksAhNYzTsxCjuD0bHLi31n3ZpuX86PDL6C7cd6V1aXhsdOhApL7ZZgsROAt084UUBf2OIJ5PnMJdHATHOjJ/0cJu+ioTz7lW8nH6ks3K+1T90R2/U7sw1rXbv0rNe2Quh4qYNVzMRK3JDgvuTuZnhxYgX7lsptMLRvX6cKydEi36MF2Od59eb41EoPH3zbWHPDyNMbFb+Tnygb/95GAHTuiFc28p+2ZE/EXSnPfG0ldB6mWbPxkeBs/+5zDF9YBNKhuS0yYKQpFjbNi6t9sOxq+THQ/j7kWFr/vjygdsf+v1nf8UjD9/20taFzonucjPXXehF7L92a7i80nvCG3A3RejZQLZqUQgUAoVAIVAIFAI3MgIlWNzIvVttKwQKgf2GQIYKQDQhXYkPduIhMTwX95sHBY8JJIcfwa8KQ2iI8+6Y3DXuOwhNXgbIXI+OJ3QgQRBOPA32cofyTvXHE2F54oSea4vQGIg0bYQdQgA5AAdhNITMQAQhOFcQufvBq2SnANvP58ncKlMuGMZshpNKQU7/IuL8X5MEtmNSpDLu7Ur2XeS9cZKh0BzDk2IWQ2loX3pV5PMU6hCcxvbdgc2zYiKIg/7Cx1OGjKKNo1smggVhgAAqdBwC2s5s4o514z0TLK/HEFFT89H89chzgueXNjE7j9cXoi37i2F/L8yO41OT71+PNlzTNR8nsIetXq8Jd4rRYHGxG/kpWiu9tUE/cpEsh5PFgW6780ir2z4eKdNb891OOFgMu8ur/U5ITScOLcxHiovham8w+JDIZXE+CMvVtd5gnLfokDvHujKdZ2UiUqTogETlvXcyzC5v2JtPCFU7+NeXDc4+PkQIQuNUHe6PnBV/ODh4i3vUH4ZgcW7UXbhXaK3dEH+uqSP27suEAtgRI2w+sBYlke2eRUyEnbltHVPMXRsMLk3Ct8mbI7G9eSO8mlBPRCbrGy8liZuzWAPzt97fjOf6Qigh/WTu/3acx/owMx4vG3ia5Ro/7WmmfcN9Ilaot/lF8OOZpI/9TxZ51sdC02bF/2k/EGJfv2nPRfC3g++7dOeLHzxz58f+6YN3vnx+5ejJI4Pl1sFO6PnH261z58K/LnIVDebnOt1YA1xzLbDU/3Datnh5mfrUR4VAIVAIFAKFQCFQCOwpAiVY7CncdbFCoBAoBC6LAMI0BQQ/NJNEIlDYjWl3uJ2rCFaeF0hH5B1iiVjh+0gL30NgIEcy1A3CFoGvOH78Q3af9kcSt9oMgzFpG4bY8SNfmAWEEGJAG5Fu3h+H1whD0lXZ3wikaDW941bfJqk1HRLH8wyvkl4VyPrxzuYZFu3S+8G4zoS8HsfJ48OQ/CeN/wDj7nardW8IFOPEvPHoO9qM9PSeuTLtTcELyXrgfNMC4K6NiiBZNyvmqKTlvxuPiFm5eSQKlofklZep0CfHZ68PM9f/bJJvZFNi7jLX37U2b+PE7cg/0QqviYgENRouL/fvCo+KOyL3SHvYHx0ahmIx3x3eGiLFkQjwtbi0vKZP5SZZ6/dGc4P5kfG8Gokvzi+trJ0JIePi4nx37a7bj+S6P8aDUBEP7gdz8dzY8JyAxRDn7i8EX2R3eur5qvvMdgoRTA//YBivAfeY91161ieujToLcU9qfV68RtRP35e2c94b5pggj8f4Rz6Sw9F/xMU7o1MWY/3pR9+bz0fCncxcNr/N2fQGM099zjtK+LYxAT0JqXVpIlzo518J+7kwIv0Ph6WwOY2h67ofSu4sJJtx4ryPxHny/4INMd+r+ZMixGYeFVG5mSbgJ3MNhvpbvxClXhv22ZP3PiceeYf5P2WzYn3+hhD5nj7qLi71j979vgtPf8XpB1/8V1dPzz2je3Glf+vaoHWwvdAMF4eR5Gaue3BtMFxbWW2dj3XhMetHrBl5b5z2IrzMJeujQqAQKAQKgUKgECgEZguBEixmqz+qNoVAIXDzIuDHJWIi8zAgX/3gteMYqWj3a+4sRzAh6hF9mb+CSGHHpc88t+P8FyfHIKWEz2F7Hfd9N3o0f4jDBdEGI2QLoiwxRNTasYowsGM18UXmwAB28KqyTxDYIgeG0FEp9ulr/Wv+ZDLuzH+R4Vf2OgTS1aCc4xxZaayrM7I5vUN8ToiwZhyM9h8diy+jSNr8ODkcL1sL8b7v+g4i1LHWhxT7kNRjD5MgCAdBFl5PEVPfECyIFXaA2/mN6Pt/woQk0vYsjv3YsP8ahiyXVJjgYU4/KYH61Hdm8elYpF6c75wPxeJciBLnO63WI+1wq+itDefDy2I+Umy3YxVrR2S05XjdxGe9+Of9gfjiheXVXkSSaiIYzIiI0Q/vmsHBCAUVz8ci1JRQkQKWNZEQZA20FvKmIHp7TyLnFLUTq428XKZxfPOkD6zBSNhciwnk/Tu/9nsjWfm/lkw4k0rbUW487kfPvqseP9NiRZzkROhQIUCNPSAPxCQ+2h615gejUXcUodyiP89G7y3FvDVPzQFjxPxN0WmEzM9d85Ok9kLgESz0HwHP7v3XhK0PrUYIYYo+//KwfxHGu0mYtfvD/O9xPdeBceUmwsV0KLyrxn+vvhjzzX0mPWZsNNFvHq2z5lnOJ2KFzSfPW1c3HnAEJF4z947a3XcN5w+/69wzX/XQAy/6qoXlYydvX7vYO7Tc690S3hTdI4cWLsbqPgqPiqMry4Mm8t0MjhydXz372GAQgoVr+z+oO1nbb6o5t1d9XtcpBAqBQqAQKAQKgd1DoASL3cO2zlwIFAKFwHYRSCIiyUgk/HgHZhiy3Q/YzMGAVPDDk1cBou73woQZQG4kEWFnph+8SAfvSWTre+nBMX7MUDvbreSMHJc76FUnd5lrH6yQNZ4TaGCE7CHseI2oTU8UmEq+HZvSdy4M0LpkzQnXtAfANIRP7ATfhIifEbj3ZTVgm+GeNCB3m3s+jft+CZOBBMucNinAJImZIqZjjsYYtHYQK7QtY+WPk7FGSSEHgeaz9LBAauUac707PAVG3iPq/ZthPxBmffsbU5VTf3P6FZP3ELOfFQYX37UOWB9muo+RzsL8hOCwEknTz4UcISdRcNfjUH0nQp9YCO+LD7baozuGa6PYnd9aC1D6TacdatToln5/tBQ79gcHF9qLkbPi1gOL3dPHumvzd77xm/tP//3/lJ45xAL3Aese3Nw7JJ8nXvyDyWcJLVHbGLqcF9p98bmQNsbPfwlDshqX4zCDaVNJtYUjdN7M0UQsIyrdNOXW4wfbQTAfiH4+EcG+7g4vmqdFbK8Xx+DsRAKTxchg0m8PWytNaxQd2/RGw2Y5BjJMT8ec1l9CPrqf2YigPCkPyCSpPfyJkux1Yf43QJJ/0xZA/x/xufukNYC4ZKMD4anKFSAwCbFmnvH2JLDyACNMmEufFEYgnC7rPSzMSdjr59+O8Gm/tXrb884+8PF/e3T2jpctPNo6cqS9Org3xshiq2kdinEyd+Hi2j394WAphIvRQqwBa73RschhcTEEr9W5bvf0wnz7wYtLa8ZFKz1zrqBJdWghUAgUAoVAIVAIFALXFYESLK4r/HXxQqAQuJkQuAyhjchhSBykOoLpZJjdxnZOIieIEEisjwxDRCDr7NZDTmb4GwSHXZZyXSAnEU9+rCKqnDt3Te5XscJwmfauEB4F+UWsQBD4DGGAfMmkzMibDI0BM6EWksDeTExwnZ0oKURlvbOfcnd/9sdMk6o7AcRenGMD4Wca1/2Kcf6fZiyZ6zmeM/yZOW9cy2NxMDBIEcLYEhoKWWYNcB7PrS2IM+sMUdQaI5b9+HwbxI/Pnc570YXT19Bf2mDX/veFJcn+7ZtURA4bCYV/Moz3gN3LyP/94G0xXF3rr7QXuueC1D4TiYXu6nY7a0FMXoqAZR9YiTBP+jUAOdGO6C+Rs6IVysXhufn2SqvprLaa4cVOM/zAfLO2dPjSQ2vP+aPvaY6/8/VCL1kXCT3pNfGOeO6e8Alhrw77qg2wNJY2WheJDl8WxkNCXxCS3IcIEeMQZZdJ3kwYSaHNjnKeBTcNIS5PSavVLLRa7cORV/1w3Hw+JFxgnh+kM6y7rU7rbMhq0S+jbvT7xfCQunvQDA+GaPGBIJ7NUQIcMQER7l5ufOuj9WtahnbjIWFO83JxP+QFY+6nuLe+260rfy3MvdFc05/3hZl/e5LQfn2FZvF1CBKbldxEMZ0HhmcYr9gMubbRd1NI9hkB8J+FEYysWY+cecXfvnTuxX+l8+jwwNGl/tw9y5fWntG0BndF+Ldbl9d6cyFMHGu32rdHp7e6nd6jMciW5udaxw8fmH8kYsw9srbWH4aqeenI4fnVEDbGSdZLtJjFkVV1KgQKgUKgECgECoHNECjBosZGIVAIFALXHwE/JpED06EfkA+IIQXZgBhCziObiBdii/uB/KIwpKPieOIGghIpZI1PocPz8e7XfepZkb2UpIwf9UhWbc0E5eP4/WGEDHjZjZox+jMcgt2LPs+kzXnenXxMAsO14e61unqOfFKEaxiH4glSedz35Wmxk11wQ5zLWDdOMxdNjqWxGBFmTJsHCEaE8p08LMTEn3xm3OW4TwEgw0sZf+ZLhlEb76ifsSS26qxt7wyz9lnnkLZCF4kHv758QbzxmWHfFcbj4r4wxC3vsiftSN/gu9fzLf25FgvBxWjwI6Ph6M+Egor37pDWYjBoBbk/jEhQ7XZ3Pijv4Wg1xIy5uFucnu+svafbW2ode+zU8NbR2aVDyw+uHnznzz6r3Vv64gkG+lXYJ2S0HdxIckTqyU0aPC1WwN+Ob+soIpUAxHPP+il00HZD6vF2IZow/bk+7NT1xH5Xr02sOHZksbu6OjgUbjNHFubat671B/dGXx6dX+h+cHW1/7RIsu6zQ91mtNDptg5ENouDkVjn9vC96EZorzPhZXM6OuU9MT7MV4IT0WKr8D7GFNx/PExeKxsfhIj622EEpI0KIZOI9elhcsMg0QlTKfLvKlb78OS5IWEsPIUJsWVDifWG98RLN2iT+7+1LAsvWflGzFPPrXHnT7/y7zeXTr6ifX7+9vYjZy+2emsr8+eXeiFADw+G0HViZXVw26A/mh+2BscHo9aw243lLbwq4rsL0fG3zc11ViMkVDe8eCK0WHMxEnFHRu5B/p+5D6GuKhcChUAhUAgUAoXAzYhACRY3Y69XmwuBQmCWEMgfvX6wIqmS2FZHP3rt0CM6ICoQBwh3QoUdxAiFF4T5gfwHYcg63gV2ZSKb7LS0oxpZlwk19+tO8+k+y3Al41AHk/bzNkHovDUMUYCUgU/Gvke0nQxD0CJy4LBbHhbOm7vZ4a9Pk3wmUrj32tWaYWvG5PNEuEhB5on2lpAx3fU33fMM7ZShnzJpeHpQIYDtpGaEO2SytcL3eFLJ7TEtoPk+wsx8sW4QNnN8zurakGuZ+iL3hLARhogXwfri/W+YvPm18WjeKzNL1skbEsR2f36uGzukmwcHIVYEKRk84+i45932qN/rDx/rN6M/a/rDhUjGHWz1cKW91n/oWPPQ3Qf65y/c8/BbPuy2R972nKNn33lxvnfhcDMavjzaTNix3ul/6yDviO2UH42DkJ+EIvlEjBeeLu4hxk/mgdnOuRyDYPc99y7r801V5ufa7Uv9fkhNzeEgkZ8T8vQ90ZdPG6z27hkMmyMhSKxEZMLjMWMXIwvJgzFnu6FOLXRGIUC2m/f2Y0u9UFLxuXmQCdO3g6Hj9dlvhZnnvxTGK8Z44Im0UTFemLEjXFjm0Ho4PAymw+w95bt7lZR7Ow3fo2PGYfjCXhZmvphzhEIbRwirGxVCsQJLItJbwv5nGLGCsHSBp9Jbv/nvjz1oHvyzs62l5d58eF4txBpwLLY3PGfYhDYZYcRC3FoZDGL8jAa3rK6N+gfmuhK2f7DHW6vVuuXAwtzpZr673BsMBp1e65EYV2fCk2uWhds96ra6TCFQCBQChUAhUAjsFwRKsNgvPVX1LAQKgRsVgdz5bNcpYojIkOGM7LbLcBDWa6QkEp5XBcKbl4UEm8hHP0R9DzFktzXS0u5rP6q9j7y87ok0d6gTEfy5O9yuUKKOuPww8ah4j3ABw2eGwVVBxiB1d2vXaApQiCViBUIDYcfjQ8l48vrTe/o/+2q80zps7HkxOb4ebm4EUugyv9MDCyKeGyd2vxMprR/GXiReDoUiSM94bu6nCJHnSTR9RvBjmdtmnMx3fdkrr4stCM9hEKbqinD95jCiLVLVjvHpncwfMVX//zBp34/F41x83zq4NJVbYZZG1ujCpdXVo4cWzoZYMRfEdiTQjVj1rdGti93WHXPDHvFi8UCfrjnqDbqLy8eHF+ZueeyP528/+3v33nHu7S85cOH9t871Lh4MseJq2uXeYixZk+BljTRGrFenwnxuvOX96kquAXeiO4JWaKNZFcaupE3bPbZ1+uzSXKfdPtDttm8Nb4o7Qrg4GDN1GP18rNMeHQ9J8eHeYGS+Rt+NIsxP69HwrIh72eiWQOqumNbz8b0Lo1HsqR+N5wAct5sDBDGuT/0f4XvuS4Sjvxr2nyZ9vFFbEOsSdxOYfjuMx8XvT86V42C7GNxIx/nfw7zIEH1C0fHmMsb/Vpi1+HKFxxLxT3/z/rovjKh6KdYluI7Li59+dPTGt3+w1e8POytrIU/GetBut+Yj90l3bW20GOPjUnhbHIjkNyFOhldFiJjLTf9IjKl4a/hot9O5MD/fOd9pd45FTc/E68H83KAVgsWN1BfVlkKgECgECoFCoBC4wREoweIG7+BqXiFQCOwLBJIwRC4gCvyq9COWICHZJvIdWYD8PhnGewAxj7SwoxhpT7SwwxoRj7x0HgSFH9LjOO6P85itG4Es0gY/7lOQ0ckpzIjbnqFzPCdQwM0OY5imZ8UY5wkoO4lJChbq5Lx5n1VXgoq+41mB+FAnYoX+TiIvvUf2Q+x9bayyewgkOTw9jlwNmZyhoHhY2AWNyMyd78KMmeuZGyfP47XxlTlUMkGyNcJ7LUmgd68513zmFPSEIzKnYfCtYZ8b9hWbnP118b74/DwFrKG/HsKFXefDWRIuJl4Wo/OXVi8cPrTQP9y7MDi28tCJVr/XifAuJ0bD/i39uUOjw+3BSnvp0dHy+dXeCx74H59+bOl9z+0OVpuFwcVmrr8UfhlbRQoao+Qe4Z5hzTF2CKo/HWYc2OktDBCCG76E3rFXxTXgZUw5t2va6b/Z7v5NunB/vi0cVNR8HHotyOZbgzi+M6J6HY5BPAxR4lx4XvQjAffB8J6YiztFLxwouiFMdDqdZjV2zJ9ohbKxMNc5FhLVUoQJOxAk9XsHoyGxwRx+infgZQS/8byJca8f09tKf399mNBqn3EZhF8cn7Hxpocw91DC1hPk+v7snafWehs5KtzL3a/978WL1XN5Qf7mNjHgHUYAIiDBkQcTr7ENxadHzi01EcZpbmW114m1/Fj4YN4S42huEIMgfG6OxhI/F+8/FGND+KeFyG/TiZwVK6Nhe7gcAeYWQgWLUFBH4zuLBxa6g6XV8Nf58/CC26xyHVYIFAKFQCFQCBQChcD1Q6AEi+uHfV25ECgECoFEIElEpKMflciAjPnttRADfiBLmipcxyeHIZJ+LQxhabexnbDICF4aCE1iB3IjQ6FgMGeZjNzuaEiiJsnLP5xgdXKChZ3AQsVkCBPkAMFHCC0YEQxgk7H8d2PLYQomSD+iBNFE0aeur38IUYjTTAhOxCA4IbhY7oinqYy/fIP033b7uY57MgIZMi6FLPPAemEdMI4QYMjgJEmJFpHot2XeS75tHcg8Npn7Ij0sPO6ntcHcz13jSHdF3H0C5UblE+NN8w5RzyvjVBiiPr2u9mSsbUCI5lr2ePLd+152sNdZPHTpwF0Ly4u33dufO/yRvfbCrYO5Q3c2vZW7V+aOv32x1Tty6MKpz2z3lo8f7J8bixTdSHowXtq351lBLPieMF4phAqCN1zkpzDGYGIdmt5Ff61jw3j7jbBM/L6nuO9J525+kXan027andZyO+SkYJ7XYkJykzkezjKDAPZCCBaHpCeJHfMr8d58zNeDoVXEpvj2/Px8+0ivP7qwNhzcsjDf+d2VtdFSCBdXdc+aCE7jvoyx6D7Ja8JcMP8/NYzX4mYFKW9TxLeEuX8h2vXjthSy69wH13J5czRzrlhDPjrMPV2+CiGgrC2XK8TVnwrj5ck7lmgKc/POWn45/MZedCFicay6NcSLW9ut0S1z3c6hTmjRg2Y8Vh4bNSFSxP8MUdHFWP2FEY3wcq3TkSel4W0Rn9312KXB+3u94drtt0SqlBu/z66lv+u7hUAhUAgUAoVAITBDCJRgMUOdUVUpBAqBmxaB3PGcyXQBkbueJUplRAk/cJELmdPCDr8MIeU5Qt4xdkASK5AT413XNyDZjURAnCBRxIsWigHxh1TQZqQbggApZzc2gvNUGDEDWZOCBax3o6hfkn7utZ4jhNRZGAm7jZEXRChhbCTr1GfGgPqpNw+ZJKfaUzkunlTfynGxG903M+c0h1kmmU8hy5jy3Dg33wlyKYwJ+0K4JHbFZu4nSDFjkMCZc4GoJ26694yzDYnpf/H6320FWZaAbHjMXoWNmuqV9LIiCorN/0/CviwMEW+OrS/m118O+zdhklB/IEjbX5/g1xM3fg973DqVuQg8WrsQo8+cG6y84PjFP105svzg2V7nwMqgPX9r7Ln/6Naw/6yICPSCYatrtzX1MsSKS007PCra0W08K1obCxa/GOcl6iJMeU7kDm/vqwdCVdg842scN3/KdgoS657Qhe5PYo5NJx3eqWvM9HliV7xMMvOjGGYRHmoQcXuWhPkJ8aETiPfDtSJycbdiDg4X4sgT3KOiK+Yi/M8dQTrzBDwTvXx7TOal4ePK1FM8LK4EAOLFRLT4+fjeqTBhnz48zBzZrLw2PviUMGHY7gsjWqiL9eNK85pcSXWvx7HpiWLzgM0i1pTc/PCl8ZxnxVbF/2nyU8D2zWFECuvtekFww/O8+/5HmuNHFtshaA1j/MS1R2shbC0PY4bGcIL5HaFTLoZnzoMSbkdHnIhKH+4NR6GPtTtra2vzsddh6cDBuXDQGoYI1opQUeGHUaUQKAQKgUKgECgECoF9gkAJFvuko6qahUAhcEMjkCGh/Dj2w9/ajIhLDwlEI7KHKIGcRGanVwbSCeHls/whTOzw/jhJ5g1IaMMLRjwn7Kq2WxrpRgTwg5y44zkM7D5HljnWLt/EMnf5Jkm3UwMsiST1Uw9iSXrMEEsQHykkIfKeFyYZrv79nUm/Io/tlERuaJdx4HvOkyJIEQ871WP74zzpUZQhx8ztDINmjJ8KQ37n+8a8MXh7kFbeN6aQXMYPQcyceTTWhvfHDt61uW53YWGhPfcd//1tsZm36ccO71Z/OGwHUdYPsSJJ7L0k9bfbK9rFO+kHwwi7vNG+MuwzNzjBJ8V7yHK7pH8l7F+FmWPvC/L2zE6LFnHOJD3h57k5LCyc/iBaWret5y8IQ4omIfrSzmDlcGvY+5XIbxAuMu1njcYpSVpBbse+6s4cb6umPQyNYex9RbCIrnmyYAETbeRN4b7g/sAbhTBhvPh8fN+Jdu/2LnnCq375uDBr4u+G3Qxl7NUUYsPh8JYYhtLEpaIVDheExLlwgVoL8eJCzD85Ldz710LDiI5t9VqDVm80GB6Id1sR0mep1XRWopMPjpp25F8ejkN0XSuAE48LoaIIWvJevSRMEmhJ63kibVTcs/5K2OeH/WwYMt699E/jPO5TzTWEDrvWJu3U9/Wb/vC/hf8bToZ9Vph7+Wu2eZH/HsdZZ5mNCbw6/U+XG1G2c5rW8mp/HLaSQhkPj4XecCYi/R0PTwsDIyJDje6IpYCCaZzFMaGB8cCJTNsxuW+JsTY4uNDtHzy2cKLTah6IvBb1f8N2kK9jCoFCoBAoBAqBQmAmECjBYia6oSpRCBQCNwMCmwgH4zQK0f4M3YSMQMKllwCCDbGF5BLyJXdDI52QTyl2ZEghUEHzEc4AACAASURBVOZu6Rvxx2mS/Um8IfyQAIh/pJj40kgx5AnRIkPkIHBhCSfEIQKPt0oKPzsxBFP8UDfk4zjJ76Q+JyeveVQQKNTVrm/iU5KZvEXUX5vslvcaoSpci/HgWPXXvzsttOxE++sc14DAFl4KEmKvFwyMiQwNRdhSHCMPAQKcKUhGZFl67hj3HxT/3M7uubn2fFCoz1ha6YVQESFrRqNLg5FY6M0gaK9M9t1c7/wWW8TofywIU54W2io8lvXxSzbojkzQ/QnxmQTeEt9aV98W3ze/Ng2PtUVScGF29IX1JPMQWW/UJ72rXFsouFNhwsrwrHJ9x9m5zgNCnwk30wrvCevX2cc9J6Krx5vuY/kjWrRaD8b750KksJY5F/KYx8jjyZsfvzfAgeeN59YNY8B9pr/HpLIx5B6WIrF72M1QxiF9gkA+1+8PDkcW9Udjs/xtrbnmgZhnC0EvR86BECkiPFRsmT8cctSZTtNeCi66G50fcb7aS5HD4n5JkyPZ8iORufv0xUurvdXV/pqcJzsF4GQsnI7xy+uGBwyvgK8I47W0UUnvAqKgY98YxnvA/LsQ5yGC7Vj9dqqdlztP1Nm8zYTahAmCDXHiZBhvyc+7zPe19fGwbo+LhD8QdirMuHfvtjb7X0C5kv/JRpEkO5wqWtb5QUz/x8Jx4miImPcMhq07RiEoR4UXYw2/M8SvQf/x/wr6cdxa6F7DuU7rSORB6UXi7qVer38p0t70H37k0lWFE9uLPqhrFAKFQCFQCBQChUAhsB6BEixqTBQChUAhcP0RGBMb45+bjxOOyHbPM94w8i1/6I53YoalYOHHNCLK91K8cOy+IgyusAu0LxNIaj9yIb0okH9+4BMtEGQIQTsl/VBPMhNhlslkdxKn3Emdu1+JTAjF7CPhV9QDoSxEi74UP94OZOE4EJjqTexQL8SJY54T5ty5Q1p/j0mMK8StDt/HCKRgMBEucq1ITyrjyvgwJowpopeQLcaSOWEHtXXFmrIWpBbS9OHgvw8GoXo03CqWQqhYjFmFGY+tuxGrpt3KNWV0vcWKbXabNdS6KNQVsvVXw/7tZb47nSz3O+K4/xHGy8mchSfx4gmPpiA115ONKTRnfhDfI0QKUUccIhy8LMy6Q3wgRvKwyJwj1iVzG5lPnFQ+dqq+QlcRLGN9GN0WYsUfxPOTIVicCVIbSexcQvoI85T1TAFL/fV3JmPPpNnXY82wNqf3j7Zb765LmSTCftK1d3Fs5/gIbnl0aNQePRbk8p9EboET4TATzhbSVgyfFR4T3RAkljrd9gcigfLF8Gy61+aGyL4tN8FoLUjrAwfmlrvdzoWF+e7KXbdfLtXENcGa/1cg1+W3MH7+QZixu1lB6vMe8B0CvDXoXMwVHlwS2+/k/fWaGrfRlycio3usUJKKcfqiMHOdJ5AQWebt5cr/ig9tMDC3CITmPm8v6/B4g8k1CIQxHEZnwkOH8CGE2OH4z3A17LHIiSJD+6PyWvR6o07k4n4wQkEdjrHTi3F0Jo4NvavzgaXltYcvXFo7F+t570OfeWvrre8/37z46UevRDjZcdzrhIVAIVAIFAKFQCFQCGwHgRIstoNSHVMIFAKFwO4jkJ4DSUAiu/x4RgQI6YE8QGArCILcCZzho3w/Q0V4VG7EH6UZrgE5aGc0TBAFyLuMXU8Q8BmBwM7Pj5och4hAICATHDPek8jDZQdzfCTmdmuqk0feHK6L+EFs6DtkBnFCmCh9TFhJwcmOTH2IKNE+9USqZEgoZJDd4M7pOzdiP0ezqkwjEGRrvtTn6WGThKAxYkyIm06MI2oRKZDDGE477H0HYRwbcpvQKIanY/du+FW0ztu7H9YJkismQ7ManhXLg8HjIuguErq70cHqnMmkf2LSXjHnNwoRNX39vxUveD59V5j1wvwkCijmW4bbmw7JZX5bp81jZK3PiA+M0KAvrE0EBeuWkEiESmuT53eFpQcdYSlzkGS9eI0x1+d94ZzWLufy/J1hQvggW5Gk+lzJxOzpaZfnu16P7lHwhCGvj3HooJ0uU/Njo1NnqL7cCZ/zph3fy5Bn+b0N19OrzNMy9miZ9M+5hYXOwX5v+IKD8/OHI3rPsdWV6NtWcymI5dsiwXYnpt8oek8YoEii3Op1Oq2LB1pzf7bQ7X7w6MG5SwfmO0JC7eZ6Dxf3J/9jvCFM3xmvwkVJbL9R+ZrJmwTSHwtD4LufXQpBwBq0cg2E/U4Pk/H5ol4pMmqf5+ahHB1EQv8bEBK/aBsX/z/jGF6T5ry1wDwkWpj71yJUuLR+HgunsR6fD7GrNegP25EE5aEYJePQlmv9/mr870JgviuOjmHUjjB/zaFBfxAeGe3VOMHqgcX5EDZa80cOLczfeuxg5hvZRtPqkEKgECgECoFCoBAoBK4vAiVYXF/86+qFQCFQCIzjkUfBVfgR6sdzEhL5Yzp36qco4fjcYY9geCJsy+S7u0loXM8emw65hJyzi9xjxoZXN2QlAsFOZ7s9kWOIFGIBHIVksVsxwzhkKK6datc09p4jfwgS+la4F7uNhaI5Gcbzgpjx8ZM+1KfqaVf2qcl37fIkaqi38YDURIYQY5xT7GqPN2Kukp3qkxviPOsI0xxnT4y3IF6NH2R1ktfEstzpn+HjEOOZsPuxcbzzx5MfpI2ximtdj534O9VP2qK9xBrzx/wn+H3qFhf4tPicKcQA5PqrwgiIPxlmrSA4OL9zIv94dxEueEiZ64zAwGNCCCiCoxBPCFzzX/gmHhjECvNf/1i/xzlFJuf0nvXrVJg17xcmz5H+1g/X/6Mw7SNOOV7i8FntsxSRjD1Cy66EpdlIUIg5YQ4oud7nfMl7SXrFTb/v+Gu+hwrbFNc3RtShH0rDsfMXRpe63QjntdKbD3L5YnhadFu95tmhQSxE+J/VdqfzUHg+RSb11tHII/NouF48ECLHmVa7eTRcMi4cWJzrveYl9+y214LzG1eId2NfHgf3Uu243BwyNr82zLj/d2EEKve6syEQeH5ZXLcKuTb5/qYPcY31ZX3YRPPXe+YrEca9lshAnOHdSLCQT8ZnlytEGJ5Y1hT9SxC2MSI9VOTDyU0jW1V7088JxRNvOvW+EGPk/hAqWoPR4EiMkafFaxm0I+pTsxLC82PtGCxz3QgkF6GiIr9FhPQbXZzrdB8KzxzedKeXlnqrRw4ORuVdcdVdUl8sBAqBQqAQKAQKgT1GoASLPQa8LlcIFAKFwGUQQJIkGTEmocOSUEdGZdLczLswHQKK8HHNJMuM906SS9qPaECq2NlshzHyL8NoIfgdi5jwSBRAHCL4MhyT50iUjC29k03PcD1JZti9md4SyBDkZnqHaIO6+Y76jBMlT+qqTd7zGUIF0Yf00yZCjOfpkTPO5Dr57EltuQGTru9kX90w55oQXLmr3nphPBD0EGuK10g1ZTqk2H7zothOn2lrelMRNv9l2NvCCH5ftY0TECJ+Zuo43zMX5b4wXxHvr5t8jrBkknkTRbnC8IywRp0MM1et1eYw4ZG3i3nL24XwITSUee+crkGgQBL7nGcFQSKFEGuBPs77gyrM7Lof4WfUl/hiLUYME4G0ZdfKJOyT6+b9IPHZaJwjhZPIfpL3xQ55FqU3lDl4R5DJkfa4Ezvkhxya7lqMxBS99vBgSIbhcdEMIh/3+bm5zmrkTF49uDj3vthV/1DTHp2dm+tePH54YeX40QO7IvZs0hnqnrmY9Jl7JrHcvSyFvY2+SnD/vskHXxePhDiJp917rT/pKTgtGu30eDCfzEX/K1gHzEWmTeagMenzF4cRY9T5EyeVMA/TY2J9vaybXx5GdPQdc1TS8mzbTodqNHadczlu7xfDDe5M+MK9Oxrhn73IPdS0Q5C4PQSts8Nh0478JtFPo3Nz3c4HY6Ccn59rX4z8FeM1/8TRA4MLlzhdVCkECoFCoBAoBAqBQmB/IFCCxf7op6plIVAI3DwIpGiRybf9qPeDNb0oMgTQEzuib0JCGtFAhGCZSBuxgiRELPKyQATCDLmI/EviCLHo+3ZA2/W8G4JF9mGSx0hjhA+vCKEmkD6KOqinOupvxIk6IVjUUXuQKIg+n2ur+PwIWOfWfo/u5enFMau7rCdNrofdRGBCsvYn3hbWDuPGePIceZdCxlgY3SFSdjebdK3nTu+FN8WJ3h4mLBxPhb8RlnHrt3ONf7TBQchO5KbwTuY4fBGZn7HBsULqZMi6zAlgLvMGU7f7wniDWBOsD4QKQgeSGJGOdNR3uf5vp86zcIxxx5skPU0y99Ju1i3HehLi43vnZiGdJp4QKXCMvSHCxrvbd2h+pIeJdTsSJo+T2t/fD1miP+g8emCh81is4LfE5vmT0dG3xc3jkW6nc3/kq3hnCBwPLS7MXQzh4mx4ZOTc3U3sNjq39eNUGFJeUmn9KTTZdA6Yzer07yfjVni27wkzP4wB+Vjcp923ifatiYfE9KaNJ51zGx4Y6U3j0b3yQ8PcF913CY3PDeOZxBOEpwgR7RVh5uO01woB0f13uph/fzfM/xfWDef93rBTYeNwcbsR9moiQqdocSE84ubb7aYX4kV4VjbxvHUgpIv2IAZUfDbstNvDGCdrIXD1D3RbD3fanfcvzLfm4wTj0GRf9AnP3m3vnHWw1ctCoBAoBAqBQqAQKASuHoESLK4eu/pmIVAIFAK7hUD+QB3HipqUJL9v9h1yuUscSYCUQPAjHHgs/EkY7wVEBTICEYIYsasXyYD8cyySMT0VksTd6b5EDGTCW4+5M5ZAkbulkQjCxSBIEJ5i3QtJ4d5sN6hdoK8OkwzY98TKJ3ho95vDEKBIJOOEN0aKWDf7GNnpvtwX51sXw3+9t81Y+NwhAnYm8bgMoQmLfhCi5hDClWAhrEsKAdYLIoPHKyni3TNlqzAyKVbk+TOknXj/iFuvrUtCyyBDs//GpPtukKFX0tBrODY9QpDGdrYjgndtfZp4V1jT8x66odfZ+vZMiOEnEqxPxobDrkkATjFEiLWoGwHqg5GPoBWJkBdjF3yMwdHBtU5zsdNqHVrpD7uRUOlEbEB44OihxUcuLa890GpGHwiPC95zvchBML6HSJq8UYlQP9fQTXEzISdsXgYxf9y3iBfG6g9Nxus3xePlknI7o/74ixPjaUGo+9kwYdcyP4wx756nDwgamY/L98ck+0TQyP+Jcgw5d3rSuMerC9HP88+dnPNH49HYM8edV66a9fli0rvGpdaLFV88qQPByfWIHvpSna9pfLhYlsvkYMkQd/5nWQthQgiod0Uk0TvCWiGADcPr4kiEGnssBIuL8Xkv3roYWSweWesNH+72W+ci78mFxfluiRXTgNfzQqAQKAQKgUKgEJh5BEqwmPkuqgoWAoXAzYLABp4S08TOjv0w3ud45q5ZOx5TdHh5PM/d0rwOkAlIQCSFXdCIBe+Jp43Q4GWBfJkWhHYaluy7zB1AbLC71KO+VAfCA4JSnb2PTBHOirDC2wIxdDKMCOM1QhXZQqSREJUgMx3OxHP39RS3drpNdb4ZRmCLpMC7RhLPMCRPqloQsgi7C0F8ij9PyCQImosIUqSmUFHCvexFMfeJjPpFyCfrBDJ4faLe/d5vCN5nhsndQUSe3+UY+ukpkULFleJnPKTg0dkpL4uJkOI+5J5lHB6JnBarw2Hr0f5g1Dt4cO7h+UiYvLzae978XOdUENEPra0NJN++dCjyzPTDArfrTTgnptrw22HuSeaOhPYEObh90mRcbzaHhHBkBIx/HfZfw9yLzYdPCYMR7w33ayJXehWZHwQNobUoM+O5EmYO8/hwr3cvNdaEZnMfdK+0GcA937F/YbNKbfA+jxDt/J9hQsllSEZiBZFlx/8f22r9jjGU/0sMQ5QYxf+Ly7F69IeD0cqoGd0T74yG7eGlECfOxdg6FSHFep1u+/ylpbWL83Pdwbvvf+RK58IVwFWHFgKFQCFQCBQChUAhsPMIlGCx85jWGQuBQqAQKAR2D4EM9yDGNBMPPsOm2KHM4wBxj8ggBCA5kCF2QBMJCBsM8YEA2M2Y4EkQIJpcBwmjDsgWdRLr3m5TQspXhglX477MECPCWGijkDN2oyJfpneeptChjXBBIGUi3gwhFm9VKQQKgURg4q2wHMKFhMLWAesFrwveF+aS+UkM/OrJd6wTiHCP5u1OFEm8zX0eVdYwYaDGhHAmD95GCJydqMdun4MoYw1DaCOAN3YP2IFaTEQBfZlhha6GoE1S3riwDkucfU2eSenVNAnTlrlHxiH9Ynf8BwbDwdzS0uixyEXwaIT26Qw7o4cj7E/sjh8shGAxvkfNWCgfGGWopR+M578eRow6FUa8eB3cwqa9Fjbq4W+INz9qctwz4vFkGDGA96DwaD82+ZLxwzvKXHGMEI/GU977Ycl7gojvGIKI87lfKlt5gGTdfiqeEDzeEvYjk+c+43HxG2HEGe2+XsJRijfauxJj47EQuyK/div+r2g9MGqGc/2Bl83Z8LQ4HWOr1xk1vch70nvw9IWdCm+WWNVjIVAIFAKFQCFQCBQCu45ACRa7DnFdoBAoBAqBQmCHEEAaIguQiYh5ogRSRI4HRIOdlhlyCcmQ8dL90BcmAqnhfUkyEWcpVqTXxjVVc5NcInJhuz6xgseE6xItMs+G+iNkCCrakyIKcs9rnhc+c4z3fFcYqc8KQ6IgZpBrDGmkLcLduNa2wqFcU6Pry4XAPkVg4nGxGgKBOfPHYUK+ZE6ZXGsQquastcUas1WxpshJcTJMcuL1AgfvDru3vy9MTH3zm8eU6+74ru2tKrsHn8PR2pQhsGC8myXXvGshlfWD30fprbEj94c4n7oRLIjL7k1Id9da6fWHc2HW/jNxv1h66JGLER2q6YdoMZrhnfHao1/dT917mJBP3xjG42E7OS54QJoDWYRqeu3E/kk8EvN5WhD0PjmMt+F04ekh15P7IrHkaguR4u+E6Q/3V2KITQLms/vues+nq73OVX9vInzJrZKCHPGkG94WEm1/sNVpw98g662s9ZfiP4lxzpMbOQzgVYNZXywECoFCoBAoBAqBfYFACRb7opuqkoVAIVAIFAITBJKI8qMd2c/LwA9zpJ+QSUgLO6cJE3Zi2jmNPEH4u+c5TsgJnyNKiB9sN4u6JhmZ8eozXjpS81VhiE3kj/opHxtmd7L31BM5IRcHwgap8wVhCE9Eq3Nrp9AaSIv04pjGajfbV+cuBPY7AuYoYlIemVwXfimeCysjVI3iM0Jphm1DMCNcPRIihKr5rjDrCZGRSOk9xxMfJfuVTDtzAZi71gEhoRCiN2KxzlqvrGO8xhD1u1l2SqRFVGdoqBbvjR0gfqc9P9wHjAP3MGt7FvkGVvuDJ/IRjZOsy2+wRcig3cR0q3O7/+hfZszzknhlmHBKhDi5pf7pJicx14gR7tUbFYIh26y8dN0HvCyJ+JcrvDdeMjmAMMEz47+F+a7/Ecxn45SnVSa5vxpvnS2qcXUfp3Dh2zEu0mNnFLlR1HcstE4lkr+6i9S3CoFCoBAoBAqBQqAQmAEESrCYgU6oKhQChUAhUAhsC4EUKexMRfAjw5AjSQwiH5Am07kpPj5e+1GPFEFCiV2PhLDr1w9898E2N4jwkNgVUmLieeESGaYp65f5JhCXyDzkaIYiIcQgTtSdB4mdpuOkm2FCXCC6xOxmcMikvq5B6MhEpJXPIsCoUghshsAkRFSGYjLXCJ4p9vFWsmuc4OA5QVA8e2Khnd/C1lhzCBknJ8/NRV4Z5qg1CWGr+Dx32XvtfMjeG9GzIuGGFwys03axW892s+yUYKH/9ctO5zmarl8+J1jkddbXf1fuSVfTAVsIauN6hreS+5M5JLwSgd29StuIAkIbul+tFyA2EyuutJr6TEg3xdySN2V9ETbxP4WZt3Jd/JcwnhRENfM2PYHG3glXWoHdPH6TpNzq6B4/PX4IGaoyrn9+b4YFr92Erc5dCBQChUAhUAgUAvsYgRIs9nHnVdULgUKgELjJEMgQHRmmwQ5V3gS8EoRseWEYsh7pb+cmIcOPdmIFcpEHhvjWPCx8F5E4Dp20W2LFBv2DVLFzVx3VldnZeTKMSKG+3pOLA/EjDre6Il/s2v61sE8Kcx7f027FOYW94mmBPIWRe3wnhJIm2nctIVIml6iHQuCGR8A8mZ4rvCXMv8yNY956j/DJM4Loae4piPkUIDxmPoUUJIgYjkXqOudMEaK71LPwuS+MJ8rSbibc3gEPiGkI1gsLOw3P+nG2XhjZl2NjEmZN286GeIE1f2bYybAfDyO6m0eSX7s3fVoYD6SdKhle0flSrPjpeG6u8mQk+Lu3mo+8LLz/jjDz0n3T/wLpUbFTddqx82yVlHvHLlQnKgQKgUKgECgECoFCYEYQKMFiRjqiqlEIFAKFQCGwJQJJItkJaUckUv7lYXao2snrnibUhh2bdvTaTWnHJfICUeh4xASSBJHic2TFTu+i3aohuXtTfbVJ+Al2KgypQmBRN+Eu7EpF+hEutFu7CBLOQaAR19v37g4j0NwXJnTN28KQokiYweMOJLvjQbJVY+vzQmA/IHCZHeTjXcyTZNjEhgwh5/3ptWN54q3xlOZO8mT4rrJTORFmGta3vv+8dhJZrU3pbTLTdV5XOfeLrRJHb7s9NyHhnGEMCeu/GnY8zEYCHkuw/ZkwoZncs20k+IQw92avfe74qylCuRFG5LdghEXX5YloTBIp3BfdT/Naw83m7tVUoL5TCBQChUAhUAgUAoVAIXDtCJRgce0Y1hkKgUKgECgE9gaBDHPEEwERRqRI4QKRn0QIMUJIiF8Is5tT/grEBM8KZCMixG7oJ5JuXwdCH9lJiBDjmxEo7PgksCD4EDgfFib0jPfUW3vfHWa3KsHiL4WJj8/eHmZ3qHAbzwkTekVIDiRphhzZl7t2o/5VCoHrjsCUoDE9j7Y1p9aRodv6znVv8LVXgDeK9deudrk7CK37qaQgdbP01472zWTME/qm8ze5zwnB5F7Oy+G+MOHWfj2MR4axQiRyr8v788viuXv7z4a5J0qyzavyq8LkhXFfJ+h/b9hvhBEknMMmBf8XuL5ruj96PzcMXCqRItCoUggUAoVAIVAIFAKFwIwiUILFjHZMVasQKAQKgUJgQwSQDUgIOSwQ+feFCfVEuGCICwR9kmO8LYSNQmzYVWnnpR2XSCi7LgkZux1XfaOGuL62EC0Qe8gVhAryhuigbj4XtoonhefEB8cIb6GNhBcEDGLHccggYgUvkvzcdzIXxkb1qPcKgUKgENgNBOyWt7ZZi98R4aCuxzp7Le2yRlcovWtBML6bosDEQykxJVi4bxHieRQSFHgF8oIgWri/Ey3cy5h7ts+JHClqGFfGF5HiZBhRw7lcw30x85CMPTMnguONnC/mGnuqvl4IFAKFQCFQCBQChcBsIVCCxWz1R9WmECgECoFC4PIIIDqQFIpHJBiCnzDBq8Jr+Sp+JwyxwSNBaCThH3hlIDw8plCAFEHu527OvcQ/d+66NjEFyUJAQcwQLIgrH5zUz2s7R9VXslDtcQ/nleF7vCw+PEySU+LMH07ehwksTk8SixcBt5c9XNcqBG5eBAjF1llrmHVtP5byrtihXlsXci1xzcdLIWgYK5mnylXd390bv3PyvvscEz7RsT8YlmGe0oMic4Pk/bz6b4f6r05TCBQChUAhUAgUAoXAXiNQgsVeI17XKwQKgUKgELhaBJLMSK+CDBH1QJyQOCFUErJeLGwJPdODgSeGMFLIft4YBA3eCHZ3Zlz5q63Ttr8XOSQ2OpaOgGRBwCBX1IvA4pGQQoCxa1RCbfkteFe8IoxHheNPhQlv9dpJ251HSCmix5snFxRWyv3+TFxrqXJZbLvL6sBCoBC4egSsY9Ywj2w/ljHhvcMJvfcjDntR5/XeD+mRk495A81cVl4bX1ccom0vGlPXKAQKgUKgECgECoFCoBC4NgRKsLg2/OrbhUAhUAgUAnuHAGIfOYH84iUhjJLnvxZGsJBA+/lhJ8OEhrKz90/DJKP2mUceFnJG2JlJwPD+dfU6mAgIEmNrC3LG7lBtExaDGKHNRAc5K4S90iafe3x2GO+SjPn9w/Fcou4XTT7P3BeEDOdqrkO+DpetUggUAjcJApOE2whlnmPWseu6xm4H9k2SYtcO/e2AtwPHbJH0fnzrWneZFC524Op1ikKgECgECoFCoBAoBAqBWUOgBItZ65GqTyFQCBQChcBmCCDAhEIS9kiuB54WzwhDxCPkXxX2kjDkGELf8UiNPwvLpNQ8KuSE8LlwScIuzRKZlnG9eVKkZwhRwnOJRn3+S2EfEvapYR87qT8sFIKN5xKTvjpMGCkJb+Hgnj+9S3XylXooBAqBQmBHEbC+Wm/kHvhA5K+YeeL/W75fzuenlPF6WR4WOzo26mSFQCFQCBQChUAhUAgUAoXAlgiUYLElRHVAIVAIFAKFwIwgkCGgeBPwRpBkE3HP6yAFiF+I58ixZ4Z9WBgPCkyUHA9yP/CyEAP7j8Ik83Se4YyESVJvbSSq8A7hNUJ4IED8Shivkq8PI1IQMeS1UHyuLYScjwgjbigfEyYhKVHGOW+bvL8cXhZr0eZZEmomVauHQqAQ2M8IhHeF6luPeYsRWc95L0SL/dasDWP47bdGVH0LgUKgECgECoFCoBAoBAqB/YhACRb7sdeqzoVAIVAI3LwIEBjs2pWTwj3sZWFIfUIETwoJpjFj7wvjjYCo/wthRA5JPIkAEnRKSu074ma3ZihMEtFCnYRyQvgRIogvwqrIz3E8jIfIdOFBQcyQ5DYTkvvc92ElZBS8fi8MmzhObjpDbV7XnHpZCBQC+xwBIqo113q2X4XRsYBc3hX7fCRW9QuBQqAQKAQKgUKgECgE9iUCJVjsy26rShcChUAhcPMgEMS6xmbCbTt3hYU6GYbAFxoKMYbkJ1TwqTXL7QAAIABJREFUMuCBIGySMFDECu/zxvi5sA8Pk9Da8TwOkGmXZsTDIjt1OnzKxXjTLmWiw2dP2jvd+TwxeFIoBBiCjLbBiSeJpKR3hMHqF8OIGLD0+X4lEqfbX88LgUJg9hCwtliPiKMzHw4KfJXDYvYGUdWoECgECoFCoBAoBAqBQuDmRaAEi5u376vlhUAhUAjsCwRCTFDP0C1GnhAnPNrBm7kpPjKeS7It+TaC3usXhCHuJX1FziPN7g3jhUDQOBUmVJL3ncuxs1JyV7K2nJnUX54OgovPHgh76aSyGWdFPg6eI58Y9uthRBkixydNMIDD3WHw43XxWBgPlH1BJs5Kx1Q9CoFCYEsEMnSfNZVgUaUQKAQKgUKgECgECoFCoBAoBAqBK0KgBIsrgqsOLgQKgUKgELiOCCDCeBAg6QkUd4Uh4HkQyOcgf4NjeF0g5N8d9tDkGO99XBiRYj6Ml0Ym66aGhC7SmiXyPhOHE1MIC9rz22GfM2m30FjeE/JKmCg5LoR7Ili8POz9YQQaoaLgwMPEc9/JXc+z1N6oVpVCoBC4QRCwLhEsrF1VCoFCoBAoBAqBQqAQKAQKgUKgELgiBEqwuCK46uBCoBAoBAqB64wAbwleEoh3YY7kdiA+IPYJEQpvA6GUiBpyQMgHwVuBlwEBw2cIf48EjsGMiRUJMdFCCCehVeSgUGc5OtQbDq8KI9jwNCE++DyLtvLE8MjbAg6OkeOCIRNXhdua0bZPNaWeFgKFwD5CwDpDqHhCrNiHCbf3EdxV1UKgECgECoFCoBAoBAqBQuDGQ6AEixuvT6tFhUAhUAjcUAhM5bBAsvMiIEgQIBD6p8LuCXtGmJBIvC4IFH8SJhm3hNQI+peEIfQl40beEzmQ/u6Ds7oLeDo0FM8SnhR/NGnbZ03a4n3tIt78cRhPCse9Kcz3eZ48GkbQIeAQbBTt52lBEKlSCBQChcBOI1AeXDuNaJ2vECgECoFCoBAoBAqBQqAQuEkQKMHiJunoamYhUAgUAjcAApm7glfFc8J4FxAwCBSZo0HSbUIGQt7xCHlhoISRIlAIA8VDgWiRuStmmVjLxNjaQWzQzheG8brwmtjyzLAPC3tj2C+HfWkYgYaAo63vCBMSy7kk4vYdWFQpBAqBQmBHEZh4U8zymrqj7a2TFQKFQCFQCBQChUAhUAgUAoXAziNQgsXOY1pnLAQKgUKgENg9BIgQRIoPhhEs/jRMMmnvCZuExJerQV4LBP2nhBEneCEQKDIskuOVFAR2r8bbPPMkufj6oyUbJzCICZ/5N7wm0hAmtJnHCUGCB4U2EjdgIrn294e9New1YUJEMRiOM5lXKQQKgUKgECgECoFCoBAoBAqBQqAQKAQKgUJglhAowWKWeqPqUggUAoVAIfAUBCZEPuI+Y6MTH+RlOBGGoOctIH/Fe8MIEbwsfCbk0cdOHoVLQu4LK0XMQOo7VrbtWd8NTFQRAkshXAgL5fXzwwg3QkBpq8+Unw+TdJs3xXsmbfYekcNxQmRlIVzMevunqltPC4FCoBAoBAqBQqAQKAQKgUKgECgECoFC4EZGoASLG7l3q22FQCFQCNx4CCDqeRgI+USkkKdCIVLcFsbDAlHvc/kckP2OJ2zwvOCJoMj9gLzPXBizjFTmsvCoHQQbQsQPTzB4djw+K+wPwn497LlhvE+0UW4LAoXcHWcmeBBtFOcrsWKWe77qVggUAoVAIVAIFAKFQCFQCBQChUAhUAjcZAiUYHGTdXg1txAoBAqBfYxAEvdECGIDAp5AwcOCtwSvCTkqkpBH4iPsCRWOIVzwzBAiiqiB+N8vhL16EldSZEgvk4+YtI13idBQp8IeC3vVpO0w4oEh54Xva3d6VQz3gXfJPh6uVfVC4MZF4NDhI0fvfvozT/Z7vd77Tr333YN+3/papRAoBAqBQqAQKAQKgUKgECgECoFrRqAEi2uGsE5QCBQChUAhsEcIpLjAyyDDG6WIgaT3Ps8KCbaR8oQL4ZNeEUakkMuBwCE01Jj43w+E/VRIrOnQUCAnWhAgJNZ+NIwgcVeYe7uQUNopFNbTJ9jwuMhE474/M/k79mj81GUKgULgGhEIneLY3/uWb/t3n/65X/BF3e7cOLzcpYsXzv+37/3Of/sfv/2f/eN+KBjXeIn6eiFQCBQChUAhUAgUAoVAIVAI3OQIlGBxkw+Aan4hUAgUAvsQAUQ7MULYI4929spZwaPCewfDhEAiYvCseFcYgUO+B+Q+Yj8TT+8XDwvdlHXNhNnaJIm290+Fyc1BkJBsmwcKLIgWRA1tzxwXYw+U/SDWqGeVQqAQmA0EYs1ofdt3ff+PPv9FL/2Y7/iWf/hNv/WWX3rT4sGDh179Wa/9S3/t677x7z3rQ5734X/na/7yX5yN2lYtCoFCoBAoBAqBQqAQKAQKgUKgECgECoFCoBAoBAqBXURAzu0pa8fzA2Enwm4Ne0HYF4e9Nuxzwj4u7Blht4Q9J+xjwp4bdixsLqwbhtzfN2Wq7a14zmBweNKmg/F4R9jxsHvCPjrs5WHPC7s9bHFi85Pvpuixb9pfFS0ECoHri8CnfObnfsFb339+9Gmf8wVfuL4mn/8lX/HXffaaz//CL7u+tayrFwKFQCFQCBQChUAhUAgUAoXAfkegCIv93oNV/0KgECgEbhIEEPZTxf2L9wSTfJtJvE2EkHxb+CNeBZcmzx0nbJKcDpkLYl95GaxrPyhgoL3aphwJAxKPE3h4rv1eJ3j7JhTWdGfX80KgELj+CHzbd//Ajz3v+R/5os95+UcSgZ/infaff+wNv7wYLhdf+ppP+OjrX9uqQSFQCBQChUAhUAgUAoVAIVAI7FcE9tXu0v0KctW7ECgECoFCYMcRQJYJbSReulwOwiNJOi0ckhBInguLhNT3+k/DCBhPxFe/AUIiZf4OggQTAktybSKFNjNhoITQymTd+yJvx46PljphIVAIXDMCz/+ol7zsPe/8g7dvJFY4+c//9I//yHM//P9v7z6gs6i2No5/Si82QHrvAVIIvfcuKE2pCihFEVRAQFSKoNKk9957771LT0ggIUAgoSO9SC/6zYOOdxjeJG8aJvLPWixk5pwzZ34zuWvds+fsndctQcJESkfHDwIIIIAAAggggAACCCAQIQFqWESIjU4IIIAAAjFAwPzCVwvyWrDXzgkFLrRgr10HCk6YgXkt3MfqRfu/i2/b2c17Uros+xfP5i7Kp8f/AwGaGPDKMQUEXl6Bt5IlT/HE+AlJYPHsqRP279qx5cH9ewoi84MAAggggAACCCCAAAIIREiAgEWE2OiEAAIIIPCiBUJasP97od7ccaFpKTihQIUW1sy0STr+dKfBf3Xh3sF9xaaC4i/6deJ6CCAQToFbN29cfztl6jQhdTPiFHcDA/wOhnNYmiOAAAIIIIAAAggggAACzwiQEooXAgEEEEAgVgsokPH3Yr019ZH5FbAZyHhitPnjvxqsiNUPkMkjgECsEDhxNMA/e+68rq8aP7FiwkwSAQQQQAABBBBAAAEEYqUA/4cjVj42Jo0AAgggYBcwAxcKSjj6gxgCCCCAQMQF9u7ctilR4sRJPAoWLRHxUeiJAAIIIIAAAggggAACCIQuQMCCNwQBBBBAAAEEEEAAAQRCFdi2fvVyNShfrVYdqBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQACBf01g/obdh1bt8j8Z3gmkMGpfJEvxdsrw9qM9AggggAACCCCAAAIIvHwCcV6+W+aOEUAAAQQQQAABBBBAILwCSV97/Y2K1d+t67V7x9bzZ087FbgwUvS9MmfNDu+EiRIl3rdz++bwXpP2CCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggMAzAslTpEy1L/jqw/6jp85zlsatQOFiB87c+rMCqaScJaMdAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIhCXQd9TkOQpaKM1TWG11vtWXXbsrYPFW8hRvO9OeNggggAACCCCAAAIIIPByC1B0++V+/tw9AggggAACCCCAAAJOC8yfNnF03Ljx4tVu+NEnznTKnssln9JHXb965XJY7ZMYOafCauPofJy4ceMq9VRE+tIHAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEYqnA4i1eR1bvPnzqVePHfgsKHHzds9+QkdMXrR48cfaSLQdPXtl44MTFgWOnL9Af7dBo/tlXXez93qnX8MO9QVcemEGLN958K1mXHwYMm716u/eQSXOXZTEiH/Y+2XPlyTdq5pK1+4OvPdpy6NTVYqXLV7a20Vx6Dx47NZ9HgcKhUSdJmvS1qOinMV6NEydOl94Dh5euWPUd65hKiTVw3IyFDVu0ae/MY69e+/3G05Zt2r0j4PwtFTrXmCXLV67uTF/aIIAAAggggAACCCAQmwXYYRGbnx5zRwABBBBAAAEEEEDgBQssmjVlfOp06TOWKFepmv3SKq7t4uZR4E/jRwGDN95Klvzu3Tu306TPmCljlmw5smTLmTv526lS2/vldfMsGMfYKvHHH0+eZMicNfuctb/6fNCs1ecJEyVOrMX/MpWq1bT2KVisVNnpyzfvyZw1R65Zk0YPvX/v7t1uPw8ZbW2jQIUCIaHx9Bk6fvq4uSs3RUU/jeGav2CRBsa8rTtQ3v+w5WcKViho0blX/6GV3qldP6Q5KeDx47AJM/Tn5vVrV4f37fnNjs1rV2nMMpWq13rBj5rLIYAAAggggAACCCCAAAIIIIAAAggggAACCCAQcwXeTJY8hXY1/DJ+5qLQZpm/ULGSql9h323gqM9cI0AxdcmGndpZoR0Fm32DLxcuUaa82iroYU35lDZ9xsxb/U5fm7dup6/aq02D5q3b6VqvGwfM8T9u16mbdng42gmiNgocqE/3/sPHW+cU0X4ao0nLtl9pzKat2nXUv/O6exaS1aAJsxZXe69+I+/TN/9QMCIkNwU01EZBDrONgjMas+q79RrG3LeCmSGAAAIIIIAAAggggAACCCCAAAIIIIAAAgggEEUCCYztEZ91+vaHzNlz5g5rSKVi2nPi8v3XjAhBSG0bffzpF1pod7SjwtpHBbm1SN/6q296DBgzbb7SO2XL6ZI3pHF17V+PXPg9XYZMWcw2SjOla1nTO6ndiGkLVzkaRzsZlNpKfewpoyLaT9fRjg2NmT5Tlmy6xpw1Ow7MWrXdK168+PF1fuUuv+Bxc1c8s6PDnJ8CNHJo2/n7PtY5f965+49eJ68/Nkp8vBHWc+E8AggggAACCCCAAAKxXYCUULH9CTJ/BBBAAAEEEEAAAQQiKRA/foIEwybPXd7o48++ePWV52tT2Idfv2LxfPUJra5CPo+ChS+cPXPq6uWLv4U2Pc8iJUprB0WCBAkSVqzxXr1v23/S5MSxAH9HfYqWKldJtSrGD+3X+9yZU8Fmm1z53PKruPed27d/1zHtqnDzLFQ0wM/H29E41YzdCpmz5ch17PAhXz8fr71mm4j2M/vnNuZxKuj4sbOngk/UMQqTq85Gjw5tmj169PCh2hj1weM5mo+R+SpJj4EjJx4/ethv3OB+P1jbFC9bqWqAn6/37d9v3YzkY6Y7AggggAACCCCAAAIxXoCARYx/REwQAQQQQAABBBBAAIHoFdBieb78hYq0blCzYlDgkcNhXW3X1o1r1aZwybIVQmrrWaR4aV+vPTvDGkt1H4zSFU9Ub2LFgtnTft28fnVIfT5s80WnG9euXpk9eexws412hFSs9m7dFQtmTTOPZc2RO48KeAcG+B+0j2WUyojb6suu3XV89ZL5s6znI9pPY8RPkDChanTs27lts4I5Rmqpb+dMGTci8Ij/IZ3XLosURv0O1aawz6lOo2Ytleqqd5f2rczghtokT5EylYIgB/bu2hGWI+cRQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEIjVAmYthyq16jUIz42o1oRSHjnqo8V3pUay1mIIaWylYFLbPccv3UuVJl36kNqlTJ02ndepG0/ad+35s9lGaaGUZmnhpr3+2qVgHq9Vv3EzjZkley4X+3gKDuic/thTT0W0n66Rxy1/QY1Zs36jj+o1adF6m/+Z69aaGpqLzlvnr37aXbJsu0/gxIVrttnnqrHURwW7w/NsaIsAAggggAACCCCAQGwVYIdFbH1yzBsBBBBAAAEEEEAAgSgQaP1V1x5KwbR22YI54RlOOzEyZsmew1Efj0JFS+j4gb07t4c1prEZwlVtlhu7Ky5eOHc2pPZFSpWtqJRNKxfNnaFdEnUbN281d91OH7X/rHHtKvfu3r1j9s2WyyWvdiqcPnki0DqekZEp3iftvv5Wx4wMSzfsu0ki2k/j5crr5qG/Aw76eDX+pO1XU0YP6W9c4rp1TvrvoONHA6xzUlqtDJmzZp81YdQQ+72XKFepmo757A97p0pYzpxHAAEEEEAAAQQQQCA2CBCwiA1PiTkigAACCCCAAAIIIBANAqqxoF0GS+dMnxTe4a8YtSm0q0FBAHtfV8/CRVVzQTUZQhv3jTffSpYiZeo0ajPXSJ8UWlvVurh65dJFpUhauu3Ase/6Dh27c8uGtQ2rlvS0Bzp0T2dPBp948vjxY+uYtd5v3CxZihQpr1z67YJqV/xp/FjPR7Sfxsjpks/twf1791RwW/c1Z/KYf9JW6bzSTenvY4f9fK3XrPpu/YZKc7V53cql1uNyLVa6QmXV6girDkh4nx3tEUAAAQQQQAABBBCIqQIELGLqk2FeCCCAAAIIIIAAAghEs0A+jwKFdQn/gwf2h/dSCRMlSvzH058nT+x9VfD6oNfeXfaAgL1d9tx5n+6uCDjk42XWeghpHh4Fi5ZQTYc+Q8dPV4Dik/rVy3b+9KP3rbsYzL5KFWXfXaEaEtpdsWDG5LFvvJUs+SHvvbvt14poP42TM08+96DAo4cbNGv1+fTxIwbdvXPntnV8o7zF010fwYH/22GhdFAlylasum3jmhWq42FtX6JcxapKKeXL7orwvpq0RwABBBBAAAEEEIjFAgQsYvHDY+oIIIAAAggggAACCERG4K0Ub6dU/2vGzoXwjpMxc7bsly9eOK+QhbWvik9r8d7PZ//esMbMldf1aRqltcsWzg2rrepb+Pt672tas1yRj+tWLe21e8fWkPq8bdS7MGIap63n6zZp3lqBiu2b1q5U8OKg977nAhYR7afrKPhibIqI7+KWv8C8qeNG2uemdFMnjgb4W4tqZ8ySLYfm5LXr+XupXLPuBwr4OAqshGXFeQQQQAABBBBAAAEEYqsAAYvY+uSYNwIIIIAAAggggAACkRS4bxR+0BDJkv8VuHD2J5kR6DBSILlrF4W9T9YcuVyUzuiwUcshrPFy53XPrzab1ixfHFrb+PETJFD6qX07t21WKqfQ2iYwtn4kSZr0tauXLv5mtkuS9LXXW33R5ftZk0YNTZ0mXQYdP3My6Lh1nIj20xgqCK7dEDmMoMWC6RPH3Ll9+3fr2PLIlDV7ziN+vt7W4+YOk8Ajfgetx1OnTZ/B4PXUDgxHgZWwXDmPAAIIIIAAAggggEBsFSBgEVufHPNGAAEEEEAAAQQQQCCSAmZ6IrO4s7PDKe2RCl+rALa9jxGweFqrwV7Q2tHYqkehwIE9eGBv+7pRE0LHHj188CCsOSZOkiSp2ty9e/uflEytvuzy/R9//vHHlFFD+mfN+VctCWNzyDMFviPaT2Nl/7tw+OPHjx7Nnjz2mdoVOq+dFApa2Gt6pDVyUDmaS7uuPX8+f/b0yYcP7t+317wI6/45jwACCCCAAAIIIIBAbBYgYBGbnx5zRwABBBBAAAEEEEAgEgJ7d27bpHoQDZq3aZc5e87czgyVK6+bx0efftk54JCv93aj9oK9T9r0mTLrmLVQdO587vm1Q8LaVmmZshi7MbRrIqzr3r3z+9MdC9oFEVbbBEZKKrUx1vrv6W9du/HHn305om+vbneMSuCqU3HzxvVrKpBtHSui/TSGipfr781rVixRQW/7HJUOSseCjh05bD2XOOlrr+nfRpzjkXncrUDhYkqpdc8ogqFdKgqC6NyrceLECeveOY8AAggggAACCCCAQGwXIGAR258g80cAAQQQQAABBBBAIIICKvT8w9eff5IwYcJEE+av2lKoeOlyoQ2V192z0KgZi9c+efzkca+v235sr1+hvtp5ob8TJU76dKdDjTofNJm1aptXgaIly1jHVrBCuw5UcDus6auAtQIBZgols71SPzVv26FrMyOAYh7TQr/530aWpmT9Rk2ZeyzAz3fpvBmTdfw1I3fTJSNIY79mRPtpHDMgsXj21AmO7kUFt3XcuIVz1vM3b1y7pn+nzfBXkOftVGnS9h0xefbgPt99rcCFr9eenapxoWfTf/TUeWE5cR4BBBBAAAEEEEAAgdgu8PT/TPCDAAIIIIAAAggggAACL6fAzq0b17Zv/n7NPkPGTRs3d8Um7XjYuGrZwgA/H+9rVy5fMuIPcdNnypKtYo336tWs2/DD+8bOha5tmzU46n/Qx5HYqaDAYzreqcfPg65evnSxYfPW7XZsWrfq183rV1vbaxeB/u27f89OZ+RXL10wWzslFKDQtfMXLlayXuMWrVU7opcRdDHHuGVsn9AOivc//OSzD1u376QgQIdPGtVWAWu1eeXVV181Skzcsl8zov00TpbsuVxOB58I3L1983pH95It5187LG5cu3rFet4otr1F8/q6V7+hG1ctXdi0ZbsOm9euWGLsxPBXXYzfjUlNW7pxlzHlVwf07PqlM060QQABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAgVgto50GbDt/0XLXL/+SBM7f+tP/ZHXjxrr7yV0ql0G5UuyamLF7/q/p7n775R9+Rk2YbmZwS2/t89V2fAYu3eB1RYWln4FToe/kO3+PmvLxOXn88eOLsJS6u7p72/u2/6dVX7bYfPnujeJkKVaznfxw2Ycb+4GuPlNoqqvrNXLl1X5lK1WuFdB+TF63bsW7/0Wd2V5htW7bv/J2cNN8+Q8dPV+qnspVrvKt/6x77jpo8R0XDnTGiDQIIIIAAAggggAACCCCAAAIIIIAAAggggAAC/ykBBSVKVahSo0bdBk0rvVO7fv5CxUqaRamdvVEFGJSyKaT2BYuVKmvWfnB2TNW9UL9ipctX1vgh9dOOBAUkHC30614GTZi1OHmKlKns/SPaL6z5K61TqjTp0ofUTrtAcrjkc9N57RgZO3vZBq9TN57Ua9KidVhjcx4BBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQiFKBfB4FCq/c5Res3RWLNu17pkB3lF6IwRBAAAEEEEAAAQQQiKECFN2OoQ+GaSGAAAIIIIAAAggggMDLI9CwRZv2kxat3X5g764dp4KOHzvsRDHyl0eHO0UAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAIFoFVDarAFjps1XvYomLdt+FT9+ggT7gq8+bPTxp19E64UZHAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBCQQMYs2XIs3rw/YLNv8OVCxUuX0zEXV48CSgnlUahoCZQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAgWgVyJI9l8sG78ALy389eCJ9pizZzIs1aN66nXZbJEyUKHG0ToDBEUAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBA4OUWSJQ4cZJl230CNxw4/lu6DJmyWDX6j546b/bq7d4vtxB3jwACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAtEu0KbDNz2V9qlMpeq1rBd7NU6cOFv9Tl/r2mfgiGifBBdAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQACBl1tAaaBUu8KuULhEmfJ/BTKq1Xy5hbh7BBBAAAEEEEAAgZdV4NWX9ca5bwQQQAABBBBAAAEEEEDgRQvEjRsvntJABR7xP2S/du2GH31y7+7dO7u3b9nwoufF9RBAAAEEEEAAAQQQiAkCBCxiwlNgDggggAACCCCAAAIIIPBSCDx58vjxwwf377/+xptvWW/YxdXds/I7td9fuWjOjAf37917KTC4SQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEPj3BAaOnb5gb9CVB55FSpROmChR4uJlKlRZt//oud2BF++mz5Ql2783M66MAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACL41AqjTp0q/YeShI9SrMP16nbjypVb9xs5cGgRtFAAEEEEAAAQQQQMCBwCuoIIAAAggggAACCCCAAAIIvFiBpK+9/oZqVri4enjevH7t6rL5M6YEHPL1frGz4GoIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggEAEBN54K1nyCHR7IV1Sp02fISoulCBhokSZs+fMHRVjRXSMN958K1l23e9lAAAgAElEQVQOl3xumbPlyPWK8RPRceiHAAIIIIAAAggggAACCCCAAAIIIIAAAggggMB/TiCvu2ehA2du/VmmUvVaMe3mPIuUKK25FSpeulxk59Z35KTZExeu2RbZccLb/9U4ceLUbvjRJ7NXb/f2Pn3zD92P/sxcuXWfgijhHe9Ftp++fPOez77+rveLvCbXQgABBBBAIDoEXo2OQRkTAQQQQAABBBBAAAEEEEAAAQSiVsA1f8EiGvHRwwcPonbkyI9WtvJfQRQFLiIzWj6PAoWr1KrX4P7du3ciM054+6ZOlz7jtKUbd33fb9i4ixfOnendpX2rDp80qn06+ERgHrf8BXPnc8sf3jFfVPvXje0gcmMnyIsS5zoIIIAAAtEpEDc6B2dsBBBAAAEEEEAAAQQQQAABBBCIGgGlKNJI/r7e+6JmxKgbJX/h4qU0mluBwsUiM+rnnbv/qP63f791KzLjhKdv+oyZs2pHx5/GT/M6lUv67t+z0+yfJUcul7Zff9/n3OlTweEZ80W2zZXXzUPXO3E0wP9FXpdrIYAAAgggEB0C7LCIDlXGRAABBBBAAAEEEEAAAQQQiHECSZImfa1B89bt4sSN+8/He8lTpEyVKWv2nDFusg4mlDOPq/u5M6eCb964fi0mzdfIlpTY3IEQmS/9CxYrVbZIqXIVdW9379z+/UXco96JYVPmr/jjyR9Pmr1Xqbg1WKHrexQsWmLz2hVLrlz67cKLmE9ErpErr+tfAYtjRwhYRASQPggggAACCCCAAAIIIIAAAggggAACCCCAwIsWqPRO7fqqSdDqy67ddW3VLFi4aa9/r0GjJ7/ouYT3eprr7sCLd/uNmjI3vH2ju33hEmXKy3XFzkNB+jtL9lwuEbnm1CUbdpp1Izp2/3lQRMYIb5/u/YeP33P80j1zl4K1v4urRwGZZ8icNXt4x32R7XsPHjt1f/C1R/HixY//Iq/LtRBAAAEEEIgOAXZYRIcqYyKAAAIIIIAAAggggAACCMQ4gS1rVy49eyr4RIu2X3VNmTptuvc+aNpCi+tzJo8ZHuMma5tQVmOeKvx8+OCB/TFtrp5Fij+tW7FwxqSx+tvNs1DR8M6xeNmKVZVO6oif7wH1vXM7+lNC6Xoqsj1mcN9eR/0P+ljnHD9+ggQ9B46cONY4d+Zk0PHw3s+LbO/i5lHgZFDg0UePHj58kdflWggggAACCESHAAGL6FBlTAQQQAABBBBAAAEEEEAAgRgnoAXdcUP79dbCf+de/YaqXsKy+TOnnA4OOq46BjFuwpYJ5XZ199Q/Y2LAIn+hYiXv37t3d9m8mVM0x4jUsWjToVvPP4yfuVPHj9QYd25Hf0qoL7/t3f9U0PFj08YOG2h/9t/2HTLmxrWrV6aOGTogJr8XSseVJVvO3McO+/nG5HkyNwQQQAABBJwVoOi2s1K0QwABBBBAAAEEEEAAAQQQiNUCSqt08/q1qw8fPnhQofq7dXUz79Rp0PTd95s012J51cIuGS5fvHA+Jt5kHtf8BVQU2ghYeMWk+cWNGy+eW4EixQ4fOuB19cqli9rBojoW4ZljiXKVqrnmL1hk/YrF8y+eP3vmr4DF79FadNuzSInSCrR0bdui4ZPHjx9b59uyfefvipQsW7FR9dIF9F6E515edFulstJ7be5MedHX53oIIIAAAghEtQABi6gWZTwEEEAAAQQQQAABBBBAAIEYJ1CsdPnKX/fsNyRLjlwuDx/cv68JaqFaX9f/dv7cmUMH9u2JqcEKzVX1FLQbILoX8sP74FyMnR/6yv+Q977d6nvQ+LtKzTofaBfLA2PbhTPjaXeFgjHjh/bvbdaLiO4dFo0/+exLBVfWr1g0zzrHek1atP64XcduLepWLX3tyuVLzsz/32yT192zkK5vBCy8/815cG0EEEAAAQSiSoCUUFElyTgIIIAAAggggAACCCCAAAIxUkD1CIZNnb/itFGL4MNa5YueNf7j7p07t+PEjRtXX9DPmzZ+VMAhnyjfuVCgaMkyedzyF4wsir6gz53PPb+/r/e+yI4V1f21U0FjHvTau0t/K/AjVwUynLlWyfKVq2tHxqY1yxcHHvE/lChx4iTqd//enTvO9I9Im1Rp0qUvW6l6rblTx4207qCoXvv9xp1/6D+sy2fNG8TE1FuO7jWm7ryJyHOhDwIIIIAAAggggAACCCCAAAIIIIAAAggg8FIImAvhSvezL/jqw5x5XN1nrty6z/v0zT9q1W/cLKoR3mvw4ccHztz6c7Nv8OXIjp09V558GqtB89btIjJWipSp0yRL8XbKiPQNq8+QSXOXaW66htoq+KB/awdDWH11fvryzXv0DHLkzuuqf9dt3LyV+hcuUaa8M/0j0qb1V9/02Bt05cHrb7z5ltlfacH0XkTluxCd7ua8F27a679kq/fRiDj82320Mydjlmw5/u15cH0EEEAAAQQQQAABBBBAAAEEEEAAAQQQQOCFC7xmrFDvOX7pnoot6+Kp06bPsN7r2Hmvk9cfm6mIompSLT7v+I0W3ictWrs9smNqMV1juXoWKhresV4xfpZt9wn8rNO3P4S3b1jtNfZWv9PXVuw8FGS2VU0LGf88YtKssPprd4Xuq//oqf+kZVKg4+m9GjUtwuofkfOvGj+rdvmfHDhuxkKzf6svu3bfH3ztUY06HzSJyJiO+kSnu3k9Lfh7nbrx5MdhE2ZE1bxf5Dg9BoyYMHHhmm0v8ppcCwEEEEAAAQQQQAABBBBAAAEEEEAAAQQQiBECWqyu9E7t+vHixY9vTkhFi7/58ZeRiZMkSRqVk9SCdbacLnmt14ro+N1+GjRKC+rxEyRMGN4x3AoULqYAQIVqteqEt29Y7bUrQmP3GTp+urXtlMXrf1WQJKz+2l2hBfesOXLnMdt+3K5TN42pXSVh9Y/I+SKlylXU+OWqvPNe8hQpUw2ZNGfpjoBzN4uXrVg1IuOF1Cc63c1rKoAVmZ03UXm/4R1Ladrk3uWHAcPC25f2CCCAAAL/bQFqWPy3ny93hwACCCCAAAIIIIAAAggg8LeA6hWsX7F4/qNHDx+aKEf9D/r8/G3HtqppEZVQKiJ94liAv/VaER0/r3uBQsZQB81i4eEZp2ip8pXU3nvvzkjv9LBft0DREmV0zGf/7l+t5w56792lHStGxqVkIc21RLlK1ZQ+as3SBbODAo8cNtslSJDgaVDmnvFAwnOfzratWbfhhzdvXL+mgNLCzfsOlzFqWVy9fOlihkxZs0VFcMmcR3S6m9fIndc9v/7b78D+Pc7ef0xpl8/YQZMk6WuvR8d7GVPukXkggAACCERMgIBFxNzohQACCCCAAAIIIIAAAggggIBDAS18hyd9U2g7J/Qles48+dz9ffbvjQh39lwu+c4bVcavX70S6Voa9uvnL1y8lI757ns2YOH7dwHuvO6ehUKas+pIPHn8+PGYQT/1tLZJYOQ50r/v37t3NyL3G1ofOZc1dlZsWLlkgYIlwYFHA3ZsWrfqxrWrV7r2GThi6tKNu95MljxFaGPovHZPpE6XPmNo7aLT3bxu7nxu+R8+fPDgqP8hn/BYOXsP4RnT3lYBIRVfD2kMcweNnxPvtQIbEZ2LUpRFtC/9EEAAAQQQQAABBBBAAAEEEEAAAQQQQACBGCHwapw4cbr0Hji8dMWq71gnpNRKqn/QsEWb9iFNtGnLzzsoVY/STYXURou5n7T7+tsN3oEX1Hb26u3ejhbLVctB563FoJXKqE2Hb3qqBkCpClVqWK+hheKve/YbMnL6otWDJ85esuXgySsbD5y4OHDs9AX603fU5DnNP/uqS1Qgq/7HNv8z13VN63hvp0qTVnNWgXNH19HuCp3v3n/4ePt5BQ50LjwpuvSMhk6et3z41AUrzeLdjq5bplK1mhrbUfonjaH0VL+Mn7koJJvmbTt0VWoujaE/eg9UR0Lto8r9reQp3laNlYkLVm/9tGO3XqE9JxWNV1ottUn+dqrUSh2mmimfd+7+Y0i7RUK7h5CuVb32+42nLdu0e0fA+Vuq/6HfC9UfcdReu2r0XH89cuH3PScu39c7brZ774OmLUbOWLxGhdoXb/E6omLr5nupOiZ69vbnrqLcGkfvjMbR7+WHrdt3mmYEl3Sv2iFjn4fa6D7X7T96Ts900IRZi+0ehYqXLvftz0PGhOarudjf7aj4vWEMBBBAAIHQBUKMdgOHAAIIIIAAAggggAACCCCAwMsqoEBBg2atPk+dNl2GbRvWrJDD+x+2/Ez1LvTfClxcuXTxglJM2Y0uXfztvI6lz5g5q1JO2c9r18SQyXOXFS1VrtKmNcsX37x+7WqdRs1aftiqXcdhfXt+Y22f19gJoH8f+jvtj0ehoiUGT5i9RMENpZ2qZRTkbt2gZoX9u7ZvUTstoLu4eRS4e/v271psfeOtZMmNDRZBadJnzBTPWLVVnysXL16I7HNNnylLthQpU6fRDgWNaR3v8sUL5387d/a0OXf7tT7t+G0v7QwYN6Tfc4XAjYxQT1NCObPDQl/Pf/vz4NHvNfjwY/MaSiXV+dOP3nd0f1rcvnP791v7ft22yX5ez3jVorkz3qnX8EMFmuzPzcXV3bNdlx4/HfE7eGDz2hVLyld9p7begcMHD+yfNOKXn6PCXc9WC/gKPmh+nkVKlF67bNFca8osc95alNcujkWzp03InD1n7vFzV2zSs1Zqs/yFipU0NvnEH9znu6+t9xnWPdhNdI3eg8dOVcBCz3m48W5my5U7r34vjHhbPB2z9klp/LJMmL9qi96L5QtmTnXJ5+H5qVHsfeXiOTMunD1zSjtT1O/u7d9/V1DrlpGaK3W6DBn1Xr5i1JdJnCTpc3VkFIDS74veMRkrMFW4RJnyeqdTpkqdtn7Tj9tsXb9qmTkPvRMDx01fULpitZr63fzz//78s0rNuh9UrlXng5UL5/xTa6XZp192tr+31nvJnc89v+7lm89bNNq+ce3KyP6+0B8BBBBAAAEEEEAAAQQQQAABBBBAAAEEEIiwQJOWbb/SV/RNjSCCBlF6I31dr6+1q71Xv5G+Dv9x2IQZji6ghWz11UKyo/O9Bo2erP5V363X0DyvxdE9xy/ds6eH+nnEpFnbD5+9oeCDFm/15fqcNTsOqFB1zjyu7rpOv1FT5jq6jhaudd6+SyTCKJaO2vGhsfUlu6Px+o6cNFs7O+znTBvtAnHU76fhE2fuC776T42RkOaqhWl9qa85jJ29bEMOl3xu+vJ/k0/Qpbadv+/jqJ++uNe8QhpTu1U0XvuuPX+2t+ncq/9QndNCu84lSpw4idwd2UbEXYvwu45dvKPnq4CAgl163/Re6N7s88liRCs0n7qNm7fSboUlW72Pqo/mJYPdgRfvKuBg7Reee1A/tdd7qkCdOU7BYqXK6rrWd1fn9Dy020O7MLTYr2NmUfbyVWvWts5Du4v0rnf4/seBYb2Lek/2Bl15YMQyXlOBdK+T1x83/uSzL/X7oHs1U4iZ43Tq0Xew5le74Uef6JjaaZeR7sVso7nuPPrb7ZB2SRmxk1fnrd91ULszUqdNnyGsOXIeAQQQQAABBBBAAAEEEEAAAQQQQAABBBCIVoE+Q8dP18KndhJo4VdBglmrtnuZqWVW7vILHmd81e5oEkrJsyPg3E1H6WTMBXv7ori+PjeDI9YxV+w8FDR61tJ1+rp86bYDxxZv3h/wupF3x2yjRW6l63E0j0Yff/qF7sH8Yj8qwXoMHDlRY2tXgKNxtRis8+kyZMpintdC8MJNe/21KJ8sxdspHfVTSiadD2uu3/UdOlbjK62PxlV7BSp0TIvN9v5a9Nc5fW0f0tiak9oobZG9jYIjCiCENS+dD6+7Alt6Xzb7Bl8204gpcKXFec1H74z9uhVrvFdP5waMmTZ/q9/pa2mNaIXZZsS0hat0TjsdrP3Ccw8KoChYYQ/+6N3WvIyyEm9Yx27xecdvdM1K79Subx4305kpFZe1rRloq1KrXoOwPBds3OM3ft7KzR981KqtPchn7+tesEhxtTF3QZnnFbzp0P2nX8x/63dNc1UdE0fX144SnZdjWPPjPAIIIIBA1AtQdDvqTRkRAQQQQAABBBBAAAEEEEAglguooPGpoOPHzp4KPlHH+FpbRYJ7dGjT7NGjh0+//ldqm5BuUQW3/Q7s32tPOaPUNp169h1y8cK5s+OG9utt7X/QKFQ9fdzwfxZVdU4L6FrwP3Rg357PO/f40fi4P33HVk3q3rp547rZV+l0jCxHNx3NJZ9HwcJKxXP18sXfovpxeBQsWuLhg/v3/X289zkaW/ej49bi4zXqNmiqnSGzJo0aeu3K5UuO+ikllMYNbb764l87C5Ti56duX336h/Gjr/arvfd+I/XbuWXDcwGH4mUqVPnjyZMnO7duWBvS2GZhcuPD/edSEyl9ka5h7rAIbX7hcTfW/d8cMnHOUu0FaNPo3UpmKqrqxi4eBcpUmHzPji0b7dfTDgsdK1O5eq0+Xb9orcLqZpvbt2/d0n/f/v3mM++Fs/egnQsKSB0/ethv3OBn03YVL1upaoCfr7f1nVPdihZtO37z6+b1q60p0nL9vdMiMMD/kHX+ZqDgkPdeh4E2s63SnmXL6ZJXKbHade3x05TRQ/qvWbogxB0yX3br3V/PcOhP3f+p0aJgkHZhBAb4/RPEci9QpLjehWMB/s8FtmTe8osu32sOC2dOHhfVvzeMhwACCCAQtgABi7CNaIEAAggggAACCCCAAAIIIPASCejr9izZcubet3PbZgUZPm7X6ds5U8aNCDzy18KrdlmkMOoMqPaEnUULnlqwPuj914K99Ue1FpRiZuSA3t85U6NBX6irv+pRKE3QyP69v7PWM9BYWkQ/HXw80NHj8SxSvLSv156dUf3otJCcOVuOXKqrYQZw7Nc46n/IR4EHY3G4mM5p0fizTt/1VrBl6uihA0Kak8Gd8EEoAQt9Hd+5V7+hunbPTm0/NoNCStNl7ubY62CBv0ipchX9fb33GbGdGyFdW2M9fqw7evDA3mbPjs0bdMxe5Dyy7korlilr9pzffdGyqRms0DukHQsaWzUyHAWksub4K2Cxb+f2zfY6KkmTvv667sH+jjl7D6qnoh0bvbu0b2V9vir2rkDegb27dljvu26TFq2VsmnUwD7dzeN63qrJ4r3n123WYIrOqzbHlUu/XbAft1uagQ3Vo7h6+dLFMb/81COkZ6f3Qrt9po4ZOkB1PMx2KvyuuiVb1q40gkJ//bgbbRWMdBQYq1HngyZ6t2VO7Yqo/l8OxkMAAQScEyBg4ZwTrRBAAAEEEEAAAQQQQAABBF4SARUz1qKxgg613m/cLEnS114bN6TvPwWizTRRZ04GHbeTaCdG4iRJkvrsfz5QoKCDghxrly6c4wxlPiNgoUV0FYs+YXwOPnPS6H/y8Kt/Dpe8T2sbHDvs52sfTwvOqdKkS29fXHbmumG10RfqaqPF6JDaauHf+BB/n9L0qI1qgijAogXlkHaEqN1fOyweONxhoeCMUkHdv3//XjejGLKuoT56Vq3+/ipeXmaBcnNuCjCprsTu7ZvWh3ZvGl/1DRzNb+PqZYsU7KhnLM6HNkZ43CvXrPO+AiDzpo0ftWXd/xbUtWieIXPW7LrOQe99DnchZMme82nAYsygn3ra56OA0rlTJ4Psx525B6Uxe5p+ae/O7Yds1y5ermJVnffZ92zAQvVM1FbBFV1T6cvM4uF9v+v0uX0enoWLl3LmvVTqKPXVezO8X69ujgJJ5tiagwIQi2dPnWAea/3VNz2U3mlAjy5fWgNVedw8C5rBR+vc9OzbdOj21HP3tk3rzfcrrN8HziOAAAIIRK0AAYuo9WQ0BBBAAAEEEEAAAQQQQACBWC5g1hEIOOjj1fiTtl8pFY01DVO2XC55dYtBx48G2G9VX3pr0dxMiWSe126JLMZX8cvmz5wS2sKrdTxXj78CFlr07/f91+2UxsZ63izGfOzwoecCFmZtiQPGwnNUPw59oa4xvfeEPrYWsXPlcfVQgKf5Zx26Kg3U7Emjh4U2n9B2WDRs3rqdCjkP6NH5CyMD0j8L8nUbNW+lBX7tKDh35lSwfReFvtTXIvrubZtDDViYtUH09b99jhp7zpSxI1xcPQpot0ZI9+Csu4JaHbv/NOjkicCjv/zw7dPC7vrR7p5PO3zby9wdEeDn422/loIGmbLmyBkceDTAHlRQ24xZsuU4duR/KZDM/s7cQ8nylavLctaEUc8VRS9RrlI1jWUNxqVJnyGTdoisXDT3aQF61b6Yu3anT6Hipcp1bNmojj0wkDJ12nTqo4BIWO+lnrXayGjjqqULQ2tfrEyFyts2rFmhZ6/5j5y+aHWbDt/0HDWgz/dL582YbPaVe+p06TMav7p+9vHe/aBJc7MWSHTsTArrfjmPAAIIIPCXAAEL3gQEEEAAAQQQQAABBBBAAAEELAI5jQLNyqejhXbl558zecxwK5DqMOjfjnY2uOUvVFS7Iexf6ZerWrO2+qxbvmieM9halM7rUaCQCkpvWLlkgaMFXiO9v5vqN6jWgH1MV8/CRTUHR+ecuX5obRRAUW2FsBZ1tZiu3Q+DJsxarJRBk0b+8vO9u3fvhDa2dlgoJ5O9jQqHtzEW8gMO+Xor6GOeV/HnTzt266UaBefPnjp5/O+0Xdb+BYqWLKM0Qb4O0nRZ2+l5699KF+RojtPHDv9F6YVafPZV15DuwVn3Vl927a7F+yE/ft/ZmpqoaavPO2hBf+v6lct0jeNHDj9T/0HHUqVNl0EBmD2/bn2utoXuQXUxHL2b6hvWPVR9t37DG9euXtls2fGhftp9UKx0hcoKCFlroii9k87fM4AnLlyzbeyc5Rv1u9O4RtlCu41sVc+/l4WK6pjv/t2/hvUeGoHBfGoz1wgU2evBWPtqB4YCDXpuvQePnbpki9eRPG75C3b4pFHt8cP697G21e+ufrdOBQUetR7X/SkNl2rW6HhIO1vCmjPnEUAAAQQiL0DAIvKGjIAAAggggAACCCCAAAIIIPAfEsiZJ5+7sZ55WCmcpo8fMciaE1+3aZS3yKvc/vrC3X7bWsz32ff8YmyRkmUr6OtvM21OWFyZjYtoMV6BAaXDcdQ+p4ur++ngE4GO6mG4GYW/tcsjtIXesObg6LzSJimljgovhxV88P278La+lL/02/lz86dPGhPWNeMnTJjQyPT0NNWT9eejNu07Kegx9OfuXaz39GnHb3u9lTzF26ON+gYyc/RMPIuWKK30XrIM7frmF/2qv+GonZ7fvKnjRxU2nqW5u8Xezhl3zVfv1gEjtdLW9aueBib0o4V3Fa/WcaMu+2ndp3YX2K+RMUv2HDrm6F4LFS9dTueMou97wnsPWsgvUbZi1W0b16yw7+YpYaSD0g4UX1uqMxVf13V6DRo9WQGYHh0+bd6gWilPBe0cXV8+em+MGNtzu4Ks7RVAMNJe5dbv2eol82eF9tzc/56DUWumW9kqNd6dOGLgT++UcMu2ee2KJfZ+6TJkzqJj+r2xnnuvQdMWbxoP5tct69fomkeMwFhY7yrnEUAAAQSiR4CARfS4MioCCCCAAAIIIIAAAggggEAsFchuLLAb66XxXdzyF5g3ddxI+20oJdSJowH+9oLTqh2gdDw+tq/HtfiqIIhSKGlHhDMs+fIXKKx2KxfPneGoVoaKgSsVzxEjcGAfT2mFdD0/n/17nblWeNpoUV9f9zuTakqplX47f/aMxp8wbOCPjoocPzd348Ye/V2bwjynND51G7dorQDMnu1/Fb/Wj77ub2CkidKulWtGVWbtRtEOAOuY2uHh5lm4mKMgkv3aqq2g4I+jNEtm21mTxgzTYv57HzRtEVH39z9s+ZmKUo8f0q+3OYaCBT0HjpwUL368+Er/lTufe37tZNBuBft1zLRFjlJXqSaG+jiqoRLWPejdfeOtZMm9jDiK/ZqVa9b94Gl9EO+9z9TUUJ0U7cjo1KpJ3XdLeeTQ7hd7sMM6lqsRsAg4dMArtDZqnzVn7jz6vdmzfcsGo077tdDe0VRp0qbX+UG9v+1UpVCu9KMG/thdO2Ec9UmZOk06Hb9w7sxp87x+X1p+0fl77aRS0OhpwXgHhdfD83tCWwQQQACBiAsQsIi4HT0RQAABBBBAAAEEEEAAAQT+YwL6SlxfkmthfsH0iWPu3L79u/UWtYgaUqBAX4+rra9th0XaDBkzq99522J6aHSqeaHzmoOjdtly5c6rxfiAQ8/XOMhq1MrQ9Q4bNTii+vGoHoTG9NodcsFt6zWNQMEOfc2+ZM60ic7MRQWy7TshylerVUdBiwUzJ401x1Daox8Gj5ly8fy5M326ftHa3B1hGJ+0XkfpvbQzwx5Ess9FASB9na9UTKEtVitIoFRHpStWfcc+hrPu79Rr+KECK9aUSQq8qDbG0J+6dznqf9DHyFzkev7M6WfuxbyeEVNIof9WoMA6BwXMVINix6Z1q0ILDoV0DwrUabxAW/0LLeK75HP3VFDFnirJyJiWXPVEVNDbmWCcnpMz72XuvG75NZdNa5YvDuu90RzUZt60CaPsu6HsfZO9nTKV3q+b169dNc+pIHySpK+9Nm3c8F9y5XHzcBQgDGsOnEcAAQQQiDoBAhZRZ8lICCCAAAIIIIAAAggggAACsVwgu7FQrFt4bHzlP3vy2GdqV+i4vkJXMMBRbQj3AkWKX71y6aK1ILT6KAWQ/r7soJhzSFz5PAoW1sKyn4+Xw10SOXLnc1Nf1W6wj2EsnD+tsREUeORwVD+OvO6ehfSlvY+RtsiZsft+36ndR+9VLG7fjRJSX6WcMjYwPJO6qVT5KjW0GL513V/pkxSo6Td66lzjY/kMXT9v3lCpmvRcdM7IPPV0R4f5k79wsVL6mt++M8B+/ep1PmhiLFq/PmfKuBFh3Zd2a6hWhHZJWNs6454ley4Xo9xC1rNsjBYAAAz1SURBVC1rVy41U1spjVPH73/6ZfvGtStnGsWuFZxRzQ5zd4p9PsaGgKfXvXfvzjP1QOoZu1AU8LHW+AjpXhzdg1EaI5PaX7xw/qy1X7uuPX8+b7zUCoLYa2O8bkQLnN2NoGCg0pw5815qh4nmsHPLhjVhPQ/NQW0eObErQrZGRqrb5pgpjC0XSsM1YdiApzuAVJD7opGPK6xrch4BBBBAIPoECFhEny0jI4AAAggggAACCCCAAAIIxDKB7LnyPC30u3nNiiWOUu4oHZTOBx17PhigdDdKW2S/ZX2ZrmOJjFRK9nOZs+XIpcVp63F97Z/DKKitdDgh1aAwaygcPxrwXMHttOkzZdZ41uLIWgBOlDhxksg+DgUsVJ8grDQ95nX0Jbt9J0Boc4hjRCzsNSzyuHsW1C4NIy5xXZbf9B44oljp8pV/6d2to+ltpCbKoHHtxc7zFypW8pgR1FGqI7Ootv36Wkjv8P2PA7cYhabtqaP0bLSjxtrnFSP1lAIo9rRGzrjncc9fUGMd+rvGRDajcvqAsdMXGCmKTn3/ZasPdS6VUXXb0b2YczDv0RowUXH4pq3bdTx5/NgR7bCwztfZe0hs7DJQP6u/W4HCxZReTEW1tTNCgTy1UdBIfxtr/78b8ZNnAjchPV/tNLK/l0pvpbRS9j658rp66Jk7EzzQHNTfDOSE9n4p/ZM1zVbXPgNHXDOCjAoUmfUtnLlmZH+P6I8AAgggELIAAQveDgQQQAABBBBAAAEEEEAAAQT+FjADEotnT53gCEUFt3Xc2PxwznpeX7a75i9UxFyItp47czL4hP6tmgvW4/r3nDU7Drz7QZPm1uNaINYujv27tm8J6cGojRZeLxufw9vbaJeCjiVKnDSp/q5h7B6YtWqbV4GiJctE5kFrsTerkavIe49z6aAici0FJIwNFs/ssFAKJAU9dO67vkPH1mv6cRulyppt1JMwr2HEeBLov+/e+f2ZFF7GDouS/r7e+8bNXblp+JT5KxQMss5Li/lDJs1Zaix63+7T5YvW9jl3+2nQqCmL1/+aLMXbKXVOX+TXafRRS1+vPTvtu0accf8nndP1q1dy5XXzmDB/1RbdV7tm9d8xg0Dmvdz5eyHePqdTQceP6ZiZwkm1O3oMHDlRqcyG/PR9Z3tqJmfv4eaNa09rRaTN8FfA622jOETfEZNnD+7z3dcKXOieFfjRnPuPnjpPbTQX7W6xumo+euc0J+vcFYyyvpdKDzV7zQ7vhi3atLffo+5NtS6ceYfsHmYfBat6Dx47VbsmzGP3je0V5n+r8HkFI93YLz9066hnqTRjOnfJtsPEmTnQBgEEEEAAAQQQQAABBBBAAAEEEEAAAQQQiHKBacs27V667cAxc1eE/QIDxkybf+DMrT+Tp0iZynpOOyV0vP03vfrOWrXdy17jYOSMxWt0Xl90Fy9TocrH7Tp12x148e6GA8d/0yK4dSwVZVZbLWiHdIObfIIubTl48pkaBmbbqu/Wa6j+P4+YNKtTj76DvU5efzzMWKwP6Z6cRczjlr+gxq1Sq14DZ/uEt93Oo7/d/mX8zEXWfos37w/YH3zt0fIdvsd1/UETZi02v/A32zVv26Grzg2fumCluXiur/d1rF6TFq01hv57zKyl66u9V7+R/nTu1X/ojoBzN5f/evBE5uw5czuaa836jT5Sv0Wb9h3Wdbf5n7m+69jFO9pNY2/vjHsVo3i1xlu1y/+knr/G0sK6dSwVNd/qd/ra9sNnbziqlaHg2Gbf4Mtr9x05q0X3UTOXrNWY9gCBOaaz96AAgvfpm39MXLhmW6OPP/1i9e7Dp2SkGhYaX++sfjf0HMx3s0ylajV1rs+QcdP0Xiv4ICtH81EAROPrd6zVl1276x2Wg5kyzZyvAgzqr7oezrw/CqLsDbryYObKrftUdLxG3QZNR89auk5jzF37q49qmJjjaH46PnDcjIWayw+DxkwxzymAqHOFS5at4Mx1aYMAAggggAACCCCAAAIIIIAAAggggAACCESrgBY9y1SqXiuki0xetG7Huv1Hn9ldobbKzb/nxOX7WvBUcML8WtscR2mFtMCs8+afaUs37jJrL1iv1+WHAcO0mKoFXkfzUOBBC9aLt3gdcXReuzO0K0DX0Th9R06arUXwyMJpIXhf8NWH9gBLZMe19t944MRFzdd6rHzVmrV1XAvcCgjp/uzX1P2NnL5o9Z7jl+6ZuyHMAIICLXKevXq7t9XfHM/+rKxjy9p8Hrr3sbOXbTALfNvn4Iy7dqlongpUTF2yYadZXN0+VtnKNd5VMKVj958HOfJVwEVBHPMZd+8/fLy5w8PePjz30LJ95+/0zjwNQgwdP12BIc1F/1bgq++oyXNU68O8hsbWDhWr64wVW/ZWqP5uXUfzVuots60Ce47SdCnooHuz7owI6x1r2qpdR+scVu85fPqjNl98bd9Ro9+pLYdOXVVbBcasabUyZM6a/Wkww0jRFdb1OI8AAggggAACCCCAAAIIIIAAAggggAACCPzrAvqa21HOfU1MdSXMGhiOJqoaElr81cK/i6u7Z0g3o5oKSr0U2s0a9ZGzhBTQMPtp4d76dXlk8VQnwb1gkeKRHSe0/tptIOOIXsO6aK/dAQoyWBet9Xw8CxcvpQBSeHacyFEFm52ZV1S5K1gQ2hyNUheZtLgfUm0O+1ydvQe9V2aNFKWZUpDG69SNJ9qpEtL9u7h6FNBctOgflpGCe28aab5CaqedMRorrHHs5+WgHSmq12LfgWNtq2urdoij8RX4Ce0+wzsn2iOAAAIIIIAAAggggAACCCCAAAIIIIAAAggg8H/awaCUQFBETCCfR4HCK3f5BZspsSI2Cr0QQAABBBAInwBFt8PnRWsEEEAAAQQQQAABBBBAAAEEEIjhAvrCPldeV48AP1/vGD7VGDk91XqYtGjt9gN7d+1QUevDh3ycKoAdI2+GSSGAAAIIIIAAAggggAACCCCAAAIIIIAAAggg8G8JKPXT08LNRlHqf2sOsfG6ShulwvKqV9GkZduvlE5LabVUhDs23g9zRgABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEDgXxWoUeeDJgpYuBUoXOxfnUgsurgKky/evD9ABd0LFS9dTlNXbQo5ehQqWiIW3QpTRQABBBCIxQJxY/HcmToCCCCAAAIIIIAAAggggAACCCDwnEDOPK7ufzx58sTIZeQLT9gCWbLnchk/b8Wme/fu3W1aq3zRs6eCT6iXiqzL8Yif74GwR6EFAggggAACkRcgYBF5Q0ZAAAEEEEAAAQQQQAABBBBAAIEYJJDDJZ/byaDAo/eNBfgYNK0YOZVEiRMnGTp57rL/e+WVV9o0qFnx3JlTweZEPQsXL3UswO8gjjHy0TEpBBBA4D8pQNHt/+Rj5aYQQAABBBBAAAEEEEAAAQQQeHkFcuTO43rU/5DPyyvg/J1/1OaLrzNkzpq9d+f2razBChUuL1KqXEVfrz07nR+NlggggAACCEROgIBF5PzojQACCCCAAAIIIIAAAggggAACMUjg9TfefCtFytRpSAfl3EOpUbdh05PHjx3Zun7VMmuPgkVLlpHlrq0b1zo3Eq0QQAABBBCIvAABi8gbMgICCCCAAAIIIIAAAggggAACCMQQgey587pqKkplFEOmFGOnETduvHjpMmTKEnjE/5B9krUbfvTJvbt37+zevmVDjL0BJoYAAggg8J8TIGDxn3uk3BACCCCAAAIIIIAAAggggAACL69Ajr8DFoEB/gQswngNnjx5/Pjhg/v3tZPC2tTF1d2z8ju131+5aM6MB0YBi5f3beLOEUAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBCIoMB3fYeO3ewbfDmC3V+6bgPHTl+wN+jKA88iJUonTJQocfEyFaqs23/03O7Ai3fTZ8qS7aUD4YYRQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEIgKgRkrtuwdN3fFpqgY62UYI1WadOlX7DwUdODMrT/NP16nbjypVb9xs5fh/rlHBBBAAIGYJRA3Zk2H2SCAAAIIIIAAAggggAACCCCAAAIRE3g1Tpw4OXLncV00a+r4iI3w8vW6eOHc2QZVSuRXzQoXVw/Pm9evXV02f8aUgEO+3i+fBneMAAIIIIAAAggggAACCCCAAAIIIIAAAggggEAUCLyVPMXb2i2QM4+rexQMxxAIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACL5vA/wOFkJLcZvyoMwAAAABJRU5ErkJggg=="},{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO3dd5wcZ3348c/MbO97e72frqr3YklWsS0bN7ngEmxTgjGOAzghvwAhBEggIaTQk5CACeCYEMA2ljsuclOzeq/X+97t7d32PvP7Y6WzZZ1Oe5bkk33P+/Wal3S7M7PP7t1895mnfB9Jp9Pt0zStHkEQhLOQJKlZUhQlmslkzJNdGEEQLl2KosTkyS6EIAjvDyJYCIKQExEsBEHIiQgWgiDkRAQLQRByIoKFIAg5EcFCEISciGAhCEJORLAQBCEnIlgIgpATESwEQciJCBaCIOREBAtBEHIigoUgCDkRwUIQhJyIYCEIQk5EsBAEISciWAiCkBMRLARByIkIFoIg5EQ32QUQJsZitaHX69HQSMRiJBKJyS6SMEWIYHEJM5isLLn8CpauWEXTrDk4nQ5SyQSRcBhZp8NmsyPLEp3NR9m88Q/84ekniMZE8BAuDrEUwCXI5i7go/d/nrVXrmHnppfZ+torHDqwlxH/MKqmnbavTm+kbvpsrrzhw6xZcznf+sL97Nl3aJJKLnxQKYoSQ1GUKKCJ7dLYZi29QvvNi1u1P7r7bs1o0E3o2Ir6OdrvXt6mFXock/4+xPbB2hRFiSqyLH9F0zQ9wqSrnrGIv/+nb/HFe+9g86YtZDLqhI4P+r0Y8yqYVmxjOKHnRw//DmMmyKFDRy5SiYWpQpbltGizuIR85st/z/f+5nN0dPVO6DhJVnA4nUhAOpXEk5fP/V+4i6d+9RB3fuw+/vDCK2cck0zEiUajF6jkwlQggsWlQu+kscLO1h37J3xoYUU9f/X1v0OSsj/LOgNz587Brk9TVDODv/3uj8845sSeTfz7D390vqUWphLRZnFpbJLBpT312hZNugDn8lTP0n7y859roNc2vLpl0t+b2N7/m6IoUTEo6xKhJUc40Ozj5puuO+9zFRaW4vX2Ys4rIeL3XoDSCQKIBs5LyK5tb/CnX/0XZs+oo6+7k+Hh4Xd1nqqZ86jKM+MNa5QXWNj40sYLXFJhqhENnJeYkYFuHrj9Q1y5/g4+97XvUFyUT2fbCbraWhnw9jE06GNo0MuIf5DBgQFCweCY5zHoFdIplbkLl7B3+zYAdEYrD3756zzyo39gYCjwXr4t4QNCBItLTCad5IXHH+GFxx/BYDRTWVtPZfU0ikpKqZsxmyV5a/EUFuHO82C1WuluO86zj/2Kl154cfQc6bSKosgsX7WKb3/mBwBcd9f9LFm+kq4Dl/O7x54e45Ul6mfOwdfbzvDwW8HEarMTCYfGLqwkY7GYiUYiYz5tsrq44ZZbeOZ3jxBLpMZ930aTBZvdytDg4PgfkDB5RAPn+3eTFZ1WP3uh9t2Hn9I+/elPjj7euPgq7aHfPqX99OH/GX3s9k9/QfvDzhPas1v2aU++sVubPb3utHPd/5Xvaj9++Lfab//wmuawGDRAs+WXa4+++Lqmk9AcJbXaN779rdOOWXfn/dqXvvwlDdBu+PiD2rorlp/2/N/86Nfar55+Xbvh+qs0JFn77N9+X3tmyz5twdwZp+334U/9hfbYy9u0n/z2Oe3fH3rogjTyiu3CbqKB831OzaQ5cWAXf/dXn+eq9beOPt7b0cKMBct4/H8eGn3sdz/5F3btP8LffuYjPPbk89TWTxt9zmgv5NorF/PZj99B93CC4nwnAFffchevPfm/pDUoKqnAZra+7dUlbvvIPTz+v78EoGZaAxLK6LPl0xfTUKjj6adfxGg2ce1HHqDcnuYHP/x3li1bMbrf8uvu4qoVc7nnust54O6b+fY3v4l28rm111x/AT8t4XyJYPEB4CkoJugfGv05NNDBieZW9u3dO/pY46K1VDgy7N5/hNLScvp6ekafu/Xjf0J4oI9Zyz9Evi5KS/cgisHCnR/9OLu2bQYgv6iEUHRk9JiGRWuo9ig0d/Rnny8+/flb7voET/32f7Dnu5BkG5/4+J18+2+/itlkIxQLAyfbUb74ZR76/j8QS6S48WOf40PrVgHQtPhK7r7nzovwaQnvlggWlyJZx813fQJPnuucu5bWNPE33/wHfv7jtw+wUnny8ce555P3AWC0uvjS17/J97/5FdIZDavVSjwSA6Bm1hJuum4t9uq5fO5z9/Hlz95HRoWP/9nXKPE40DIqIHHVdeupqKjNns/i4Itf/TvSyWw7hM1TwtKli6k8+fyMxVeweGYFGzY8jcdTxA13fZLf/+x7jIRi6PRGNC0DwCf/399RUZxHNBxCZ7Sw/tbbUdMZZJ2Rv/jK1/jxv/7jBfpAhQtBzDq9FEkyt33yQT58x50M9bWzb9cOOtpa8Q0OoGkaZquD8qoa5i+7nNIiNz/+9tfZ9uaO006hM1r5zi8eJdB9jIrG+bz2+5/xi58/DMC1d32G9euWsXnbbtbfdjvf+LNPUDl/HbfeeAXPbNjAzMWrKbKp/G7DS9x33yfo6h9GDXThqJrPYOs+ps1azLMP/4DG1bdjTvmpaJzDHx7/Nbfd88dsevUVFi5ZzFceuIe2zl6+/fOnmFnl4Lar15JIqzQsXM03vvFVmtv7sRDkuY3bufdTHyeZUdC0NC//73+R8jRSXwDf+Po3JuHDF8aiKEpMBItLmCTJVNVPZ9bc+VTW1GKz2ZAkSCXidLe3cGD3do4eOYL2jmnrpyh6IwuWriDk6+Ho0WNvPzMrr15PWbGHV59/Eu+AD4AZC1cwb95c+jubee3lF8moGnUz5uG0Gdm9402MZgcLl11GT+tR2ts7UPRGFl62Em/HcTo6uiirbqCmppK92zcTPllzqahtQkqF6ezsHn31htkLcVj07N7+JqqmUVhagZqMcdVt99FYU8aMOU186sPXE4qK3ByXCjFFXWyX1HbXA3+jbTrYqs2eUT/pZRHb6ZvoDREuGbLOyLLVq3nk377NgcMnJrs4whhEsBAuCbfd9/+Y1VjD8NDQuXcWJoUIFsKks3nKuOPD1/PrRx5BlsSf5KVK/GaESXfzRz/Nc7/+L4KROBLSZBdHOAsRLITJJem4/obr2fDoo+gUAyl1/DkkwuQRwUKYVBVNCwl1HcAXiGJyOIi+bRSocGkRwUKYVNPnLmD/7u0AFBUVM9gnkvVcqkSwECZVQXEBAz1dgER9Qy0tza2TXSThLESwECbViH+EorIK5q26gaT3CEOh+GQXSTgLMdxbmFRWVyHf+reHsChpvvWlz9HW2XPug4T3nJgbIghCThRFiYnbEEEQciKChSAIORHBQhCEnIhgIQhCTkSwEAQhJyJYCIKQExEsBEHIiaxpmggYgiCMS9M0RdY0TSQQEARhXJqmibREgiDkRgQLQRByIoKFIAg5EcFCEISciGAhTEmSJNr1J0oEi7OoqW9k+ZqrqG+aOdlFueAUnY4FS1dcsPPNWbD4gp3rYlJ0Om7/6L1c8aEbWXnFNbg9+WfsY3c4aZo1dxJKd+nTTXYBLlXVtQ288vxTlFZUXdTXkWUFVc1c1Nd4p8WXXU5GVS/IuSRJIr+o+IKca6IURSGTyf2zy8svYM+OrTQfPXzWfarrGujr7roQxfvAmRI1C1mWcbnzJnRMJp3GYDTS29VxkUqVVTWtFgCD0XhRX+cUSZJomj2P/p7sBWGxWs/rfG5PPiN+/+jPK9auw2yxsnDZhau5vJ3BaESSJCRJwp1fMKFj6xqm09U+fo7PgsJi/L6BnM7nnODf1PvdlAgWeoMBu9M1oWP27tzG3IVLR38uKa8EwGS2YDAaMZktyLKMwWjC4XIDYDAYKS4tz/k1JEnC6c5DkiQKi0snVL53a/aCxRw7uB+/bxC7w8mNt92FK8+DxWpDp9NRWlGFxWrDefI9udwnn9PraZg+C8h+QxeXlqPT6amuraet+RhWmx2Ara+9jNVmY/ebW7Da7FhsNhwuNyaT+YK8R7vDBZKE0WTG4ZjY77SgqIQ5C5awcNkKJElGp9NTXlXDnAVLkBWFhctW4vbko6oqM+bMx5NfOO753Hln3sZ8kE2J2xC93oCnoBCDwYjRZCIYGCERj5NKJkln0gAnf05gdziRZJngyDCeguwfy6qrrkVVM1isNhqmzyKTSSPLMs3HjjBjznzKq6r5z+/8I1detx5N03h+w6M5lctssZBOpzFbLEyfPY/rbrkTu8NJNBImGg1jszkIBQN4+3oIB4MERoaJRsOEg0Fi0QiSJJOXn5+9cJwuYtEooBEJhwgFA9nzRCKjr2cwGrFa7QRG/MiyjKwopNPZ97L08rUYjUZq6hvZs30rTpebg3t3UdswHYvVSjQSZsg3iKIo3PmJT7Nv55tMq2/CYDSyZMVqTCYzG377CMtWXcG8Rct4/Ne/ZPa8hciKws6tm1i++kpUVeWFpx7HaDRRWVNLJBJGzWRQdDpUVUWn02G2WDGZzVitNiw2O/FYFEVRSCaTxGNRikrK2Pr6Rmx2Bx/7kwcZ8Q+RSMRRZAWD0UQ4FCCZSNDX0423r4eO1hMMD/kA6OvpYseW10c/j5r6GSxduYbfPvwQV127np3bNtE4cw51TTPQNI2GmbPZ9vpG7A4nsqKgNxgwGIyoqorN7iC/oJD2luMX6K/00jclgoWmaaOBIi+/gKLSMlLJJH7fIIl4nEBgmHg0CsCi5at45fmnAIiEw1htNtRMhp6udmRZprSikg2/eYRZ8xZSXFqOt6+HSDhEeVUNNruDA3t2AmC12XHlebA7nBQUFaPT6XHleTCaTOj1BjKZDCVlFbQ1HyMRj9N89BAvPfMEiqKgaRoAik6Pze7A4XRhsztwezxMq2/EZLEgSxIgEQoFCAz78Q/5CAeD2YslmSQRj512P19ZU8e1N99OZ1sLNfUNeAoK2b97B0cP7sPvG6SgsJj9u7djtlhpO3GM0opKps+ay0vPbmDdDbdw9OB+SiuytatwMMDBvbuorJ7GFdeu56c/+GcuW30lFdXTiEbC5BcVExgeoq5pJj/5wT8xrb4Ji8XKgb27AEgk4rQcP0JxWQU1dQ2YrTZsdjuJWJxUOkUkHCIWi5JMJtE0FVnRIcsybk8+5VU1WK02hga8vPnGK6OBWQOkU/+evE0xGk2j719vMJBKJk/7u2iaNZeXnnkCTVVRNQ27w8nBPTuYu3Ap/iEfb7z8PJqWDb4OlxuHw4XeYEBRFBwuNyVlFUiyjHaB2n8udVMmWJgsFrZvfu2c+xrf1nZgNpspKa+it7uDxplzef2l5052uWn4Br0sWLKcx371cxYtv5z8wiJefu5J/L5BACLhEJFwCICjB/eN+VqXrb6Sgb5ejGYzqWQCTdNIp9Ojz2cyGfyJeM730OPxFBTy9GO/pqezHbvDSf30mVRWT6Pz5D280+1moL+XopIyZs5bwKaXX2DZqrWUVVYz6O3DN+hl5twFFJaUcWDPTqbPnsfhfbtpPnqIZDJBMhGnadZcopEwLccOE4/F6Gg9QSadpqqmlpee3UAw8NZqY6qq0tvVMeE2Ib3eQH9vN4qi4HTnjQZWyAYKyP6+NSAWfatWVVPXQGdby2nnikUj9Pd243J78Pb2sP72u/nFj7+P21PA5ldfJJ3KLqWYyWQYHvKN1lAgG5DW3XDLlAkUAIokSV8FlMkuyMWkN+ipqqmjrfnYOfdNp9PMmr+Iypo6erra6WxrZcmK1TQfO0wyHqOzrQWL1Up/TzexaJTuzjYcThf9PZ3MXbSMVDJ52kUxnsaZc2g5dphMOj16a3QxLFy2Et9AP90dbaPv0enKIxaLMnv+IjpaTqDT6dGA5qOHMFus9HS1U15ZQ56ngO2bX2P1uusYHvKRX1hEUWk5g/19hIMBAiPD2XOmUjicLrx9vQSDIwSGh0drb6lUitnzFxGNREYD6LuVl19AT1cHqqoy6O3P+XxFJWU0zppDZXXtaA9XYNifvY1JJliwdAW93Z20HD+CxWqjvmnGuI2hsixjtlgZ6O89r/fzfiFJkookSQmyQfkDu+l0Os2V55n0crxzk2V50ssw0W35mqvGf0+KTgM0SZY16SK8P4vVNumfwVvvVZn0MrxXmyRJySnRG5JOpxnxD03oGKfTSWVlJXa7/SKVKlsVfy/IgO4CDViU5fH/ZBQlW0m9WNXzaCR8Uc77bqgTGOPxQTAlgsW74fF4WLNmDTfddBMmk+ncBwA6nY7i4mLmzJlDbW0tBoPhIpcyNzoZrigF/Xn+tmVZPmfQTSUTo/+fSvfzU8GUaLN4N/R6PUuXLqWsrIzh4WH6+vrG3d/pdLJy5UpuueUWFi1ahKqqBINBAoHAe1RiyPYHnCmjQaEZyqzQFRlzl5xomsZA//ifg/DBJEmSKmoWZ+H3+xkeHsZoNFJXV3fW6rckSTQ0NHDHHXewfv16SktLicViqKrKyEhuDZ3jkYB8EzQ6od4JLsPZQgLIytlj/i4fTHeB89Ko7ADZz85gNI9bbuHSMSW6Tt+NdDrNc889RyQSIZFIYDKZiJ4ci3GKLMs0NDSwfPlydDodkUiEeDxOW1sbO3fuJBgMnlcZau3whbmwphRUDSQJ7HrYMwQb2uDRNhh529ABNZM+67mSajZgNLngzfPvib0g3PlFzFq8hu72E7Qd2X1aN6hw6ZlSwUKSJPLy8tDpdAwPD5N8xyCddxoYGGD//v2YTCb0ev0Zz5vNZioqKlBVFZPJxGuvvcbBgwfxer3nPPd4DDLcXQd/ORd+3QzrnoGBWLZZutgMCwvgukp4cDb84AD88jikc7jOOsPQ4HzXxbqgZEVh8errWbj6Rnraj+HtaiESOv+amHDxTKlgIcsyZWVlrFu3jqNHj7J79+5x2yI0TaO5uRmTyUQsFjvj+XQ6TU9PD8FgkJGRETo6Ooif51iJYjN8Zmb21uOG56HtHcMIOiPZ7fftMM8D37sMbqmBB944d3uEqkFEtmEwZkgmznw/b8kOPJMk6eJ+20sKyUR22H3mPZ55K0zclGrg1DQNs9nMwoULqa+vZ968eXR0dIzbtqBpGqlUasyLJpPJ4Pf76e3tZXBw8LTRl+ei0+mw2+1kMpnRLtQSM1xZBvv98NMj4EuMf47+WLbm4THBvy6D/UPQPU7AyPMUcPn6T1A/fwXd7c3EY2Pv/F4khtE0jaGBHkaGBji44zWGB6fG4Kb3K0mS1CkVLACCwSCJRILy8nLMZjMWiwWv10s4PHb/vSRBUwXctFLh5jX5rJ2TYmG9itkAfX5IpbUJffsajUZqa2u59dZbeeCBBxgeHqa3t5dMJoPDAMdG4PBItgdjjNKc8UhGg20DcGg4W8uodcLhYQilTt+v1gF/f7mDuus/Tc2cpQx6+2g7fijncgMoOgNWhwuT2U4yGYPzrHXEo2H6OpsJjfjOvbMwqSRJUqfUbQhkB0K9+eabdHZ2snLlSlKpFOXl5QSDwdMaMO1muGYRLJsBs2fNpGzeA3gqlpGKB+lq3sZHdHG8ra/zzPOv89JulePdZ39NSZJwOp2UlJRwyy23cOuttzJv3jwkSSIajXL06FF6enrojZ7teJn6mfNxuj0cPbCT0Ij/jH1e74MPPQvfXAybboL/PgpbvBBIwhVl8NF6eLZ3iP5Dx5i3rAiZ3GtBALKio3HucuavuJpIJMjWPzyKt7t5QucYm2jUfL+YcsECslXg3t5eHn/8cUpLS0+7N5eAVXPg/lvzqZu+DM1xGSXTbyej6UkrOgqqZmItmEs6naJizh8zb80ubnnlazz90mF+9jyE39EUYLPZmD17NsuWLWPt2rWsWbMGq9WKJEn4fD4OHDhwzrEYJouFdTffTWF5HcWbN/LCoz8lMcYtxFAC/nQTzHDBPfXwtYXZrtYDfvjLbbCxJ0VR98/o7mxHzaQpr6zGP+TLaVSkTqentKaR2pmLiEWCtBzceYGCxeSTTi6fo2liENl4pmSwOCWdTtPZ2TkaLGQJblsN91xfSfll38bsmUNJSTmKoow2hGYyGVKpFA6Hg0BAY0SbTsM1/8t685cpL3ief/o/Dd/JHlNFUZg+fTpz585l2bJlpFIphoaGOHToEL///e95+eWXOXr0KJHI+C2TiXiME4f34sgrQdbpMRjNYwaLU5qjRv5mVxpJyyBLkHrbNdDT2c72za9id7pIppI5t0+kknG6W4/Q3XaMTDpFb8e5J+VJsozLUwQaDPsuncFcis6A1V6Axe7BmVeKxZGPpEkEhroIDHUTGO4llTxLNW8KkyRJSmiadgkN1Zk8H10HH7upAVvTX2MvXoSmaVRXV6MoCj09PSQSCaLRKK2traxbtw6z2Uw4HCaRSBAO+und8TWO7NrAV38Bw6Hs7ceMGTOoqqqirq6OaDRKLBZj3759tLW1EY1Gc27vMJjMlNU0EYuEGehpO+uYCrPVxrwlq9A0jX073iA2Rq1BkmVuvvOjFJWU8tKzG8bNSfl2eoOJ0pomYuEgAz1tnOsWwubI47ZP/xUms5XHfvZPDPZ25vQ6F4uiM1BQUsuCa+ox2TyEBmuQdSYUnQ6QSEZDjPS1Eh4ZoKd9N6GR/kkt76VEkqTUlGvgPJvVc+Cv/+wm1LIHqZ11BR6PB71ej16vp6WlBaPRSFlZGZlMBpvNRjqdxuVyYTAYMJlMGE0W3BVrUaKHKLG0sulAtqvS7/czNDTEnj172LVrF/v378fr9ZJKpc5dqLfJpNOMDHkJB/zjVpftDifX3flpZixcSTQ4TE/HGLcKmkZ5ZTXbXn+F2+65l51b3sgp8a2aSRMY6icSGs6pzLKisGj1jeSXTiMc8NPZfDCn4wwmM9PnL8flKSQ0MjShpLxnY7a6mb5oPQ2LL2fmVSO4K7wEBxXSCSfpdBJF0aFKPvIqhzBZHJj05QSGe0inLk7agPebKdkbMha3Db712VpcM79ApzfN7NmzMRqNmM1mVFVleHgYt9uNzWYjk8ng8XgwmUwYTmZNikQidHR0UF5Rhat8DTr/Y3gHQ7T0ZttHYrEYiUSCTCZz0UcpapqGp6gUd34xXa1H6W47Pe2brCh4ikrxefuRZInmY4dZc/X1HN6/+4KXJZ1OEYtGMZjMtB7Zja8vt5pF5bQmbv3jz1M3axHR4CB9PedXI7HYPMy+7DbcJTWomp7e4zp6j8volAZQdUhIGKz95Nf0oqkmGlf1EAurkChn2NeFJsaAiGBxyt1XwnW33Ie94kMsXryERCKBwWBAkiSGh4cpLi4mkUjg9/sJhULYbDYURaG7uxu73Y7BYMBms6HX65EUE4ODw9RYtvD8Dki9x39nmXSa9hOHOH5gBy1H95NJn16DKSyrYf3dn6Fx9gKaD++mveU4V123nv27t49mhrqQfH0dtB7exUBPa86zUI1GAw0z5mFzOGg/tp/ezvEzco9HkmRmLr2R0ul1FDU2o6r9ZBIVSBSCqhutOaTiEBpKomkt5JVrOIpjRPwailbOiK+Tqd5rI4IFYDXBX30sj7JFX6G8eiadnZ1s2bKFpqYmIDv7VFVVwuEwBoOBdDqNxWLBbDaTSCQwnkxNr2kayWQSi8VCSs4n2PY7fMNxms9jrJHTADNdUG6DGW4wKhBPZ+d5jCeTThMOjpAZY5CYTm+gad4y7M58Bnra8fZ04h8aZO2HbuTgyRyZp0hk82BYdOA2vjXFPZeh5W/RSCXjE5quHg2H6Wk/xomDOzl2cM95BTG7q5jLbqmkamE79oIAjgIbFgeEBt3IsoKiN2Awa8QSz1JQM4jZmSA8ZCM6opDRhshEC4iFo8Rj5zfP5/1uSo6zeKfbV0PdzLUYHTWoqoqqqixevJh0Oo2iKKNtFvX19QSDQfLy8vD5fKPjJjRNG508VlpaSjKZJL+omv76T3L3ld/ljQMQmeBtr06CO2vhk42gyNAXzT5WYctesD89Co+cgPC7uIYCQ16e/b//oqy6gfbmowCcOHKIa278MHqDgUwqSbkVri6HpYVQboVSC+SZsm0wGQ32DcGmftg9CB3h7DDz1BixwGi2YrO78Pv6JhQsNE2lu+PM2oRRhsUF2a7gQI7vvai0EVd5EE2KMdxrZ/D4XEyOJIou26avqSrhQA/ppIe+w9OJRk5QMb0STY3iyncSK+rH1V/ByJBYeGjKBYt3zne4Yh44imaj0xmIx+PE43GsJxfeOdWtWFtbi9/vx+VyIUkSJpNpNCOUJEmYzWYaGxuBbHdpf38/SdNcVi904bSOnBYsJElCr9ePJsbRNO20XhGPEb40D8wK/Mkb0BI6OeMUUCSoc8JnZsBj6+D2FyF4lotGkiRqGmahaRodzUdOW/XM292Gt7vttP1btjzLv/7JLTSe+A21Tjg+Ai90w8PHoSucDVoAhSaoskO1HT7RCI0uSGayk9le7MlOVjtl0errmT5/BZv/8FuO7N48ZjllOfs5jrcqm0y2ZvWNRWDRw50vnXXX0+j0JuxuN+GRQVwlBXS0LCKVMJAa1KFpp+a+ZNDpzRTVuUlGQyRCc9DYjat8mKHuGOlMGruzHklWpnzbxZQIFhaLhYqKCoqKinC73QwODtLS0sLAwAAOq4bZWc9wKIROp8PhcFBQUIAsy8RiMVKpFBaLhYGBASwWC1ardfTCzmQyyLJMJBLJJsF1Zqd0GgwGkhkDFlc1ZuNeIJscp7S0lJqaGqZPn05jYyMOh4Oenh4ef/xx9u/fD/EQt9bANi882XF6dV8j+/PREfjzrfAPi+FXV8BHXobwGL2oBcXl3HT3/WQyKR7/5X/Q3X7ijH1ksjNY766D26p30jb/w/z7s79hYzf44jBWXaAlCFvfNsXdIMOcPPhUE3xuFrzUA9/bDz1RSEQj6A1mqhvmcHTv1jNqFwajiZXX3I4KbHvp98Sjp3fzykClDf52EVxeAk+1wzd2Z0el5sJkdmB2QSI4m75jCZLxOGZXkERERU0XgSoj6bxUTD9KSUOSTErF23qEfc+VUliTJB2ZSSKYQVYiSEhTvNViigQLq9XKggULWLZsGel0mmAwiNvtZvPmzSjyCJlUBF/Ih8lkokAHMnkAABRkSURBVLy8PJs5enCQeDxOUVERgUCAWCw2mqpf97ZFcU41fJ6aGAbZwJDnyUdKZAd66fV6Vq1axcqVK2loaKCgoAC3201RUdFooAn4vBSEQmzxwpHhsS/UUzIafGVHNmD8bDV86vUz54IUlddgc+ZjNBnRvyO9n16CBQXZC3xtKTzeBmuehMVKC9toYDBxArPVSjKRIJ0ev76fVGGnD3Zuyk6E+8u58ML18JMj8LMdLxGPRwn4B8a8DTGaLFQ2zMbmcNPTdowTB7ZnH5dhVQl8enp2Zu2GdrjxuWygnMgYy3Q6QSwo4yrtIp0oQmcwEguATm8nkwFJBlQnGmFCQyr2fBNFtQaqFvg48FIZEibyyyrwNu9Fm/KhYorMOpUkieLiYnQ6HTqdjpaWFnw+H11dXdy8PIWreAZ5VVcRiUTIy8tDVVUMBgMejyc7O3JoiKKiIux2O8FgEL1ejyzLqKpKNBolHo/jdrsxGo0cOXKE4uJiwkE/tpFf8pMnQwyHoKCggNraWmKxGHq9PhsgAgEOHTrEa6++yvGDe+gcSdIVya3dXQM29mbbFb40D0LJ7Lf+qQloiXgMu8vNQE87u7e+QjqVRC/BvHz4zmXwsQbY2AMPboENHeBPQFdnO9ffeicD3n7+6N4/p2JaPW3HD+fcwBhOZ29dNvZmA9Fd0zK0trezp2MQdYw3lUomyKTiqKpK66GduNUgt9XAt5dm22xe74PPbs5Oxx+IT7w/Ip1Kkpdfi5ZZRiJip3b5Fvrbj5EMl6PTm9E0FUkyMtThIpUwkE57cRUZcZdqtO/N4C6YTyoRJdDfxmDv1Fl5bCxTpoEzEomwceNGtmzZgizLJJNJYrHsil3DIQgPHsBa/9ZH0dHRwaFDh7j22muJx+OjtYhT59I0DY/Hg9frxeVy4Xa7sVgsaJqGzWZDkiRSoRYCw/3Ek29NXuvq6hrtXdE0DVVVSSQSDA0NkU6lJnwxqBp8cRtcXwWfm5nNqrXTl62ZDMQHib7xX6iSjltKwsxww5qSbI/Kc13ZOST+d0yBDwz7sdkdWO1OCsqqKamcxu6tr9J6bGKzU4+OwG0vwo1V8MV52cDx38eywSmYyl70sgQGWWXkyBs0jGzjWw1JriyDXYPwL/uyM2lzvd04O43BvuMUVM4gmfKjN6aonqcy0ref4a4q9PoqkCQMpgIiPidmZz/+3giZtITNcRloGtHhAYLDfUz1rlOYIrchwGjj5Ts9tRXKi18jVXaChulz0TSN8vJyZFlmeHgYnU5HdXX1aM6JVCo1OqIwGAxSVFSEyWQabceoqqoiEAjQvOM/GerM4D+ZvCaVStHRceFXZFeBpzrg2U6ossHyIlhSCOurNBJqjLQKw4nshfeNXdn2hnfesrxd89HDoKZ5/rFf4vYU4u0dZzrtODIaPNEOz3TC9ZXwJ9Phn5dBXwQSGTDpsgl+QGMglmRjTzbZz/GRiXbNji/g7yEaGMRpraZzfwfzr/NgMGlsf6KFQFdFttdLp0dWwFlkRGeIERzMkE6G0NI64kE/QwPvfpzHB8mUCRZn8+x2uG1VhOihh2mc8V2i0Sg6nQ6LxYLf76e6uhrINmYGAgEqKytHA0ddXR39/f1kMhkqKipGezZ2bH0RXWgrv30V4uf97XgmWZazK7+8rR0go0FrKLs9cnKE96kpYhO59vbv3s6yVVfw6P/8jLdWD82BJCHLyhlzVlJqNmg82QH5xmzS4RJLNk3gUCLbLRxIni1/x/lLJsL4ek9gduaTSdSRTrbj703g75iJTpFRMynSyTiyotB3eDqls7ZhNOXjLOmi72AEb88RYpHchrd/0E35YJFIwYYt8BH77wmOfJlURh5tf/B4PCiKMnq74fF4CAQCuN3u08ZhGI3ZlbX7+/s5fPgwQ0d/TjygsjW3+VkTkl9cwewFS+nvbqP1+KFxlzx8N9efb8CLOy8fSZJzmrJtMluYVt9Eb1fH6FKGY1G1bLvDwCRMtejp2IPDXYI5L01kJMXmXzlxuCtAkjCabWTSaTRNJeJ3k4q5aNvhIupP0XlsK96ei/BLfJ8SSwEAz7wJQz4/0b6X8fv9qKqK1+tFkqTRRtFTbRUjIyPEYjHC4TDxeBy73U5eXh4DAwMMDw8T7N+NI/kaD78IyYnllzknvcHEzMVrWHHd3axd/1GcLs8EzyBRVT+bhatuwOHOH3OPVDKB1WrL+YzTZ8/n3ge/xMce+DzGHBdjeq8l42FaDr9K3yGVF36gR9ZqSCfjJONhIiODqJkUmqoy0tvGrkcN9B7xsn/Li/R3HxIZx99mytcsIDvC8j+ehJlL/kDRgrdGb55K0mu1WvH5fOTl5VFVVTWaudtsNgMQjUaJRCJERjoxDfyQTfvTbLkIX0jpVJLBvi6Gh3xkVI1YfLyku2dSFIVFq66hbuYi8gsLeOmJ/zljSHgmkyGdSeecCGZkeIhkKk1hSQVOdx7x2KWZByIcHODw7udx5ZVjdwUxW13Iih40DUlWSCVjhANehn0dRCPDU34A1lhEsDhpdzP8/Q+f57v/uoaEvBKTyYmqqkQiEfR6PU6nk0AggN1up6urC4vFMjoIKxqNMtBzCP+uL3Lo2CD/8eR5p6cck6apHN39BoEhL5qWIRSY2L10JpOmp+0o5dX16HUKiqIbc/5IagLLGHS1NfPk//0Ch9NFOPRerr42celUHJ+3GZ/3VKNOtlVHQhJZsnIwpZPfSJKEy+UiFouN9pRcu9zJ33/1s7grVuMNmCgoKsXlcmEymfD5fNjt9tG2CgDfoJftL/2ITPcvOXDcz/cff2suiNPppKioCLPZTCaTQZIkwuEwfr+fWCx2XmuLvFuKoiO/uJRYJExwjFyeAH/8p5/nkYf+PeegoSg6ZEWeUJA5HzITG5wlnD9JklJTNlicGqhVWlpKJBLhxIkTo12ic2oV/vLexcyfP5eEvglX2QoceVVYbTb8fj9Wq5Vw0E93y3aiJ76Dr2sXT26F370Oqbd9UVdWVrJ27Vrq6+tpbGxk2rRpo9m1+vr6+PWvf82mTZvo6ek5497YpGTnXyzIz+bUTJzsAu0IZQdfdYbHHuZ9IVx78x28uelVRnwDOA0wKw9m50GBGdyG7ELLI0kIJmHvUHYJAm/s4o9EcOrhqvJs9+oB0UHxnprSwcLtdlNVVTWaYbu5ufm0jEx6BZY0wYpZsLDJTEHlMvJK5+PMrwVJxu89xq7NT/Dsa+1sPgSDYyw9YrfbWbBgAevWrWPGjBk0NDRQXFyMy+UarVU8//zz3H///QwODqKToNgCd0yDdeXZiWPHAxBLZwczFZuza4RU2bP/f7IDHmuDLf0TG5sgyzKadvYlDJauXEODMcTyxC6uLDs5pHsQmgMQTYNByc4JKbdmJ7ZV2mCvD/7tUHbU5YX+1pfJLuH45flwIgB/sRXioknhPTVlg0VlZSWNjY3Y7XZaW1tpbm4+67ohACUemfm1GkVuDUWBUBQOtsPhjnO3Tej1evLy8vB4PNTW1rJgwQLWrl1LRUUFHo+HJ554gn/+53+m4/hhFhVkByqlVdjty35bJ1VQdDosVgfRSIhMOoUiZaeNX10O9zZlB1n9457cLlS9wcjcpauxWCzs2foqoeDpUa7cCp+/ejq3LmviqQ2/56dHs9/kibOcWAasevhEA9w/A7YPZMty4gKlf6iwZieSXVUG3zsA/3UYYiJQvOemZLBwOBxcfvnlFBcXk06n2bRpE62trWf9llUUhdraWtLpNO3t7aMDst4tRVGwWCyUlpZSVlaGwWBg9+7dDA4MoEhn1hAkSaKwvJbl19xB88EdHNq+8bTp3GYlu3zhX8+HV3vhS29CZJzbE4e7gI/++T9gtlh45ff/za6tr6Cg0eiEG6rg/unQnHbzf8ar+cWvfpPTrYXBaMaZX4wS8fGRihCfmQk/OggPHR2/LONx6OHDNdnh4keCOr6538i+viiq6MqcFJIkpabUOAtJkqiursZoNJKXl8fBgwfp7Owcty/dYDBQV1fHkiVLRns/TlEUZTRTVq4ymQyhUIhjx46xceNGXnjhBQYGBkanoL+TTm+kuKKOpgWrWXPzvbgLy057PpaB/22Gyzdk2xKeuDo7ZfxsErEIvZ2txCJRSs0qn27SeHgtPH9ddnTlva/BrU9HiBvzcgoUkiQzb8U1XHXrp8hvWML3D8pc/Ux2Svkb62FtyVjrqJ2dLMGHyuGlG+Dzc+DPtkh8K7CCsrV/TGX9rAmcSbjQplTXqSRJBAIBvF4vzc3NNDc3nzPLtl6vp7CwEGB0MtkpDoeD2tpaTCYTzc3NeL3eCQ/iOVdNJZ1K0tN2BG9PG3q9EUXRjTm6cjgJf/oG/FEd/N+V2faDXx5/65tdkSDPCNMcUeaceIh1cgF5RW3s1eDpTvirN6Enkr2NkeV0zt2geoOR0uoGisunMTzYw+Fdr9IayibmuasO/nMVPNYK3z2QzZFxNjLZGbFfmAtLCuCHB+HnxyCUkbhqaT1VTQvJqBpdLUfInGUZBOHimlLBQlVV+vr68Pl8JBKJnBYylmWZ4uJiQqEQDoeDwcHB0eeSySQ2m401a9Ywe/Zstm/fzp49e877VuXtNE3F19fBb374ZfRGE5Hg8FkDkkq2lrFzEP5lGdw3Pdv4ORCHegcUmaE3CvuGfPzlBh97h8ZuKFR0OkLnWCXtlFQqyd7NL5BJxWk7vBP1ZCOxBvyqGV7uya6Mtvkm+PlR+G1rdvHmlJoNYGVWmO6G22tgWVE2t8aXtmVXij/1ro4d2I7V6cHX13lBP1thYqZcm8VEuVwu7rnnHoqLi/nNb37DgQMHTnve7XZzxx13sHDhQjKZDD/5yU/Ys2fPJJX2LRLZVHQ3V2d7KwZi2YbTh09AW2j8Y+0OJzX1jezftX3sc78jNaGi06M3GEnEomMObjpVlr+en+0KzmjQHc727LiN2S7hR1uzga57rHwekoTZYieZiJ2RrVx4b0zJBs6JKigo4L777kNRFJ5++ukxA0FRURH33HMPK1asQJIkHnzwQbq63r8JXj0FhUQjEWLR8ZdVnCgZsBugyQVWHZh12eS/g7Gz97YIl4Yp18D5bphMJuLx+Li3LF6vlyeffJL6+nouu+wyrrvuutGEvu9HoUDgggcKyN4mBZLw5kA2m9YzndmahAgU7w9TIq3e+XA6nVRUVDAyMsLevXvPuohxKPRW3X737t0cP378giy7Nxner+UWLh5JklRxG3IOiqJQU1NDXl4e+/fvHzPb1ikGg4Hy8nISiQQ9PT3vYSkvjLz8QkrLKxgaHKCv5/17GyVceKLNIkeSJCFJ0ge+Jb5qWj3Dfh+hQHZUp8jlIJwi2ixydCq57gddV3sLVdPqsNrtrFp3LSazmZLySowmMxXV0zCZLciygsWaTUqsNxiwWK3kFxYBUFE9Db1efO98UE2pcRbC2VXW1NHZ1oyiKMiSTGdrC02z5pKIx8nz5GO2WLFYbRQUleD3DTDQ30dxWTnllTXEY1HaW07gzvPgG/CSSr33U++Fi0/ULAQAHKND2SUKikvo6WzHaDJz5MBePAVFHN6/G7PFit2RTQo0d9FSejrbUdUMg95+zBYLJovlovSiCJcG0RsiAGCx2SmrqGLEP0Q8FsPhcjM0OEAkHMJoMqOqKk6Xm7bmY9kkPsEAgZFhujvbyWTSmCxWqmvraTl+ZHQUp/DBIXpDhAtCURRmL1hCPBbl6MF9k10c4SIQDZzCBWEyW3Dneejr7pzsoggXkahZCIJwTqJmIQhCzkSwEC4JnoLCsyYRkmWF+ukzx3xu6eVrsdrsACxesQqb3XHa85U1daxedy16w9iV56ppdehOZmoXxieChTDpLFYr937uC5gt1tHH7E7X6P9deXmj+TUk+fQ/WVmWKSmrQJJlmmbOJZl8a2l4RdHhcufReuLY6DIF7zze6cojPU4CpHfuP5WJrlNh0qVSKfbtfJN0OoU7L//kwtRWUskkFTW12B0uNE0jnU6z8opr6GpvHR1RW1hcCpKEJ7+QSCRMd0cbFqsNp8tNWWUVRSVltBw/Qk19I5qaYdmqtXS0nKC0vJJEIk559TQy6TR2hxO9wYDJZMbpzsv+63Jz2aor6Olsp7SsEiRODkKLkU6lMJpMYy7S9EEkSZIqgoVwSUgmE1TW1FJaXonN7sRgMlJcVk5XWwuz5i9CpzcQDgVQVZWB/l4AnO48FEWH2WLBaDSRjMfx+waZs3ApDTNmMTzkY+/ObdQ3zcJssTI0OEA4FMRisTJn4RJ0Oh1FJWXo9QbMZgu9XZ1U1zXgcLkoLa8imUgQCWdnEzfMmEUiHqe0ohKjyURBcQmyrBAKXtqrsF0okiSpoo4lXDJKyyrpaGsmFo2QSiZRZIVoJEI0HCIcDGA2W/H2vTWbt7yymq72FuKxGIf27QIJmmbPRVUz9Pd0o2ka7jwPA/09xOMxisvK8Pb2UF49DYvVRl9PF90dbSQTCYb9PppmzSEWjaDXG0imkgz5BvAPDVJQXMLW1zdSXFrGob27AGiYPov+KTYzV9QshEtGNJJdmT4eiyFBtpqfSeP3DZJOpQgFR/AUFDE85AOyOVXDwQC+AS/pdHp0lmxfdycGg5GyiioikTCBYT8Opwu/z4fD6cRkNnNgzw7isShFJeUcPbiXqmn1dLQ2s2zVFbSdOIpeb8A/5KOgsJiBvl5CwRFUVcVstSFLEj1d7Yz4hybx03pviRGcwgdWw4zZtBw7PKFEPo0zZuNwudmx5fWLWLL3JzHOQvjA0jRtwhm/DCYT4dAFWkrtA0iSZTmuqqpxsgsiCBeUJJ17bUkhZ7IsJ2RJkj74WV2EqUcEigtK9IYIgpAzESwEQciJCBaCIOREBAtBEHIigoUgCDkRwUIQhJyIYCEIQk5EsBAEISciWAiCkBMRLARByIkIFoIg5EQEC0EQciKChSAIOdFJktSsKErdZBdEEIRLlyRJLf8fou286UTlJUcAAAAASUVORK5CYII="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydCcBNVdfH9Zb0Nr/NyZh5zEyGkAaFBqWJ0iDJUKJEhBAVCSljCCFFkkZliCLzPIekQaVRA1Lf+l13+67rnDs8nune53+yu/e5Z5999v6dc/bZe6291sqWTZsIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIZDCBYzL4/Dq9CIiACIiACIiACIiACIiACIiACIiACGQZAsfYdsqpp51OOumUU0898aSTTs5xwn//mz179uOPOy579v/YRp79+/ft2/39d7vWr1m57J8DBw5kGUBqqAiIgAiIQJYmIIVFlr78arwIiIAIZD4CeS8sWDhnrjz5jj3uuON2ffP1zs83rV+rCVrmu06qkQiIQPoRaPNot9579vz26+gX+j+VfmfVmVKbQK68+Qvs+vqrLxFApnbZKk8ERCDzEShfpXrNR3s8M+jdN1+fuPevP/8sVKxk6Tz5CxTKeUGevGede+75KCZirfWQZ3t3Gz7gqR6x5k+LfChR+o+cOI3PB+5sVD8tzqEyRUAEREAERAACUljoPhABERABEcgUBKrWrHNl+259+l9YqGjx0Ar9/OPuHyaNGT4YQd2+fXv3ZorKqhIiIAIikE4EKlWreemwSW99RP9Xo3ju0/ft/euvdDq1TpOKBMpWvLj6qKnvz1u26NN599xQ95JULFpFiYAIZEICx+c44YSBo1+dXqVG7csjVc/0GH/88fuePda1/0k///ff+/f/Y9u/ltxx7OvVqW2LTetWr8zIphYrVab8hHc+XvLrLz//VLNknjMysi46twiIgAiIQHITOC65m6fWiYAIiIAIJAKBeg1vbtJr4Ihx1PXbr3d+uXbF0kVM1goWKV4yf6EixVq069S9Rp0r67VsfN2VTJISoU2qowiIgAikBoHq1vdRzpYN61ZLWZEaRDOmjKq1L6vLmc85L+cFGVMDnVUERCA9CTz94uhJTlnxw3fffrNkwfw5G9asXP7F1i2bbKy74/td337zy08/7kZBkZ71OppzlatctQbHf7NzxxdHU46OFQEREAEREIFoBKSwiEZI+0VABERABNKUwHkX5MrT9ZnnR3CS53p1eWT8iMH9UVa4k2JO32vA8LElLipX8clBI8e3aXpjQHinTQREQASyAgGsz2jnkgXz5mSF9iZrGwsVLVGKtm00gWWytlHtEgER+H8CxKPgr39tu7FO5ZK23ubHROdTqmyFyrRhy8b1axK9Laq/CIiACIhA5ibwn8xdPdVOBERABEQg2Qnc+0CHLpjNvzZu5JCxwwb1C1VW0PalC+fPveuGK2rs/uG7XdUvveLqS+s2uD7Zmah9IiACIgABYvoUKFysBN9XL1/ymagkLgF811P7tSuXLU7cVqjmIiACsRKYMn7UMPJuXLtqRTIoK2hLiYvKV+Qzo11TxXoNlE8EREAERCBxCUhhkbjXTjUXAREQgYQncPzxOXJc0aDhTaw+GzW4fx+/Bn371c4dzz7RqR37m7Z48JGEb7gaIAIiIAIxEKh3wy23u2y4EYnhEGXJhAROPuXU03LmypOPqklhkQkvkKokAmlAoFS5ilUodtlnn36cBsWne5Gnnf6/M3LlzV+AE69fvWJpuldAJxQBERABEchSBKSwyFKXW40VAREQgcxFoEiJUmUQ5AT9+X4ZqXYfzHhjMgG4S5evdPEFufPmz1wtUW1EQAREIHUJHGNbvYa3NHGlfrVj29bUPYNKSy8CRUqULsO5UM6bwmJJep1X5xEBEcg4AoxXOfuyRZ/Oy7hapN6Zi5YqU871Y6awWJZ6JaskERABERABETiSgBQWuitEQAREQAQyjMCFhYoW5+S7LfJgtEoc+Pvvvxd8POuDfw4cOHDKaaefHi2/9ouACIhAIhOoWuuyum5V/u97fvv1j99/35PI7cnKdS9asnRZ2r9j2+ebuZZZmYXaLgJZgcCxxx13XPFSZcrT1hWLF36SDG127aEfs27sl2Rok9ogAiIgAiKQeQlIYZF5r41qJgIiIAJJT+BUsy+nkS4wYbQGP9Wlfesb6lQqsUFBS6Oh0n4REIEEJ9C4Wau2rgnffr0zogVagjc16atfrOTBlcnrVi2XdUXSX201UASyZStcrORFjG2/3rljeyyLchKBWdGSFwX6sTUrli5KhPqqjiIgAiIgAolN4LjErr5qLwIiIAIikMgE/jazCepvXqFispj41aIWkhK5zaq7CIiACEQjgPXZxZdceoXL983OL7+Idoz2Z14CRUsdFPStX7Vcft8z72VSzXwILP/ykFFQdstywNI/ZC2b+1Qx8yFQulylQPyK1csWLUwWSMVLlw1YjKxZvvizZGmT2iECIiACIpB5CUhhkXmvjWomAiIgAklP4Osvd2ynkTlz58l33HHZs//99/79Sd9oNTBDCJjA5QI7McKW70zI8keGVEInFYEYCTS9/8FHyLr3rz//ZJXuN1/tkMIiRnaZLZtdvhPzFyhclHqtU6DazHZ5VJ/YCfD+LGzpv5aWW0Jxoc2HgAu4nSzWCFhEu4Dbq5cvkcJCd74IiIAIiECaE5DCIs0R6wQiIAJZkUBwNdoJ1nZWoe2DgVaiHXknWNC+wGrT7NmPPz5/oSLFNq9fsyor3i9qc9oRCD6Lx9oZSlk63tLX9tsyex4DK0TDt5CVpLjNPJRHz2/aXSOVfDiB3PkuLFi/4S23E+tgyYJ5c2pefvU1TrkrVolHwNyolP3PscceS8DtDWsUqDbxrqBqHCRwjH2SSlraYek7kfEnULpcxYCFRbIoLMy6ogLt2bdv795N69as1LUXAREQAREQgbQmoBgWaU1Y5YuACGQ5AkGBJ/3reZYItHlKloMQY4O/+/brrwjeR/byVarVjPEwZROBeAmgqOA5PNMSq0SjbSdbBuKr5IiWUftFILUJ3PtAhy4IuCeOHvq8Lc4/ifLxg57a51F56UOgWDDw7vYtmzb8vmfPb6l11tP+d8aZZ597fs5o5R1jW7Q82p+1CNg4NYcl3ovxbCj+uZcY354Yz4FZLS/PJopn83r69/rVK5clQ/tLBV1coazYv39fYCFWVtmY11k6JvjJ90DSJgIiIAIikLYEpLBIW74qXQREIOsSYFJ3hqUClgICJ23eBObP+uAd9lSrdXldMRKBNCKQ38pFWcGK0LUxWFcgmMG64t80qo+KFQFPAnnyFyhUr+HNTbCuGD98cP9zc+bKTcavv/xiu5AlJoESpcsFViavXpF6blSwupm5dNPXMz5dtbVKjdqXe5E565zzzh/+6oxZi7b+sPeGxnc1T0x6qnVqEzBBK/P/0yzFOzZlXIsbqPWW9qR2vZKpPGdd8fmm9Wtx65cMbStb6eLqtCNZLEbivCbc++dbcq5F4zxc2UVABERABFJCQAqLlFDTMSIgAiIQnQDuoBA0sYItlhXd0UtM0hwfvTt9Kk2rVL1mnZMt+naSNlPNygACIdZORAb90dI6S9HiVzi3F1hXaJyUAdctK5+y1SOP93LWFb/8/NOPCJ3h8c1XO3HBoi0BCZS4qFxFqp2aft/bPtbjaVwpHn98jhwP2ncvLP1HvDK1YtVLahMfqmLVGrUTEJ2qnDYEeK+hrDg5qLyI9Sy8R4kzdrYlWe1EoJZs8Sv+Y5tTwqxduXRxrDdMEuXDjXpxSxdZwnpemwiIgAiIQDoQ0EQ8HSDrFCIgAlmSACu0t1jCz2uWMp2O92qvWLxgPq6hELxcdvW1N8R7vPKLQBQCKB4Q+uayVMgSz2akDVcXCGZ4bvXs6vZKNwK4Drq8/vWNcBuEdQXBtk86+eRT8Bn+4w/f7UpJRVACn3v+Bdz72jKAANcvz4UFCVScbU0qBqrNmTtPPtecXd989WV407h3nNCUfUsWzJ+TAc3XKTMnAYSvLA7BTWI8igfejbhKJOh2PMdlTgppWKtSZStWpvi1K5clhXC/YNESpU6ylwltWrdy+ZI0RJdZi8bi1lndylVoZr1KqpcIiEDSEZDCIukuqRokAiKQSQhgAs6KbjbP4L6ZpJ4ZXo1/bHvnjcmvUJEGNzW+M8MrpAokGwEm2SgqWBXHylBcWkTaXOwK8gWeXQXcTrZbInO2h1XzxBt4ZeTg57CuOOOss86hpqar+IaAzfHWmhX4r7w9d/GIyW/PjvdY5U8dAkVLlinH6mTzCvPH5g1rV6dOqab8CApCt2xct6ZnhweOcPe0b+9ff21ev2YV5/ts3uwP35g09qXUOrfKSXgCKO15v6F0iKdf+cXyf2vpZ/duTHgSadAA+nBnVZUs7pMuKl+5Kqj+/OOP37d/vmlDGmDL7EXyrGA5j0soKSwy+9VS/URABJKGgBQWSXMp1RAREIFMRoCVaHUsXWqJAL7aIhCYPvmVMewuV6lqjYJFipcULBFIJQJMMnn+sHRaY+krS54Ki6D7KJcfdxlMTrWJQLoQqFrrsrqVqteqs9u0Ey8PHdiXk57+vzPP4nP39ymzrqh1Zb1riYnxw/e7EDJqywACTnC5bvXypQTgTa0q9HikdbOnuz7yQNNr61zMPRNeLgqu26+pU+W2qy+p0PL2hnVT89yp1QaVk2EEsBzENSIuS2O1lEDJUcJSPUt5LeEaSpsHgbwFChUxw7bTEe6jUEwGSGUqVqlGOzauXbWCRUbJ0KYUtOE3O4ZFBOem4FgdIgIiIAIikAICUlikAJoOEQEREIEYCKCwYBUOlha/x5A/S2fZtmXj+uXmGgoINze9t1WWhqHGpwqBEAVEESvwEksoKjaatUSkFaUIZXAfxTGalKbKlVAh0QiwAh/rCvINfbZ3tz9+/z0Q0PaU004/nc8ff/ieYPFxbwRm5qBVSxctiPtgHZAqBA6ttE5Fd1BU7IutWzZNGj3seXeveFWWYL/rV69Y+s+BA9GsylKlrSokYQicYTXNE2dtkRlUsYR7Oe4nyRB8AJYuWxFO2datWrYkWZ69iyoctLDYuG7Vijjvm2TJjmIPhTNjRFyqaRMBERABEUgHAhpspANknUIERCBLEkBhwQo0VrCpr43hFnh93EtDyXZ1w1ua4Pc7hkOURQSiEeD5Q/mQzxKrSn+IcgB+vXNbQmkRLTh3tHNrvwjERKDBjbc1LVSsZOltmzeunzrx5ZHuoFNsmS7f9/z6Cy5Y4t6ckEkKi7jRpdoBJcqUDwTcXrVs8cJUK1QFicDREWB8xYKanabAj0eZxeKbOZbWWko1a6Gja0rmO7pU2QqB+BUrl3z2aearXfw1Ouuc886/IHfe/By5ZcO6VHNrF39NMvQILG6x0F1nSWPDDL0UOrkIiEBWIiANcVa62mqrCIhAehIgKCHuPBjkInSSS44o9GfOmPZa+659+p9x1tnn1L/htjtefXn4C+l5wXSupCTAc7jJUk5LuIaK5q+b+BWfW8L0n6RNBNKUgMVGPrHlI116cpKBfbo+Groi978nnRRwJ7hnz6+/xluJE+1YJ2RatypLBkmNF1mq5z/9jDPPctdg7Yqli1L9BCpQBOIkYJaHzgUUVlzH83cUq0N3Bt6df1nCZecOS1kxjkFMtEuUqVCJjM4ln3mG2rNv79695hFu/7/mTik0HhHxLo4xC7tjj/3Psccdlz374k8/nv3utNcmxHQiy1SucrVLipYsXXbCS0MGhh+DWyr7979vvt65Ix5LD95Jx9r2+549gTGQU3zzfVMwLk4s9Tvz7HPPK1+l2iXUgXZhFRbLcZk0D2NJXKJ9aUnKukx6kVQtERCB5CMghUXyXVO1SAREIHMQYHLHKjYG6Cly55E5mpF+tdi/f9++N2x18T1tHn7spqbNWqaGwsJmgMcxafvVAtgmq9/dCwsVLV78orIVmPd+/OF7M3756cfd6XfVMv2ZzrQaFrSE+4sfLUVSWCDIwT8xE1OCi+7N9K1TBROewB33PfjwOeflvGDJgnlz5s58963QBhE0m7/37dsX972Yr0DhovQJuJP69uudCFli3nLnu7DgjU3uvm/U4Gf7EPw7/EDKLVi0RCmTR+XcunnDum+/2okA84iNfKXLV7r4zLPOOXfRJ3Nn7fntV56ruLccJkHLkSPHCWZo8lOsB1erfflVta+sf93p/zvjzG+//urLGVMmjt2wZuXyaMff++Cjj195TcObO7W6+9bwINnnXZArD23ZZRLAH7779ptoZZUsUz4guCRvvNcgWtl++/974oknHTjwzwGCbsdaxvm5cue99qYmd40bPrj/73aRQo87PscJJ7DA2sKgfI2LqWhlcq0qVbvk0nPPvyDXVrMYWvbZJx9HO0b705UA7zksgHF5iED66zjOzvuURTgcg8WitjAC3P+Fi5Uozc+MzUjxQDrD+pdYFRaMbweNmfzWSSefcuqsd9+a6voYnudHe/QdVKNO3fq4G7TH9o8X+/XqOm7488/61SXvhQULN7m3dbtL6za4nkVD5Fttbuw6P9CsSZkKB+NXMIbesmFtVAsLlOUPde7V9/pbmzajjhxrupr97e9t3JAxajw8MlFeXEEVssRYUi4WM9GFUVVEQASSm4AUFsl9fdU6ERCBjCHAhBCTYWdVEbPgIGOqm3nO+voro4bd1fKhR5nkVax6SW1WZcVbO4Rk9W+89Y5GTe5pYe44KjFhQ9A1cdSQQcMHPN0jkuKCFWHDJk3/8Ocfd//Q+o4brmai587P6rcW7Tp1v+6W2++2lXJ/j3nxuacnjRk+OFL9qMtzL02chvCQydrnm9bjSuHQdvX1NzVu3rZjVyaI70+f8uozXTs8gOImljazcrfrM8+PIFCvy7/bpEpNGtSu7CdAjKXcJMvDBBOf27iCIlBktACjTEYLW0LAG1gRbatPkwyJmpNZCJx97vk577y/bQf6pGd7PNYuvF70OfwWS8Dkxs1atm31SNdeCIb+tMAG9D0ci8B+zqrth1yhWTiDAyg1B/bp1nHuzHeme7F4/OlBw+l/zV350venvz4pNE+dq6+9oW3nns/kypPvQn5n5W7f7o+2De8Lr7qu0W30bfksAC356JOaXndZVdOe4FYj6obg/fbmD7RvYH15rrz5C3DAzh3btw548vEOH73z5hS/Amh3t34vvIQAPjTPbffc/yB99qCnuneKdPIWD3XsZsudj61So/blTmFBH/tQ5559i5a8qKw7dvb7M6YhzCOwrl95TmGxxsO6gvgit9x1X+v8BQsXg40JFB9HqRMVjE8GVlq36vB4LydcfG3cyCFPdXm4dSzlde49YAgKni+/2Pb521MmjeMYBK9tHu3W+4bGdzVnxTWrwt+Z+ur4Ho8+0NxLGQL3m+9s3rrVI4/3NPlpwJUZG0qv559+4rFY6qE86UIAF6UXWML1YVSlW0iNUPajrOBYxiiBoNvEitI78v8pFSt1UTmE9PRzIwY+09O+Zudv+nL7l53PY4/jl4N/8z+eLTPC2EP/Ft7fRrojcNSEsoI89Pl8Fi5e6qJhE6d/iHWXO5bnt0W7x7r7KSysH2rzUJdefY8/PkcOFJabzYoCBQaurZ5/+fW3XdnbP9+0IVLMHM5nxhRnDLXz01fy3lptrvAusHcFY9yHujzZb95H778damGSLnd86pyEeRzPC/FfsmrQ8dQhqVJEQAREQAREQAREQAQyjgAm9paqW3rY0i2WTgsGAM64SiXQmQeNeW2G8fq33/DxvkIpv+YwWRox+e3ZHO/Ssh2//OO+o3CIhAKhlssbagaPAGvAqElvhpbL91BlgVe5TB7dMViOhOZp2uLBR8LLc65hol0uJsVz1+z4kePnr//ql9FTP5i/cPOuP/gbYWO045N9P8+bpf9YqmjpWUu9Ld0Y4g7jCAS271hL9S21t1TBUnY9t8l+p2Rs+3r0Hzom0jN7c9Pmrdjf7vEn+0Wr6bBJb31E3iXbftxPn/DZlu/+DO9f3N+Lt+3ed+U1N97iVybHk7dqzTpXhuZ5oNMTT3mVSXlYZZAX9x+uD6fvfXfhui9cH/xY7/4vRmsH+4uUKF3mnQVrt3v14Uu/+PlApWo1L/UrB0WFO27cW7M/6zVg+Nj3F2/Y6X5D4eJ3LEJ6l69qrcvqku/25m3au/pz7plLN33t8qC4idQehH3kDe37EVRSp3COXK88+QugYI1rQ1HQ8uHOPULfc67sgkWK474n6sY14pg6V13TkMxYJY6fMWeR17UuVqpM+fACWRTwRP8ho13+yTMXrJo2d9lGdz+y4jtqJZQhXQjYNeEev8HSHZYOKeCinZx3p6VGlugDOlk6i/ej3pGHk2tyb6uHuO9ZTBKN6dHur3fDLbdzLp41yspfsEgxlNP8NuPT1VuxlkDpcFerdh39xqq4YSX/oq0/7EVx4ZTkKNOnz1uxObQP4BmPVGeOHfPGzE84hv67kFnhkR9lhRufOuXz0bY9vY+3Np1kifHkxZby6d5P7yug84mACGRVArKwyKpXXu0WARFIawJn2wlYWcqKNPyQp8gVRlpXMjOWj1uoGnWurFf7inrX4lZi1zdf7YylnigrXpry3scFzB4fy4jhA57qMXXCmBH44WUS+eBjPZ5u2qLtI6wyc755w8vFfQm/YeXAKjO3//72jz3BilhWL2MmzypWBEXXNGp856L5cz7yq58rj/3rVi5b4vJdfMmlV1Af/mb1LRNNAo1T3ot9ez0eqb24JRnyypsfIBhcOG/2zI6t7rqVFdM1L7+qwYBRr05npWwsvLJAHlan48qAuBSsCF0RxVc3bjJYlUgQUlzwsIruOJuYMlbCHQBBSvnO77hGwY8xf/PJqlVWtHNOVqKy+pRy2M/vzqUPf5PX5XEr9cjDb74r97SKNbnuWFbfYwmGm6TBz/To7NU6Zw3mXENFItDmjhuvRjDEyl6OQ4GBYL+juTbCLQ8WCwiUDtiyV1wU+fWB9Llu1e5P5k/KnRMFK9Zv/P36+FHDsAgocVG5igjlKfeKBg1vmj75lTFDJkz7gD74k9kz38XyAr/lCLro23AjFe0qwsVW6M6kDuZ6fdSi+4wAACAASURBVDsWFbgRYUnyE8++OAqFQwvrj/2sEVA6c4533pj8ChYQfKevfPGVae9T3/xm7eZXh8LFS17EPvr/xZ98PAvrAqcsWvDxrA96d2p7P6ugUWLwO1Yk1M+rPN4PpcpVrMI+Z2GB4rvf8HGv8y7hHLyfdmz7fDOrn1ES3G4uWZ587KH7ozFy+ynviX4vjuI+4jfeldMnjx9d/dK69VBql6l0cXV+s1vMN2j7eTlz5eadwvEEBmc1NvyLly5bAeuRF/v1NMuPj2ddVL5y1X/MnGb96hVLw+uHIovri+VF14fuv/P9t6a8ihJj7PRZC2FeuXrty6ZNGvtSLO0KCsAZN9EfHnKFpv4vFnox5YEr41PeNcSx8NzCFBG8s3j/sYofpRrvN6yeeGf+anlxXcf7jrEurlApG+tUl9jv3pe8Y6kD+7i+/I2rN46lPDbeo7xzt1viWO4H6srvvEP5zj3NOV1e6sR53fuVczgXkP+m1/3jrKqOxloqyCDqx8U1Lr2cTJ/O+fA93DD1H/HK1NPMog7L5IebN7nBudBjzOpVGFZ5jI2xkmt79y3XUo7L9735vcMKr9+wca+736IFEW/9aNcnWejz0+4fvm/W6Kpa9N8ci1vCr7/csT1/oSLFzjFFyE6z5IrauMyXgWfmaku4XH0781VPNRIBERCB5CQghUVyXle1SgREIOMJMAFjcpfPUsCth7bYCGAyjgCeideV19xwy9hhg6KuLsbAHosMBGVMtO6/7borQt0vvTx0YF8mZrh8qlStVh3ceXjVpkTpchX4HWGVM31H6XB3q/adEDC1adqo3mfzZn/Y5amBwxBmFSlRqkykVpUwoQ/7EUouWTB/Dt8RTPV4bugYBFpDnu3dDcVK3WtvvLXP4FETEBbSbr84FAiBnnnx5VfJs2Lxwk8eaNqovnMh5SalZ5vD8dhIJ32uk6yFrOzdZgkf+55+9kMo4LcZv964ysBtDf6961uCJ0IVBDW4eSMfLnaYwJaztNASft8RyPD3ektc6+2WrrFU0RKuwFZaYtyFuynOg7Bml6UtlnChQj5cDhDzhn3UAUUGypG9JhRCIMPvuCZwio1DMTnSSyBj59Z2lAR49juYj/GDfcCT3RDweBWJgJjfXfDtSKe1MBd7nQ9zyjVBcaDvWbl04af0ibFW2eT5BBYNbD/t3h2oF33gAx279+H7iIFP93yx35Nd+Y67D5fXvPiVemH81Pfog1HA4ArIuf5wLq2iubai/8OSDWXF0oXz57Zrdtv1TuhmN/6fL5gyF4UFwnMU1OHxNRDaFSpWMuA//u2pk8a7ulHGQ/fceh3WF1MnjvFd+Vy0xEGXT59vXL/2wsJFiz/as+/z/D3j9Ylju7W//y6nQLKyx6GwIPYIimYv5Q/WEtQRBhZwezHlYJGBsoL6tGl6Y71VSxcFfKE712DlLEBtrNeJa4yFTr2GNweUMvi9f7LTgy2oC66d2Ne593NDUIJce0lZ3Nx5bri+YgcKeu6TXgNHjENZgZuqB+5sVN+5xdq0bjX91xFb9UuvuBplFmw63N/0JheHhb/XrVq2BIUF7Yu1XZaPPpL3Kn03Qm0WLGy1/o/++JAQWv1dHEQPzwpf+gPeVbzrNvuUxLuHd2g+S7z7OA5lH1Y7p1vCNVR1S7yfUB64cQfXjDhQ7t2FoooxMO/QcOumYfYb9y+KCi93jYyhUVjw7nvDEkqN/JYQGvN+5N5A2ca7GPehuHGsEaznp/bJu5XFClhr8V51Sg3e1SgxUt21T8myFStb2dmWLvxkLp9puVW0WDGUP3/W+++0e7z3s/kKFi66bNGn8xinRos3g0Wc69OHm+uqUGWFq/M8UxTzHDPu5DfGnH7twZqYvob9KIqdssLld+8wApCnJZM0LJv7n3uNe1BzujQEraJFQAREIJSAFBa6H0RABEQg9Qkw8UKoyASNgW1gdZpNmFihxkQJIRQTbz6ZMDmho5uweQYGTsQJOi5N8hcqXOzpxx9pE6vfWqwYZr497XWCvrJqNxaFxd0t23WscHGNWigZwpUVXF7ObTKczSgsEKh5KSxQJDhzdbcfn77d+77wEhO2/j27PoqygvLWrly2GIUF/uEj3T7OfcYnsz941ykW2nfr0/8sUyrM+eDtN1FWuPJcOZTpp7C46Y5mLVm1i6Du4ftuvzE03oUtoGYilc2MS3x9qqf+rZ6pS0SQQtB7ePgJREIbQKwLlBFOOcGziaAGKw1WXvuNmQKuY0I2hDrXh/2GEPXW4G/z7BOhSui23f7I50ETxQjCIRSgoyytsUTgYH5HSIT1CHX+zfoXlBn4s6bvQRESEMpYcrE7AsKZKFYmHlVInZ98XIfQ57nk+FJnVtc66xT+RujEKlt+Q+gU2o9ybRGsudgvPAcIzehvKQdBJ/dCeL9Kfvpm1wc7YWia978IznHVgVL11ZdHvOBH2HSkgTaZTDyuQCrEzEHov/uH73bFG8+G/pFzIvD6zgTYWE/gZo7V/B+9O32qU1aQ51TrrFzdr2hww80I0bE4QEEc2ibnLsoMOyLGrzALitH00QjJH7zrpgbhioAvtm3ZRF9Of8xq3XABGopcF7vjr7DYEgjjRz7f98lId3Px0gfdHW1av2YldcGyBSu2bg+3vDs09hEKJlYlw+S/J558spfCwllXfPH55o0orLF8Q6CHFQLxkUKVPaw+5rzxCPaJL+GUFbwjn+vV5RHXtv+ZqY377mdJ4/ZXDLrXmj/rg3dQnFMm903zW+rX+XL7VgS+vhvWGMS/IMPoF/o/FR40/kRjw74//9gTj5CS5xHhMiv1uR4kFMUIpOn3UO7i9oZnmryB5zetx0dR+i/HyPUdzuIOYTt9EP0V/Rb9F8J8xn7sIx/7SM56gO+0zQlFOY58JPoDyqO/c/lcfwkHl9f1aYfiNoUI53lnoFygvEjjF/bT56JsIj/XkGNJ3F+BwMzB9tAmtzkrCbcvUhyV+0KO8/pKO9lg0ThKXhRvMy1xTFVLN1tikQJjgKmWUK7CHCsv3g+4Cp1jn9xTtBV2R/T98dxXxI0gthhWWPEoiaO0y3M3fSoKU6yJ6RMb3nbnvVjXYVkRTVlBgbiCOj7HCSfwfhhtsX28ToISnJgWjI0Zk27bspHFGJ5buy69+tEfvvXahJexRgvNRL+MJRd95hdbN3M9jtiCzxdjAe4l7juuB39zDzuLV993dDzXKcL52eWsXcOzMQZDQYaltMbYKblpdYwIiIAIpICAFBYpgKZDREAERCAGAkyMcAPFhB3BGYNuTOgRfjLgZR8DclZa88kEvXgwH6u1GaDzOyvJAq5mbECPIJJ9THaZYHEOJrAM4p1rGrfPTb4CK6OCeVy13WSav5n8sjlzferq3NUwSXSm/kzwKNsJQaMGWsTlEQFlEe480+3RB/+1yYqrQLTPD995M6CwcKszI03+WMl6b9sOATdKuCAJD2ztzmUyEwSX2Zg8eZ0/NKAqwhvy3HHfAw8jGFu+eMH8CS8NGeiO+9ekV3wngK1fWxB2FShyUPg3L1hemYpVqiGsZIVtTwteGl5epDJZyduifecnyNO/x2PtCbAdem78vvP31k0b1kXjm0X2c51Zjcn9zkpx9ywc0Xx7ttiHIIaJKNfWuZnYat8R1jihTWqgy+dRiJ9A2gXORECEOx76DfKGr0bl3p5oCRc0KEcmWEKxwXPrlBu0pZy1FUEg9wjCY/oU+grn8opJOc+/K98pV8OF+k7JENq/hCpGKMP1H5RNnRF4cRyCLliz4RqCPgX3ebhbYB99HsojuHOP0+ch5EARRF1xW0E96UsRjnHNsE6hHIRSBIPm3BzjruWP9p3VofSXrIDl3qD9CEY43xfBctjvVvQ6lyX2U+ptuCfChQ4losiNZHWwd+9ero9vn+VXK5Qh7Fvj4wokUmsKFD0Y98B0KasQMN3a7L42xELAjVSPR1o3Cz3WZHOBYNhsKAqmv/bKmHBlBfucInjrZv++CbdGlWvUvgwhWSdzY+UlaKc+Ju//E0H5aSYdDG9HqKL3bBPmxXvVnIK5qJnGsWL4KzNV6NDijps4b3hZxwRXHXsFoCZv6RB3UASh7m6BwPm9T+f2rUKVFfx2nEXe5dOEg4F3VLQNpQJ+6clHsPNQZQW/1b22kVOOmruYmYfcvHiVW75KtZr8joUefvdpa4cWTW+KpqzgmCbNWj+EOyncfg177qnAuyl0Kxy0QIzzneQElPQtCO7pE+g/YEQ/ns8SfQmLB7gHGDv9LyjwpL+AIWW4sRF9jhvncB357oT7TinqVt67vIyD6FvIS//AuemT2I91ghOqsp++DsUd1jH0HVj0OTeAKLwRpFMnVvzXsVTMEn0wfQ/jPPpA+ieUQ7ik5HyvWSImDH05imn6KhePhLrSV2Kdwz3FM8h7wilD6A9xU0nfQT+JAB//+8vsk42+9gpLtOkn+53nxClIKJvj9pkA+G/bR714V7jxK1YZru8OFnfo4y371iD8R/vbMffYlW2F/RjRStXrIPuNNjplRmgWWDvlGG2COdaNvBN4XzgXVFw33oew5jf2r7ZEe7nvuMYcH9fm3EGtjGCJEFeBETIzlmT32pVLFz/c/ann6H+feLjVPX7WeqFFMa7GhSi/vWAu3/z6MBbsOPeAjIH9Fh3xvnF9N64Cw6td32Jt8BvWH7iZi4EBzwf3J88ICkqeH55Jrjnfeb4YF/C88Xxwr7q5CuVzH9NnuP2U4xaPucUr9BW84xnbueeYc3Bujqcc990dy73M4hXuna8zavFHDPyURQREQASShoAUFklzKdUQERCBTEaASTQrqStZchNJJkCYFCMgwL0CLjuYwKLUYPB8nkcbEFAyWWQyiwDSrRrmdwbtDNYZVOezNMcSA2rKYWL/sSUEeUzGGHzzG4N8BvwM4AnUx0AddxEc51Y0MQF3/oGZ9DNZ5nj3ziBfxA1hCsqKn3/c/cP9ja+7wkvgE6mAJQvmzWFVKoKeilVr1MYfuV/++02Ij3IAP+FvvjqOVeiem1MumPcoz3efc++EoAbXKpz7jhYPPIxA8cmObVuETtb+d+bBFayRfIOjrHABDHExRf6WD3fpyefzT3XvhF9fV1FXXqQyb7rj3pa4GNmycd2aGVMmjg1vpPNj/kmIH2IvEDaxc0KZw4RwyTL5Clmpx0rKfJYQ3iMUinTfcs9zjyOw2GxpuiVW0yG8eN8Sk1/2MQFGYIPQh2eLZ5MJL8Jx8iK04nieaZRVYyzNscSKT/Yj2ML6geeYZxqF5Y2WeBbpFyg30sbk3WujDwg9/jb7mxRpQ1DD80+/gOCPtr1qibojsMkX3Icwn/axWhVhFufiWPo2hEMIfXDfQp+G8AluuMAhgC/uPuiPKBvFCX1PwGVPcHMuXxBKYknCPUk5uM2iLLdSfKR9p7+k30I4B0uEZzzLuAHh+tEGyqC+CAqpB+1D0OgUvNSXa0A+nj/qxbm3B/PSNsqkf+UYpwi2r6mzoazgeceFD77GI5X615+/B4Q7rNyN5+z4ESd/NJ/jXmU6C4uNa1Yux8XSPa0ffox8T3ft8IBzz+SOI0aC+44yovdj7VqGl4nFBKtr+d3PpQj9d8v2XQLWZhNHDR3kp3Rmf6R+HAu77Vs2bcA1Shlj8P701yfFyo064AaK/Cgr6O+7tbv/Lq8+nngghyw5bIWz1zlKljnoGgZFADEqsKqbOeON16Z5vKPOvyA344Jsu77+ivs+4kbbOvcZOJRMc2e+M71vtw6BmB1uw8UT8Svc35/NnxOwCvTaCIaNGy5Wade+sv513Ge48iLmSbR6wAA3i+R7oW/PLqHWfvyGAp2gu1yTFUv8XcmEnye4Uvor68dxj4fAmX6UxFiEPpOxEorZepZ4PnjGL7NEP8M4AcUl++lbXb9OH82zzliG/o1+jGMZk9En0YfVskS/wdgHQT/7UBLgPpL+Ds7Uybk+Ig/vgtDf7E/f7TqPPSg+XBBzhO1uY1wYbUO5wfm9YrLc43EwfV/A4sU23oW0ifEg4wEs93gv0b+SiEuxya4FjAhYD3MUJLCij6TPxFUnlgv0k4wxt1vCYoJ3IPm4HpyDewm+vNvIR9/LNUNZgTKE/pj+Dd701eznvJzTWddxvfiba8q7hrz0KZw7VDBN3ej/KZ97hecKTpyDfNSDMsmH4oiyaDsbihv20fcT84FYLZ7WdsH8R3w4hUU897tfWdF+R+lAHlzgoQT/4K2pkz+d+xFjlagbLtzIRD/7ztRXD7nOCz+wULESpZ07qGUL/fuEW+5q0YZjGac7t4SuLCxBmrft2JW/iR8XpXLw5lozJuE+5H5FScF9zvud54U+knECzyb9NeMF3uVYraK84z7m+rNYhfEDygXuQ/oFxoTcY9w/bpzHPck9y9iK+5Fz8SxyjLMg5DnhvmIMw71KH/CSPRfr7RmJW7Flx2oTAREQARGIkYAUFjGCUjYREAERiJMAkzUmkgx4mSgzCGcwziouZ/5/bUiZCDCZTIWvGmUQzcSYyQmJQTR53cZgmQE652GQzoSc8+GLm4koA2smYgz6OY6yELwyIWCgjlCPQT95mSQy+XYBEBmkM8ml7tTZrUwMOf2RXwkojbsKBBUtm1x35ca1q5iYxrWhJECYhxClfJXqNf0UFpjfm9soTP+z4Tc9ktsphG/k++3Xnz0DkDr/5fhOJ1/jZq3aYgr/6svDXwgXoCHoIU8kFyes0iUPAQYx1acdFateUhtf4QRbDQVyfq48gfIw5f/NrC/CYTFpRGHB72OGDHgm1D0Jv9W56pqGtSxIOcynvDJ6uB/soLICYQMTO1aCsnKMSd2pto97h+uMAA6hAfcRE0F3vyLkcMI5hEdMGg+t9D9af9BBRQMCiID1SrBst5LfmenzDJHHWQGEWgvx3bn5cS4qeH6492GKCwju4UBZVt9QhQ0ceL7gMscSz0HAf7/l4/nKFuIShPOwkp+JPt/dc+GsCuDFOdjnXIGQ363mdW10CpTRts9ZLzFZ5nllYgwH7gv6Ea4R1+JKSwhg+E6bcNGAcIp7mzbzPDMhR+GAkC7S5voRJ4Ajb+BZ8tloA/eFl4AsyqkCuxEShW+sdkRhisLGCbJgRxu4H+ECE4RNCJYQOCCogjnXhT4LayhW0cKKa8Ax3KfsQ2hB/+VWznIcArTA6mJLMOMaIWDjN4RVLkYIZbl70b4e/YYiAdcdKGOfNSupaCXagnv64GxnnnUOgrqYt7IVDyoSIvkc9yoMIfyFFoyCfeYVadltd7d8EOUKAWQ/NDd94cdUqlrzUvcbygovVySVgn7WsZzwC/5a97obb6VPZfUtAnO/hlI/BOXs91MWz/3w3bcQ6l96VYOGWNyF95V+ZRe0GByhwc1Rfrt3Qfgx51plXR1oV/j+HGYCYp61Aoo53je33Nm8NdYffbq0b+V1fhd3Y/vWzTwHvhuxmp4aPGoiDPAR3/mBe28Pb1/zhw4KB9l4jxJI26/AEheVDwg9ccOIwvubnV9+gT/7WG40rDiwVkTBH35v0P7OfQYElCpTXhk1zMWDiqXckDw8ezyX1B+rVJ5d+hDGVs7ii76IPpvf6CNR0vL8o7BxromckJ2iUYLy/mdfqOui0Kq5fpP+mT6hhaXtwQyhfaWzNOC3SFYEcTY7ruzx9MVOWcEJaBcJSw2eJ4SwKPcQBjM+CFjahrzz6CNpI2NU+kiYItCnj6afRJlNv811wTrEbexzQn8W3CBcDt3IzxiT83L8hrBjD40vguUwZiGxoVQI3+/GCa4uCKUZz9FW3r+01Sm9uV/4m3cm15p3C8+yU2aFVTX6n6WC8StSoiiOXvrhOYqY/zp+QVnBc874N5YysIhivEjeNyeNGxWpfwy1Ol7qo8RkYc9lV19zA+VNfnnEi6F1oE8fPmnGR9Tx7SmTxn1sMTFiqCP3BO9vEs8q727e/4zHGM+578yVGO/VssS9yfvcLUjIZ9/dQgXKY+zAeJbfKANFKM8t72DuD8YP3KdYT2DZ5MYF7rnmnNwfjLcYV7Cf8f2BoNKCemgTAREQARFIAwJSWKQBVBUpAiIgAkaAAS4TXyZ/TLIZ0LJKmQneTEtMjJjAIcBgMvimJYRTmOozEGbwzOAb4RGuXpg0I+icYwnlBEI+9nMMk0UEWkxeOR/+Yz+xxKpEzsd+VpoxqWfCyWpzJn0cwz5WIDGYZ2NS4FYXogyhngHBbpiAN5j98A8mL0/0HzIawVLPR9s0X796pXND4Jk/0o/LFy2Yj8ICdyR++YgjgTAfqwMXX8Ivr1vFGh6o1eV37isQqiEQuu2e+x/ELYmXq4vc+QowqcmGf3K/8zkXTU5Id0+bgyuV8fEePkl0Pt53WJwNrwlk5eq1LmOiidBr5ltvTA49Z9Wada7sPfglrAiysdoW1y1RYHMvcm0ZAyD0RQDBannuKYQw3HvObB4rIe433AdwHyMA4J5jwoegCCExwiQE+pSH4IHJP5NCJnbcb05JgBCE8rnXuOfZxzOCMMG5pGCFK8J657oBpRrl8Dsr3DgGgQMCQ45FME951CWfJe5r/mZCiVAFgSoTTfxoI5hg1TP3Nz7QaTv15dwcwwpQ2spKziOEkCE+kp0Q+zALFTuGLeDCx2fzyk/WwCr6oHCI5y+gKAlutA+BnVPM0BfAEX7UGeYDLPF8w4e6wYy+oXYwoVhBgE1eFB1dgmXPD/7On5zTWTNgHcFk3il7ODcbq5aPZqN+CAbgjkCJewom9IsIN+m7nNDBXVvH07nvoM3crxzHfUA5CDaoI+U4JQP7+c79ywYvJzjj+h62paZ10dXX39S4oK0s/8ksqLBIQLCOgsJije7p9szgkQHXSZNfGYO1FG7eEDbZtt9kxvt///2331jt7iqHhRrfWfmOtRaC5fC6h/9NXgT2CNKJtRMtf+h++hin2F2/evnSwWOnvosS2JQrgWCqoZuFSTjHxWnAcsBPuF+peq3AanHcIPm5HmnU5B7eb9mmvzZ+TLgVR+g58dnuVvz69ePTJo19iRXE5L3ksqsaECsoFgahwjmuQWisjvDjc+XNxzNmCuuveb8esRUvVaY8ygUUOAQJ5/uA3l0f9XPXUrhYSQRl2bZY7I5IdcVqkfcKFouPtbmnMf7lQ/NjXeGUVYHy7L0YyZ+9syrkvU3+of17d4/F/z15r7v59rv5fG3cS0NDFwrgF7//yAlv4CZm2+aN6ykzFv7hecJ80uPyhWeYfpl3AM86/RnjLMY99N30H7SDfgwhJ7/TXzAG4X3B+w33WLwXeN+FWnp5VZH3ktsQVPKuo3/iHch7hHfNbEv5LGFpgAUYK7Xpj3l/4rIHAS39DefD0oW+m7rQX9MfoaRFkcCiDtrFd96zzgUNZTuhOsJ++mXeZ07pAgP6Rvo7lE+0nz4THm41OO9GNpjRB2N95dwpOUUt5dGXwou6M4bwEsLSdupBG7j3AgqJ4LVy/WskJa/fvlDFRrC6gQ9Xpvst1r9dPriQ3PvcLVZhDMw71y2I4P2xyhI86WNpe/i5Quvl+b1EmfKVGDNGshCLWkgMGXiHOCUn2bHWi8WFG3kZUxNrgj4kkuUyeYuXLss9ba7q9vy2Ye0q5itHbNUvveJqnnncwq1fvQIlVmAjHk6nJ/u/gLKCgN7dzV1VpKb5xKBwCq09dq0YC7l7lDEl4zaef8aUPJfc2/TLPHc8By6OF2OhjyzxTPFscBzzHr5jSeEWSrj5FM/1OEtOCcr8g+eWMRLH0EbGFdSHd3Xc90kkDtonAiIgAiJwOAEpLHRHiIAIiEDaEGDwzOSTiRJCQrfyi0Gx87GLq4G3LSF4cxMrJrj8zeTcmUQzycKUmoE5EyknBGYwz3FMOlE+MJllP5N1JpNzLLEKiTowoHcTN/YxKeMdgK9iVtK5lWpHNfhudEez+wkciq/a9958HeFqijc3+UH45lfIVSYcZN+k0cOej3QiVnzmzJUnH3mYWIXnZWVt/uB5UDAQZ4KJ1pBne3fzEjJZTFuUQdm2RghCWLj4QSHU6uWLP0PpguUJViNeZvvODYtfeQi9KMtie0xxK3qp830Pdex2V8uHHmUC+mLfXo97uRsJbWvwWnM/cX8i1Ec4wr3GZJ3JHvcG9wqTO4QytSwxSeNeRLCOMAOBEPcJEzncKvAb9+C1lhDgbbeEmwvuR+5vJpUcg8DHWfsgMAgIY21DeIICiMkfgpZQQRErLlEiIIxCiMJKOerHRNOtcKUM6sa9j/UBGwIm6sZGPbgW3P8IJph88psT2iBQ4ty4kKBcfnfPaLCItP+IEDQS1k7Z4YR2VMgJtuG4PWQ1LIoZNgRLgyzRTyC0hSvP+ShLbgUhwiz6KZQACPDgwspVOHF9ETZz7REQuNWplIuVAtYL9C+cHyUr9wHKFc7BPUYZsEUggLADJSr3EvXgnnjKEvcN14381NP1k/b1MEsbr6C6AUVPlC2qgD9aAfHsR5j85KCRvi42XFkoQ0leZaPAMEOp31By7Pvrr4DCBgFVx179BhP0FCVwJJc9ZSpUqUb+dSuXL/Fa/R+pPU45TJ+HSyOUEu+/NeXVTetWh6+MznaprdJ1yoNRL/T3tIqgX6p1+dXXcM65H7wz3evcxLdwig/cQUWqn/XRgWcape6X2z/neT1i225KZPpYFLm49ItdYXHQIo7tjYkvj4wUNwmFFPkQyHvVwbWHGCSX1m1wfSR3hVjPwJlyIin47fV1YfMHD8ZqGjbg6R7hq7i55q06dO0VWh8/IaPLU9h8R7nvxOuYMXUSgrqoG+942oii4v3pU1iZH9hwRdVzwPCxvM+w1sAdZAqtK46oQ0j/SH+4z/o7+g36QPoY+iNn7ca4hncDyb1L2Md7hP4GYeYUSzxbKDHo/1C657NEH0b/6RaYkJf+jzEVmxsf0X8yrqMP4n1CWS8Hv1Mn+ktWm9Nfk1ikwiebs7BzZfG3c8fp+j+OAD0Z2gAAIABJREFUd0J8N1d3wn6nQOZvZ2lCubSVYyiDOruFAdTVlU97eMfea4l7FxdC9NmBsWQwbsUXwXFCsLqHfXAO2kv94HZU40WvE6Tnb0FFtVNyu+uToioQSw0lNAtnYrXqStGJ7CBbfJMXZbc7fvzIF56LtawaderiSi0bgbF3//BdwHrUbytXqWoN9tkYdqGfW1dX3qx3p6O0C7iCe6Bj9z5Va11Wl79RpvTo0PreWJTtMbSBa+WUT6F9r3tuaA/jF+55nhvyc115PvmNfc5aiHJQZDCuYXzlxlaURT/BPU5/wHFYIDEeRiHJeIY+gueGcUlCPwMxMFcWERABEchQAlJYZCh+nVwERCCJCTDgZSDsVgAd4zOwZSIZKlRjEH3Yqskgo0PxDnyYbbUJPCvtQjdWBDmhjpfA79CK79QYdCMwwfUFFZgw8kVWGR7VhislCkBxwArV8OC0CEfwjc7vXu5KQk/Oak+EZ/zmJRTCdzkrmBHw4QP92eHjp2DN8MrIwUdMBHEThcCGsnDv5NdItwJu45pVyxuH+Pr2yu8UIJst0K3Xflax8bubFCIEa92h65MEBGciOOjJ7p28gt16lRW81k4AE8gSVFghNEbQ4dwqcS+iYOATgSWCGASGCEJYEcp9i6KB1fusNiMfQm/KYKKHggIFAlYoCOSYNHIM38mLsAdBufM/7KwinDIFIQoKC5RDTBJR1CFgYj+KkVCFBQIr6o2QHSE8dQ11sYbgnXOyuo56oJCgHJ4Pp5BhdTMWTgjinVWRfU2MLUygR6VDBTCh3w+5RLPrTvvdhJsVwIFnJLihUO1tiQk814IxI/vhDB+EV3y6saQTBDjrBvc7f4cK1ijvCEFJFIVNQlyEbdZ34JoD4fKpJrxi5boFLT0FZSmulehfcPl2rHVo9Gl88o2+ycW74Sf6PFJoo7Emc383rlez4rpVywOWTeGbC8a63JTG8UIL9cF+e/PW7RBSDTWlrVc5DW649Q5+x13UBot34ZWnfOVql7j4G7Pee+sNrzy1zZUdv1OGlzI59BjXNizRIgnChz3X5wkUFlgb4IYvWqwQzuFcAiKEnzh6aEQFuFPsWNgOT4sIF/TcXUNcU/m5K8RPPOdHyLlhzQpfi0Rin7CSGSXJyOf7PhnOEsserh/nYYU3dYz0fuJ4Yky4ciaOGjIo1lhTvI9432M1g5UJcUqat+3w+A233dWc+5d3bIcWtzfa9c1XTnka760YNX9Yf+GE907o+Lv1be7cAWGmyx+yqp5+j/cGG9+xOAtcCktOqXCoHhH6p1Dltp+iOxbFaajgM9QSwc8yL5xRqFVg6HcU/IHN2s6YkHekW6lOvf4KHf+57+HttWOpH+97hNi8k/H375QdUa9Xsmdwz/yqZYsWpHVbzX3dIatjFtjE6naVd0z5KtVqUr/Z78/g/e67YW3nFgtFci3o+mSU3M8MeXnyZfWuu5G+AUs5+r0Zrx8Zby0lfCI8fxTnnh23uMPrOQxdLOaqEMkiljz0I3wyRmURDkoS3stYaESyJEpJE3WMCIiACIiABwEpLHRbiIAIiEDaEGBFDhNmBL7psvkM6NNt9Q+rKnHDgUuJebM+wK/8UW22yBilT2CzxWSnhrsAqVTtoKsRfOv6uQdxx1euUesyvhMQcPf3u45wCeOERp9v3LC2Wu3Lr8JF0yALjI0pfHgjnLAKAZOfQIjJHooNhEc/2PkQJrHq18u3McJKNzH0mni6wKic77+2rG78jDmLXMBFlCtd2ja/I17XL+FtCq6oRMgRKujAfQ9CCTYEOCSUYs4aB0EISgf8AnPcq5ZwIYBAG8ERE3cmeAhcKAuFBJZAKF8QlOO6jL+xvmClG4oOFCNMpFH2ofAgYVXBqk4mnNzPsyyh6OC8rPBHCMP5+M4qWueOikk9q6Y5doylRZZQdKDM2M9qUvsMbDYpZRKKFQurFqnTEQIrlzeZPo1B6KTbrTR1TYwmZDvCbVYYGz+/zunWJ6X3tcLl0UvP90PJc2hDaD155oKAIrLHI62bve0T5BQhDwJp2+wxP+VUFBykDk88M5D+CIG+6Tv++t5cvhHg2q9tpctXClgZLV+8wAlgY8ZQunzlwLH/syX/nBOXIVgshBdAf+XOg29yvxNcXv+6RuzDQoMV/F75nMuoWe/N8FRohB5TuXrtQD++dsVSnmXfbdXSRQuclcVdrdp1jKawwFKEQNsUiGuraO5VcPlE3jUrlnjWw1lYkAd3WdTHr7JOsb3DLP+83jcchzD08vrXB1gO7NOtY7hiwQwIT2xjq5rZj2WjUzxt3eR/n7BC28Vi4r7FTVmsN4oTUqIYadu55zM3N23eijqweGDssEH9Bj/do3N4EO5Yy06tfB4K3EDRIavq+TO0L/JTGKRWlTJLOSiLedYYo/4U52IV3o+8V+n7eXegwJbg1iC4/nBlhGc9tW4AZ+FFedNfi/25pU8//vgcgdhVn82fw5jLd7uifsOb3M5VSz/z7L+IYeMsl9t17Y0VeDbiEE146cWBLKDxizOUWhzSsRzGsIxZGaM6y6p0PL1OJQIiIAJZl4AUFln32qvlIiACaUeACRzuaxD4IUTF/36ar7pKu+bEVrKbsG1at2aln6/y2Eo6mOukU07BOiWwebk2cSvaFn/yMQLsiFtN82VOho8tIKtXRies2rh25fLGzVq2RQHy6phhg73yFgiubkOo5bfKt0hQ+PXVju1br7ruptuYJA4f8FQPr/JwJeAmkRvMGiM8T/FSZQPCMYRq/YaNCwS+/farnTuGWXlMVmNdFRuNURSFF8EFw1d6sjrNrdJDwM9+3P4wIWb1vXNZhLUF+/idxOpllAXOhQfCD54Vt7rfufpBMeLiNbhzc4zzL40iw7nHCG/eVfbDQ5awsnjX0ljOEUE4g8UMCQsMXIbFuqo1Glbtz8IEUEL0eG7omHPPvyDXR+bOzU9ZASKUmyh7SfQ/BFXm9wY33tYUQRMC/REDn+4ZCSdu4kqY33HKijfwK3V1gu4SZcpVREHqdz4Ch1MP+mU/ywkUsbiNIt/MGdNCA/Ee1gR3zsWfzo3Yj2Op4d4xBNaOdlvR32JlgSs++ncvt1aujLwXFiqCwJ2/cWESqWyuJQob+t2VSxbS3x22YX1HHn6MJRiuxa8IWFiYi3hPixn23fvgowFXUCih5s480rUWbgE5J8JCFAYT350XsNSwGN6+iq0CIbGhZlucj3iEi8WCCpvrbrkj4Jee+w1FyYv9enWNpuyJdt20P80JsHiA2E1YbPkFHverhLP+3W4ZjnCtmeY1z8QnKF2u0sU8B1gdpXU1bW1QoM+gf0EhGuv5sCQm748WX8lZMPsdW6/hzU3cPr8FMXkvLIjFa2DD0mry2JEvvj5+1DCsk2OtU4Lkc67WsC6in0ZxoU0EREAERCAdCEhhkQ6QdQoREIEsSQAXNriWwVUOq8GTdlWxu7q4heA7K4BT44qffc55+NPPhvIDQUx4mU7gsj6CGw2OwfLDrWKd/Z63GbyFpDgYgNOEdhUurlGL2BV+yggXbyKSGX6hogeFULiIuemOZi1Z4esnQHTlMYn0Cpidt0AhfE4HNlxtTBj14sD335wyKb1XsEYIikjV3CrLcBdn7Iu2Ej/S7RJtlf8RqzuDLj+Ix4FrKAQsWHn8E2UlKc8pfs15Zo+wwEmN+1llZD0Czdo80rmmxXDAsqtnxwfvSwkBczMe6E/NwxTK74hbsdJlymOlgVVEpODVXoVcWKhocRd8GcUHsSu8rCtwK1K/4S23U8aSBfPnEGvDq7wKVarXJD4D+z4K+jcPz8c7A0UEypFobk2ubHDDzShtUZJ8MvsDlJARN/pb3FVVqlbz0hsa39m8T+f2rfwOsO46EL8CgePcmZGVIQS2Ji+uWLwsIpwinTxvTZk4FvdVkSrqrPsIcu6VD4s+5xJwkFlXhOfBZ/zdrdt34ncUTHabYLGWjcDhfkHB2e8UJXx/b1rs8aZQbDlBJe/lGVMmjJ3w0pCBXvdKtGuk/elOgHk/Vkq857jn43UbhxtF3pX5LJWzxAKKaO/odG9kep/wxJNOOpnnCYvXePvdlNTVjWcD1sVxKAdyW7wgzrdx3WpcevpuWL25RTwozv3adP4FebCAzbZl47o1t9atUS6V4lSkBElaH8NzQ8wWrPBYjEMcMG0iIAIiIALpQMBvZWI6nFqnEAEREIGkJsAqcHz9M9DFDU3Sby4IoHk0wfXPUW/OrYbFmWUl/WEbQhMLXxGYLOGWItLJGjS6rSn7UQYgYPPK6yaACKNQVEyK4MO8YJFiAf/BkSZ9LuA2wigCqr40+NnD3MSE1sG5mPIrjwCL5Gfl2m1X1yiPT+D0VlYc9cVMpwKC/oadyyrOilAG1xfRNp7TSy3Vt4Rf99Ayoh2r/SJwBAHizNz/cOcerILt1PruW+MRLIUWhm9w/j4xJMiqH24XhyGayySv4531gts3arB3IO1LLqtbH1dV5Jv34bsz/OpS5+prcLGWjbgUBAv3ymfyLgSn2b4xf1FeSunQY1w/Pu/D92bEGsh58ssjXqCMutc2upXYCn51RejPPgRvXi4DQ4+7osFBVylYzHiVV9LcN/E7yo8xLz73dKRHgzoRh4g8XtZ1/N7ojnvuDwRRNwuMcF/yKJZ6Dhg2FiUSq6DHDn/+WdeWnTu2bfWLm0G5TlECd9xnRapn6L4zTAnlLAIbVL+oYO/H2rWUsiJWehmej3k/CjfixuDSMd4YI8S+wloYy8dDcRQyvFUZXIGLyleuikVZStzwxVt1FNJ58x+0bJjtExfIr0ynkN75xdZAfDi/rWmLBx9x+/ziE7H/f2ecERhb7fn111+SWFlBE3l34GqU+x63oygttImACIiACKQDASks0gGyTiECIpDlCNC34g4Hv/isZrvGUtILQH/+cfcPXGlbNBsISH20m3Pj5BXwDx/vTNw4RyRB4H9PPPGk629t2ox8U14ZPdxrUsUqYJQK5CGI95QJo4dHWiUXm4XFwWCmlIdVxGfzZhPQ2HM7pABZu8pz1ZutmA1MCn82yeXRMs0ix2PNRGDpzyyxGpQV6qFBpw/DYEoOnleUFSiGXDDwLIJKzUwLAqxO7TVwxDgEzf2e6PhQpKCl0c7/k5lekYc4PtHy5gtaY20w13bR8obvL12uYhX32yLzb+7nQqn+jQeDbSMM94s7QbuxLCGflwsjdx4zBgj0u9GUORdVqFzVxe2ZNGa4p6s+r/bOMfdJKHyII+KO98pnBnYBCwu/QObuGGITVTEXUyihPpjxxmSvspyLq2W2+jlaEPF85orKCf+9eKOQwLKE8/D+Cj9fm47dehM4GzdixDKiXk75vuvrr3D747sVLnYwZsenc2a+F48LR/c+4li9k+J9yjI8P24XEbyyoIaYMvjjj2dDUOssPnmn+sUpiqfMhM9b3qzJaER6KCwKmDmwU77Sv8UDz8bNxCAJuITyO65yjdqX4UrP7V8TIV7QCTbAJp+Xy9Z46pUAeeGGYpn4L4wpGV9qEwEREAERSAcCUlikA2SdQgREIMsRQGBK/8qEEGGp+zupQZjlOAGZAy6Yzgq6c0ppgynDBWN9d9rkI3yK/9ds8CkbP+KRVuY2ur3Z/QirUFS8Pn70MK/6uJWmrryJo4YM8qs3yg23unjz+rWBQLrhG4oU4lK438ePeL5/JA7OwsIvgPehSeHefUfjWimllyIRj3PKwR1WeZRnuCqLpDDk+cTcHwHfTEtc16R34ZaIFzYR6oyyYuiEN2eiLMUqKh4Bu1f7zCVUwEVZztx580Vrv3PVs2XDuiOs0qIdG2ph8dr4UUO98ucw6zknzEI45+dyqGjJi8q5OA4fm0WE37lhxL49v/7i6VbKHXdP64cf4zsWEEsWzJsTrS1uPwL8VcsOBrwuUvygFYXX5tyfbNvsbQnijrnlzvta45Zq9vszpu365qsjVqejqCle+mDMIb/YHqHnd+8eYhJ5xZAguDWBbXnPcc7QY6++/qbGtzdv057fcHeFOxq+u3vAq37ueOrpFBvxCj1drA/ceME31muhfJmGAO9ChK9XWIrXFz+LcJxlBe9MuZY2CLid4+ouXTh/blpfZefKjb6KfiOe87ln98CBfzxjdGGp1bFHX2KMHdoixeSwbilQzr/WF8RTjwTMiztGFMco7LBOCbTXx01qAjZPVRYBERCBzEtACovMe21UMxEQgcQlgLCTGBYImFdbyhIr41mpid9sTONvvvNeX3/h0S4rwpTHevd/kXzrV69YGmmFF+diFapXmSgqnG/vaRPHvuQVH4LjWKHqjkd4883OL/HT7LkVKFKsBDt+N8ftfsK6AoWLFKde5Ntt0sYP3vJeict+6k5AXb77BUjNQpPCaLdGrPsRwlSyhOk+gcGxdopm4YSp/yWWGlnCz3O0/LHWRfmyEAFW14+Y/PZslJoIrPt08Y+bECsW188QY8L1K37Hur4kWkDV8ONPsc4yv5l68TsK4Hkfvf+21zkqV69ZB6UF+yIFe60TDLaN66ZYgn87pazXOVm9XKPOlfXYN3Jg316xcnP53GriU047jXfyEds55+W8wCmhI1l6YF1x6133tcGyZLSPqycYYv3HST6ZPTNqnA0nfEQR41W3cpWr0Sdl27xh7WrnGoy/cZfYrd8LL/F92qSxL705efxod3yuoJ96Z/HoVW7OXHnyOReOC+bE7g6KsvQ+ivcOzFT5GZsSDwwlHlZYvB/j2VBQ4EqKDWVVlneN46y3iPUQaewYD+RIeU0ZHLAGW7Fk4Sfxluli7px7fs5cXsfeeX/bDvkKFi4aquz0W0jD8d/v+gZrg2woVeOtS4Ll/83qS3/uLBc95xwJ1iZVVwREQAQSgoAUFglxmVRJERCBBCSAsqK6pQqWEJgm+wqkbAinpr06LhCM7u6W7To6C4l4r9397R97wglqnu3xWGAFafiG8Ma5dwq1ZgjN175bn/6mszgD5cKQ/r27+dWjQNHih3wxT7EV0ZHqawqLQF5zD77FtzwLkur2TX91/OhIvn2ZHDrz/i+3f+5ZZhaaFMZ7q/jlR9nA6mdc3KC8QAEV6fkjPxNQBJq4y9AmAnETaHjbnfeOmPzObARYCPw7tbr7VlbGx11Q2AEmPAq49mF1bGigZK9ynWWbdcUIWA5tFateUrvJva0e8qsL/S2KYvYT0BoXQ155a1x6UHGA0P6jd6Z7xnBgvwsSvcKsMCL1fxZWKBDfCSG7O3/oeXGX1KXPgIC1Byt9CQTuVS9cRt3T5uHHvOJU5A26yfph17eB4OXhm4s3xO9OGeOV7+FuTz2H9dz706dM8nMdVaJMuYoci5Ipmjso8jkrh22fH7SOCN/MY1Rxftu0bs1Ktw9rkIGjXp0OG5RBxJBw+2g/7zz+juTW0Ak9v9y+dQtKda9z+/32/a5vA0JKzuWUM/Ecr7wZSoD3IUoKLJq47vFaEvJeHWmJAPGMV7K8Yr+GxfRBkRzJ7WdqXvHCJUoFLMW2bt6wLt5ynavAarUvvyp8oQ+K4RbtOnWnzPmzPniHTyyofvn5J+KWeG5OMZ47X4GCXn0n1mj1Gt7c5PmXX38bhXu89c1E+XlOUETTt2LVIsuyTHRxVBUREIHkJiCFRXJfX7VOBEQg4wgwIUT4iV983AMFVtwn+zaoT9eOCEGYwD0/ZvIM3FbE0+a7WrXreO+Djz7OMawa9TOxRwi2buXyJeSrc/W1geCuoVvda2+89ZpGje/kt6e7PvJAJJ+9zsIC8/qF82bjEsh3c+6bdtlSOr9MrjyEem/Y6tfI5R1UgJhO5Re3+i08v5sU2nzvkCVIaB7zjnXyvQ906PLcSxOnYdIfD+8kzYurCtxdBNzN2LYphnZ+ZHlYQTcnmJJewRgDE2WJgQBKgn7Dxr3++NODhqNUeHfaaxPaNbvt+tTy603fhdKVqkSKw8D+HDlyBFy8uOCqfK9So/blL77yxvsPde7V10/AXOHiGrVcU2e+Pe01v2azsp99BHh2itTwvJzbCeJXmZIhEsINa1Ys279/3z5iCJWtVLVGeN4OPZ4ZhFIXBUq39i3v9iury1MDh7Xu0PXJJs0OV8rUvPyqBuWsXBRHiz6dO8vreBeonH0uBkh4PlYeYzWC1UK/Jzq186uHuz7LF306L4Zb51Dg653bt3kGwT09GL/IxTExd1MVnAUPK7rb39u4IfzcuU444YSA9Qubn9KJfUWOQuj5oyk4nBtGc2nl+U7ClVW/4eOnXF7/eizWtGUeArwTcV+EBSJjhXgVqlhncI+h9MBVXZaXI9zQ+K7mXF76OsZiKAK8lK+pcQtQbhFTWFJWJMtjv3OhSCdeDbHVOvbqN9iNFxlDDxrz2gyUkChBXdwhzhepLbwHsCrBWuvmpv9vVY2ighhGk96bv5xYTihITj711EReDMI8DktoFrYw75B71tS4oVWGCIiACMRAQL4nY4CkLCIgAiKQAgLn2jH4+2UFWr6sMrFDkHHvTfVqDzJlBStBnxw0cvy1N99+9/gRg/t/Ovej9/18XhcpUbpMuy69+jmrDILUPtWlfetI3Iltgd/1pi0efGTRJ3M+coFtL63b4Pon+g8JuMjAXcZbr0142a8cJmP5LIoh+6dOGDMCv9yRzukCbkdyt+FWki3+ZO4slDdHW96Hb097/cHHejxd0fwklypbofLq5UsIJp0N/++wRVmBwA93JtmPz358pBXNKbiPE/EQVsIFfErbxorQPVEaweo5JqCsYmZSinuD7ZbiXX2aiKxU5xQQQBBui0//rlbr8ro3NL6zOSvvee5e7NvrcT93QSk4zaFDWK2PsJrkFXzZZfxx9/ffoUChDxw7bFA/hEZ9Bo+agGCKejnFR3hdyla6GGvAgOJ07sx33/KqK2VcWPjgKtlIcSnOvyB3HgRW5Nu2JXJMCJS0H9v5EJh17vPckBa3Xns5ihCORwGBMBDFb69ObVtEKmvR/LkfoUxu+XDnHlgM0D9jVdL4npZtqcf01ye87OfvvWjJgwG32erdcMvtY4cPeta5duG63tf20a64FuTd0P3hlnfvNhMDv2tZvHQ5LCqzrV2xbHG0640ljovz8ccfezz7KBfXAqVT42Yt27Zo91h3FEK0r9XtDa8Kt46AJ/U78+xzz6tx2VX1Z0yZNI5rGl6XIiUOupVZs3zpomj1DN8Ph1nvTp8KKxQ57Zbedr17b1oc73LN23bsWuuKetce5BB/+fHWR/njIrDfcmPxi2IT5QMpng1FBSv7v7eEW6l4FR7xnCvT58Wyq2zFg31nt76DR5JcpRnr7jdt4sH/7zv4ad8OfbffDtvPPtuwX6OvRblMnKBBfbp1dGVekCffhfzOc56SZ5cx4mvjRg2lL8Ei8LJ61924f9/evfQXnAPL5S5tm9/hzsfCI1zm+cXDoW9+bfxLQx/o2L1P2849n+G9iGUXMYxQilAO53zysYfuX7X0YCyhBN1Q7rlA23IHlaAXUdUWARFITAJSWCTmdVOtRUAEMj8BhAQIQPNYYmVnlhF+Mrm5q+EV1RFc3HbP/Q8SkJCE4GTDmpXLEb45QczZ5ky3hAnhWEXrLiluP3o80roZ8TAiXWbcTzVp3qbdBbnz5h85+Z05Cz6e9cGJttKLFbUcx0rnnh0fvC9SGQj3WBXHuV5/JbI7KMpxMSwsvrivIsK5qBpnSppot2nBoDuqSOURzBxlD8Fuh7/69qzFn3482+az2VFeuJXUn29av7ZT63tuixSAPFpdkmQ/CsITg23hGcRyIppQxSkVscxgUspxWeZ5TZLrnm7NwJ3OAHPJE3pChDHEq6B/S4uKoIxFWRHaT3qd57N5cz5EkIzwCCGSi3nxwVtTJw9++olA4OrwjRXBLvjztEnjRvmtzEdZ4dyIzJ/1fsBliNdmMv5Dq/y/2bnDNx6QO3bYgKd7XGKCLhS9U2YtWotrFZQPtBXLiGe6PfrgjNcnjo3E9eWhA/tizYdFQs/nhh2moIZdv+6PBhQXXluRoE/49atXLkPgPvHd+cs+nfPhe+StVO2SSxHmIZDv+egDzf2UOeSFdeFiJUrzHeuHaPdBqCtDM4zxDH5MgHEsO1D+45KKMhEqtmxy/ZUuyHb4eV55achArj3vi2dHvDL1vlsa1AnP4ywsPjNFf7R6eu1HSHm1uXpBIfbahwtXb920YR2ut5x1IcLZMUMGPMN1SUn5Oib1CSz/8leUiPksoaTAFRsWhfG6tiE/gaWxGCaWBQqQLLuhPEAxwbOPS1QWwByX3f6zARrWCgdd1B3qDuPm9EeYaz9nXfGWKWBTujBl8DNPdM57YcHCuO1Daeoqtcyswp54uNU9zqIXpe35uXLnxS2dn8KCY1GMFy9VpjzKD+fKld+xDJxiY+rxI154LpJ7urihZNwBa+3UuA3Fok3jw4y7DjqzCIhAFiMghUUWu+BqrgiIQLoQQADKoBbB50ZL+DzNUhuTtwFPPt5h8ssjXmQlV72GtzQhaCmuR0LdjzgoCISWmCAeIQeKh1hgoWRoe9fN1yCUQfjj/Kaz+nTYgKd6TBo97Plo5bBCjNVqz/bo1C40qKnXcaz6PdZmoOxbaUIwv7IR+OHOyvkBjlQHZ5LvrEP88nY3dyhDJ745E6GeC0BLXvwYjxs+uD8TWD/rlWgMknA/rgd4/vhEARHRaqZs7lP/MWEOLndWWMJ3f8BHuzYR8CJgHjX+ou+hz8Kyiz4u1j4rpURft9g6Nza56741Qesqv3IG9+3RpYQF/sa1EUI03H9MtH5w0FPdAxYCXseVrVy1BvEQUCKP8QkmzXEWGiEQWBWB1vrVK/Bh77l9afvpi362DpVg0dHaTFDXzg/c24TVyQT/RvDFMds2b1z/VNdH2iyaH12oTswIE+LXpQys9dzxUyaMHv7qmBEv+An3OJ/Fn76Q/N3atbizr7n2Qph31XWNbnP1pr1PmAI2m5X8AAAgAElEQVQd5UGktpxlig3nxz2SC0JXBtYRcEKoaWFKPMcIU18ZMxwlABYof9vSbFy6DO3fp7ufALHX+MXHDO1+57Mo8a+/5Y573MKA0HoTIBfLDgJ9Exck2vXx2o/bmOd6dn64bZdefXknOatC7rf3LMbHqMHP9oklhkdKzq1jjooAK8VRUrGIZrclxqrxCl+32jG4luJdecgd2VHVKkEPRrF5ceHzTvrn33/+CR9/odxFeXuCmcLiKtD+ncjf9LX27wT7fkJ2+2KPv6k4smdHu5EtGEeIMSSxYnjOQtHs2Pb5ZizsBj/d3VP5HAtG3l1tmt5YD8W7GReXMEOPvZvWrV4Z/rwO7d+7+8U161yxZMH8iP0e7X6kxR2NcIdH30u7WUCDdUgSjUlR0BHzBVew21LwzMRyaZRHBERABETAg0CWD5alu0IEREAEUpuACT/pW/F52ic4IZxon2+bYDTe1WypXbUMLY/VWsVLlS1vcp2cp5x6+unHmALgt19//hm3SQhOIgX3i1RxBHNlKlSpZjKYPN9/t+ubVUs/WxDNOiOlIFC6YOqOv+LUCKiLhQSBdDeZ0M7LdUdoPRFsVa5e67JcefJfiI8BfBgj7EtpW5LxOHv2aFYBS49YusTSw5bet3TAnj/fJttxuLphtSHBillJF7DKiHRMMvJTm2IjgKLxgEljUHjGdsTR58JPuF+cm9DSUayem/OC3AjGTI7/ZaRYBhxHwOs77mvT/t03XpuAkMmvpqwern1l/esQRkUTRrPS9geLqI2ALdaWY+nGcaz65Z1A/5YSvhyPciZaf0q9cBs1/NUZs3CjdFm5QufTH9e9rtGtpsMoyPvIXBotXvTJ3I+iuQp0bcQVlx22e9lnn3wcS7uJ9XG8XSh8wUfLb8qIw7J0aRKI7x3YUFTYB8nFFPjnrTFPn9DgzkfdamD2/WPH/INSpXPv54Zg/cC1jHbeSPtzmranXJVql6D4+frLHdtR6vi5HTua8+jYoydg7zgWW+C+yFn9/mXvtx9iLTn4bnXZEeCiAA30f3pPxkpR+RKNQPC+Z3xY1RLuAFH4oazTfZ9oF1P1FQERSEgCUlgk5GVTpUVABDIzgeAA9wyrI8Gjc1pCcbGKldyZud6qmwgkOoHgs4cPBoQyBITF7UXAT3cUhQXuoLDIwEc3K081GU30m0H1TxcCQWH5YecywXi6KXKOppG3N2/Tvt3jT/bD1VPbu2++5mjKSutj/RQWIcoKhMgIpVG2krgGKDBYVc8+fqN/y5Yo1yetmWal8u3dyD1AjCbclmHRs8neibh10iYCIuBDIDimxAqP5wYXh7j6DczlpKjTbSMCIiACaU9ALqHSnrHOIAIikDUJMKB1wTkRmEpZkTXvA7U6/QngVxuBDMK5gIAu2mYTzz02MSVvtHgX0YrSfhHIEgSCAnS38OmQa5lEEoYXK1WmHBcrEYJDh1pUuBssqKwgCCwJC076Lz7deAOlRcC6wpJTaPzNcYl0nbLEA5X2jURxVTh4f5xrn7hA1CYCIhCdAO59sRbc6fpWKSuiQ1MOERABEUgNAlJYpAZFlSECIiACRxJAgPCNpQ2WvhcgERCBdCPglA74HI55pXdWd9mWbldHJ0p4AiHKisOer0QTghctUbosF2PtyqVRXTJl0ouGBQVjDT5R1Ia7neT68DtKC+Z8zuLigF1DXETF3D9m0varWrET4Ppvt4Ti6jd73+2N/VDlFIEsTQCFBQta9Mxk6dtAjRcBEcgIAlJYZAR1nVMERCArEMAtDX5OWZGDX3xtIiAC6UPACeFYVSzLpvRhftRnCXEt5ClE9VphftQnVQEpIhC8FqHXKeEE3wTCzWvByQEQSwyJFIFKw4PseXHKhxx2mt/tmkSKkfWv5UeRi7D6xGC/+Jf99rcdJ6uyNLxOmahoFFfbLfGZpYNlZ6JroqpkcgJBS4q/zQJXY8lMfq1UPREQgeQk4IKzJWfr1CoREAERyDgCe+zU+Dv93JIEAjFcBwuwekxYypaOMW1jqKGyJBABnrlDQhmZ7yfMlUs4wXfCkFVFDyNQuHipiwhQvvOLbZ8TYDuR8ASVFczhTrKE9URUATQBty0fSg0E1iguUHT8xysGSSKxUF1jJsB1/8PehQTblvA1ZmzKKAKBeBX/BJNiV+iGEAEREIF0JCALi3SErVOJgAhkKQIoLLZYknVF8LL7KB8Qtjg/6OREkMKG4JJJNZ8SYmapRyfljQ1RTOieSTnGNDsyPHBwyInkUz/NqKtgLwLFSgbjVySmOyjemc7CAkF0rIsiyIdbExfPgjIOxR/RnZK8BKSkSN5rq5aJgAiIgAiIQLISkIVFsl5ZtUsERCCjCSBEwO9prIKEjK5vRpzfKSuc8MT9zacLJOqsLjKifjqnCIiACIhAEhIoWjIYv2LFsoSKXxG0iOAdiYXECZYYa8S0BWNWuDEJi9Y4PnvQYiOmMpRJBERABERABERABERABNKDgCws0oOyziECIpClCARXecvkPvJVd1YVKCuyB4UvuLUg7odb9Ykwhe/8bgYa/zqLi8NKPuaYUAONLHWrqbEikAwEtMI7Ga5igrWheOmyFajymhVLFyVY1XleeGcSi4JYWXEtPsM1lCkoeKeyKIB3LG6iIsW/SDA8qq4IiIAIiIAIiIAIiEAyEJDCIhmuotogAiIgAolFINSSgvfQyZbcak+EL05hgTLDfUdZwXfnKiqxWqzaioAIZPMJnC33Xbo30pXA8TlOOKFA4WIlDvz999/rVq9Ymq4nP/qTuecFJYNzDRWv0u+v4LuU43i3Sut/9NdFJYiACIiACIiACIiACKQiASksUhGmihIBERABEYibAIISrCoQwpxqiVWjbLitONvSbkusJkWo4nx186nYFnGj1gEiIAKpQWBvs0OlHBL05hipWDupwTY9yihW6qJyxx533HEb1qxcvvevP3n/JNrmAmj/Eax4XEo/XEMFrSxYBCBr0ES7+qqvCIiACIiACIiACGQBAlJYZIGLrCaKgAiIQCYlgJAF1xQI/VBWnGnpFEu/WvrGEi4rTg/uowm7LCGgIRE4lC0uQU0m5aBqiYAIJB4B+i2swOiDjjElBsJfp0w9ojWm0NCWSQiUKluhMlVZs3zJZ5mkSvFWg3sOpX7ouzCuMoKuoTgmYNVoCoz9wRgXcZWjzCIgAiIgAiIgAiIgAiKQFgTi8nuaFhVQmSIgAiIgAlmWgBP4nWYEzrPEJwqLcy0h+EOZgbsoFBf/s0SQURJ/8+ncRWVZgPE23OKAuCDmhz7jLUP5RUAEDhFAYUF/hMKV/gsLMbnXyeQ3SKmyFatQxQSMX+HIoqzAJRTvyBTHn0BpYcdL6Z/J71dVTwREQAREQAREQASyIgEpLLLiVVebRUAERCBjCTgBCYI9BHwI+hC6IPQrbCmvJRQXbAgDEQpeaKm0JdxEnWEJBUZgX1AIn7EtygRnNw5EJiehjHDf/2PfYRRIVk0sK3GxxSeJ3zUWyATXL6tWwVZ2H2MpUZvPs3O+pUKW8gU/6ce0ZWICZSpWqUb1Vi1bvDATV9OzakErCOcSMTXcWaG0QAGiTQREQAREQAREQAREQAQyDQEJKTLNpVBFREAERCBLEXCBtwn+6VxC4f6JhDsofkeg7iwvgJPfEkoLfsPyAsF7ln+POSVFkIULWo5yAj5YopwQ/Ay1SGH/ScE8x1kZpFBFh1N4ZKmbUo1NXwIoK9L3jKl6Nqd4RenKM5YrmFBg8Hxpy4QEzs+VO+855+W84Mcfvv9u25aN6zNhFWOpknMJddSxnEIUILGcV3lEQAREQAREQAREQAREIF0IKIZFumDWSURABERABMIIIKhkZScuLYhHcYElBH24gkKQ7txFkYdVpCgy+P1HS8S4QFBzjqVvLTmXGEnt2gLFhMfmFD/schlQTCBA5W+sUP4bZM3fsMbvOQJV8rCP3/cErwUrbbXa1ou0fkt1AkngM5/+6jdLP1viueNZOivYL7l+Kqn7pVS/KdK4wLIVL67OKZZ99snHaXyqNCs+GDQ7Nftp3aNpdrVUsAiIgAiIgAiIgAiIQEoISGGREmo6RgREQARE4GgJoIhA2I6Qj+9bLeUMCvtQRKCgwDUUvsYRCKLMID+Bt3EbxeaE7AgN9wcF+kcIXo45JpEXcUfE7BrmrCkQYMECRQTs4MqGyy0UPSgrnIstWLMyHP6/W+JYynPBzFNTGBaxEdopAglMAGUp1mBYV+QLeaZQwH5gib6LZ0kC4UxykctVrnYJVVm6cP7cTFKlo6kG99ZRWxkmgeLwaBjqWBEQAREQAREQAREQgUxI4KgHuZmwTaqSCIiACIhAYhDAXZELUotgb7WlX4ICGNw+4QKK/QUsIXRH6OfcHO2w7whrULw7YXtitProa+kUPbDAQgIlBHE9iPOBogJ/+jALTSg14HemJYSp5OU4rC2IB4JCiPggWLGQN2m1PEePXyWIwGEE6LPohxhT5wk+k5Xt87Lg84YCUc9TJrlpylWqWoOqLFkwf04mqVKKqhGiZHCK6RSVo4NEQAREQAREQAREQAREIDMSkIVFZrwqqpMIiIAIJD8BJ3QPBH62hNCcT9ypsGr53KCQD2UEAj8sK36yhFXFNktFgnmxCPjeEpYFHOfcQyUrQbg54Si8CE7ObygscltC8QOnLy2hfMBahSDAKID4DqevLKGo4DtKDHcN+A5r3HTJNVSy3kFqV2oToA/aYAm3UDxzPEM8m5dbQpj8fvAZlZVFapNPQXkL582e+cGMqZO3bFy3JgWHZ6pDZBmRqS6HKiMCIiACIiACIiACIpCKBLTiKxVhqigREAEREAF/AmExGHj/INhjI4A2LorYSlhCuL7SEsqLspawxMDtCm6iEKajtMAagN8+sbTUEm6N8BnPb4e5M0p0l1BBbk7Bw6cL8gsLOKCsQPkAR5ghJF1lCaFpXUsod1BSoBTic5ml3UFWKDEQsn4X5Mo1gSPCV2KH/JPo/KwN2kQgVQnsbXZEcTw3KAzrBZ9DLJawfkKZisKCPsrFtDjs4BwjU7VqKkwEREAEREAEREAEREAEREAEEp6AXEIl/CVUA0RABEQgYQk4iwgnbGfV/0JLP1j6xhLC9S2WyOcsCxDQI6hfZGmdJdwa4YYFoTsCQqwFkk0Zz7sa90+ujShwUD6goEA5g7ssFDZYV7APBuxjRTfKDJJTeOBrnxXhMMU6g3IJXI4wlePgybGUw3mTjaU1SZsIpDoB+iT6sZ2WNgafSxSHBS2hMOQZ5FnTJgIiIAIiIAIiIAIiIAIiIAIiEIWAXELpFhEBERABEcgIAgjTEejxHsJiAGE8wj02Yi+gmGDVMiuVEbBvt4RlBRYBi4PHEIcBpQYCdgT4KDwQtCPETzjXUB4WKKFus2gXjGCAcgLFAn/TduJSIAytFvyOsodjsaKAD5YSuIiCCdyxZilpCcEqsUDYnJspyudYrDP4jWskVzZBSPoQAQhgFRFmZcEzwrPG84JSEHdDpSxhueRi7zgF4GHPkytHlha6t0RABERABERABERABERABETgIAEpLHQniIAIiIAIZBQBBHcoF3DjhJCdFf+4hCIoNMJ4Yi+gsFhvCTdRuIRCQF/LEiuWsQpgZTOCQATsPwb/RsFBuYkoaA+1aHBWkC6oOG3EigRlDlYV8IEViggCbVew5FzToPRx1hPsJx/KHqxR8Lf/uSWCnBMcGEUPcS9QfJAXhQj1gON+U6Tw/V+5hjIK2kQgSCBMwfCvKR6wsMCVGn0VfdFbweeI55Z9/M6zhpuoROybdO1FQAREQAREQAREQARE4P/YexM4ydKqzPu9N7bca++q7uruym7oDZBNERCUBlwQRQV1QB0RFdFx1Bln9HPcPvUTFcUZHedTxx0cdBhUVHQYka0BEcFGFpGtG7q6i+6u7uqq6sqs3CLuMs//5j3VUVERmZGZkZmRWeet36mIjLhx7/s+73Ijnuc95zgCjsCWIOCCxZbA7BdxBBwBR8AR6IIAu5EpiA4UBIm7ZdMyCHXIeTwnINE/JHt+eSwJuCHReR/PAwsFxXGQgxD92EW5LHZQD1B37s+0rRALZIg5tJM4+cdKrBAWEC8gQWk7QgRYIkrwN6IOCco5zkQLS9LN+TmOc0Gy4mmBpwvXJrQUYgXXn5NQ4eTqDho8XtVtRYC5RlgoBMQbZcwz5iXzjPlEebcMrycvjoAj4Ag4Ao6AI+AIOAKOgCPgCDgCXRBwwcKHhSPgCDgCjsB2IwDJTh4FCHPIcUh2kkfjAQBBD8lOIbcF75No+2nle+SyIMQRYge7mI3sh3A3sn+729fv9U1oQZjAUwIvEzwpIDcRbvCoINwMXifs4Mbb5ItlCDNgc50Mb5RpGQLF7TJw4HMIQHhR4JVCqCiwebKM7wGIROfK84IvhCufpx4VeVgUYaHcw0IoeNlUBF75OqK9FYW5QNgzC+1mIeR6imc/8a+fsql16/PkNheZU4+Rfb6M9cvyyxByjbw8n2VO9XlOP8wRcAQcAUfAEXAEHAFHwBFwBByBywoBFywuq+72xjoCjoAjsH0I9CC8s5IQx0sAg3SHrCecEWGN2JUMQf/V5WuQ518jg8iHUGfnMiGlbpaRp+HDMoQPXhuqPBYdOSqsIywElOWM4L6MUEH7IWwRKyBv8YZArODRPE/4G3zeLgMXdnQj9FDAEPL02eXxfI6wUHhTIOzgfUGIGoQiBCPLj8F1+RzGcdTHcl+Up/YHR2BzEEB0kGhhuR7My4h5wDxhPFpyaxujm1ORjZ2VeiIcMjdtDjPXmJMIjaxxrFXmWbaxq/mnhxaB/G0hir7Uhamt6KA2sbM9rOIFUXBIBM2tgMKv4Qg4Ao6AI+AIOAKOwK5AwAWLXdGN3ghHwBFwBHY0ApbYmd3HCA0IDhDvEH6QfHgJmEcBf1voIsh8PDDwHOB1CHvzIOBcw57Hol2soP5GzIIH+SQQZSA2nyizMFAIM7xOQXy4T2ZhoCB6PyJ7v+wJMgQf8KSQEPiDJU78DXa28xuhiOech+N5pA487tSwWmWz/WGnISBiMRP5aDlUmBeQjvzNvEdQY1wiojE2bawOk7cCdcGjglwVrFuIg5aHhnnM3MIzDGHjQr1Fbq9UbK3o2U4R4162GQH1oeVToib8xor1Gv1s/cdzxGnGMX1pgrCNBbsXXtIS79+LIWkTKHjD8OURA2PLkcXfPXHd5iHjl3cEHAFHwBFwBBwBR8AR6IGACxY+NBwBR8ARcAS2GwGIBQhIxAYIeDwBECzwJID0g5Tk9cMySHdI/OeWhAREPCGhCCNF4m7OYSR7+07L7W5j5/Wpm5FbCBWEtIKc5XXa+WgZogU5KiA5IWvZpc0jx+NJ8rcyiC6O5fOEhQIP8CKZNoVzcR0IMjACO4Qg271OKCieE17qjvIz4M7rfG6YiOCyev6w2xGQaJGLkLQE8JYEnnHKODZy10Ko2RgdprFKHQkL9R4ZodcQUxFXCcdmc89yz3TrTghX5jlEK8bfFBNhh8p7bLePR9q3gqDEms24pJ9YO/EIpJ/pv8fJyA+EuMz7COm3yLi/PSjDS457G59HLP50eRzjx3I8XQ7wbqSNJlLY/Yq5Qj+wHoAjpan1pMCTtWUjF/PPOgKOgCPgCDgCjoAj4AhsDQIuWGwNzn4VR8ARcAQcgd4IGLEAMQm5Q3gicjZMyyBxIH94DtkDAX9F+cgZISHwFkCo+LgMEsjCx/D+sOaxoF7cgxEg8JigvRa3nzYhPtBWiBcTHSBAIbaul7Fz+7jMQj29Q88RIm6SIWAgfrxVBsHJuSFxwBeceA+Rh3PwPueEUANfrk09KEaWOsFTAjLMD0svv7DLmP6yPjTvhM6/ix3Hjd8dHkGqY8c0UHeOO+rMeGUsm4fFsO6cNi8L1iSeMy+ZX+TloZB75n2Vx4UHZNZO1gNIbuY8AiLeVDwiHmKsFR+VcRx/W0gpn5/bMzFNcKa/CPOFwIxwTO4S1lNyBz1D9i8yiHNyCuEN+CUy7mH033NkeONw3+I+9hdl3xJSjHsA491D8vXu33axwgRM5pCFRLRPXvAURLhw0WJ7Joxf1RFwBBwBR8ARcAQcgbUg4ILFWtDyYx0BR8ARcAQ2EwGIGcgGiHXIGkiHT8kgd9ihTGgV3sPwFLCQRtRpWvZAeQyiBySQlWEKa9QesgKhADEBUpLXERwQZyC6Pq98nR235Jl4vAwPEvJVIDYgWtxaYsA52LVL1mGILwhdI2zwqqD9eGpwXkhPnnMOjoNMw7MCjDGwg1yzEDYk23ZCVIBsd5Eg0VkYM/Qzxtxh/DA36D/62cKnQerTt4wtiFTmDcelOie7/C1kzYqeChI3NrX0iDF/oU4iGi3EC/VoH5NDMT7Bp6OPqBeCK15PrGN4SL1Ltk+z/YmSCe+PDhUCooku0219Y/OUttJX9BlrAOsg85i1AC8r1jzEC+ar78jf1BFanLzdM451m7WUPkGAYj1lLf4iGQKVleeXT5ijvX53IVBw73uvjFB+eF78Q/k5+phx4l41F/ev9YVtSjBPJHCkIACZAG95cXj0UIcX4+h/OQKOgCPgCDgCjoAjMJQIuGAxlN3ilXIEHAFH4PJBoEzGrZzUucWkh6CHwGFHMmQdIaIgHiBW+Ztdy5AUkEO8DvGPVwbkESQhBKHFsE50Xl1iKEh3i61N53L/ZWcuRCQkCrtzEREwwoggQJC747jsczIIMEQKduhaIm7CZUGa0WZIMgSdO2V/LfsqGTt5P18GgcM5psv3wRZvDXYCgyl1gAyjfhZKg3Oah4WeetkqBEjUy7Xak/XiPaGd+FH6MQ2WK8JYvqB+aoWpfKkYKwf0ids1ig6rx/ZrNEBwPk2PjCFyJTBOCFMDsY1gwesIYXjuIPwxnyznC2MLkn3oPBfKXdFDIU70ORZMsMCT6UPqoy+XPUMzf09UV5+NhidEI8UcZ91CYIWoJjwQ/cQayK591rUnyW6Q4XFB3+Kl8RIZ5PYbZJ+R1TRueK9nIm/PgbByr/WRQ4R7CkISay7r9GNliEjMFdZS5hh91aus9JsL0YPz06+2Fn+5nuOx8RbZn6h+zE3mKe9fIk5dpv1rnormXcGjCbgIe8wvRFnua3xP4O9kGL0suow/29xgHnN2T+46vi7T/l95Uvu7joAj4Ag4Ao6AI7CjEXDBYkd3n1feEXAEHIFdh4AJE+woRZwg1jdCBqFQIHUg2C2OPeSchYOCfGUHM54ZkBbc34Yi6bYEEzrJ8mlYLHojhCFXCAnFDnjCO0GuQCJDrCAkQIxBZNJWBBpS60JiWcgRBAnaCeFpce/xtIDg5LzvlHENdtdDsFGPf5Kx45vzQ+TwHp4VtoPdxQqBsVmlBzHa7nmDpwTJerP8fGil/xKifFYixUOhUbkpTErWe3I0pT6dE3H6sLxsIhHeFYkQsf5uhZfqfUjV5VGRhpeqV/G6IRE7ryNiQXj+vQyCG/IVMYvxBbHO64hezCHEMRMyIokmjIuegsFme2BsVn9s5nnrLwl5S0mX1X/VKFYvVcLRaDIck41GV4VbovGiP1jPmI8vkyHOWv4LQrt1K19bvsjct7WC/BiIHHhdsCZ6GRwCzAXWSQycWWcRCr9RZt4TG72a3RcYD52Ftfy4jPvf38jwmuM+MXSi4kZBWMfnLSxXVK3Gda1OcZJm43Fc3G7zLMsR/FhP6TsTYrkfLki0SLcyNNQq6367t0iRrL001mfzgEOAQXzmuwHrNf0/rCEv19GV/hFHwBFwBBwBR8ARcAQuRsAFCx8RjoAj4Ag4AsOCAGQoZCpkDLuMIVoRLSAabOcwP9oJl0HybTwHuI8R0ojX+DzEBOQ/n+FHv8W6386d2UaqgDP1gzjmNcgvBBnqiNDCDl3aAvFI0mzL14GgQCgZ88RAaODYZ8ogMP5K9iwZggSeGJwTAQNCg+sdK59DboCT7eAFI4QhrsfxlvvDw8sIjEGXHoRV+9gAf3bbR+q5fRrN0xIsTsRHw6H8jMZKLRySUBGipfCYaF84k90d9uWL4esjKK1Y3jOLIubGwlhEr2uE5IwMUV15S/MhCy8o2rNMcUKQk7QeYpvxYQVxgjj7fypj3iFoIGYgXECSMV6Ym8MUYm3Q3TSQ80moMIGyVn1GGM1PhpP5ufDuaG94ofrrqeqpLBqVN0ylIFMJy/Z1MvtOTv/0Eis66/dqvUBP/6yMec9oQHSiv4ZCsB0IoNtzEvOIY44ghkN0sy7jyfbdMgTmzSzypyqEEQTrP5exbuOJ99vlc+6RrNuX9Xys1yrx6EgtzfIwmiV5I66kFXlUTkbaKNBMsvmQ50Xy+izXSrg8x+hX81LZju8FJk7b+OJezjrAfd3u3XwfoK5PLseZhRP7iP5m8wYbFqww12nbdrRlM8e/n9sRcAQcAUfAEXAELnME7AfVZQ6DN98RcAQcAUdguxFo80Tg3mRhniDt+dFuYaH44Q4p91kZwgTeBvyAh9TnPchVCDx+7LNrlb8XRWBsOqlT1r8TRiMlLKEuggGeDxDVhBOhQE5AgvEe4gFeFRTLPcDua3bWQrw8UcZOW4htSGXCPyE68PrzZBAefycDH/JggBG7TBE8EH0gNj4pM4y5HiG0OFdXcacM2VVWyR/Wi0CHYGHfvxCvCP2DGFAV5fQFoh9Py/CaeGGehLrCB92Yz8nToRLG9fxKvdZQKCHmx0Ul10hXqKig3fxBx4VcvR1p1En0CBI8itnAexI5lkdW7xmBKAExBoHGuGPsMqfeISOUGJ9E3IAou7DL2z0slrtD/cy6AwGJTctu0axjDj5Bs+55QhMCetAFsvI9MkJK8fh6meW2KK7lIWNWhrycn0Ym03eI46zLCMHMBcqtMhJls1avpzB3/ouM+9oTSut2HtZ07guEAews36IXuO+xZiNOWd6hFT2gdlv/y0MiklDRaNSr4+ON6llIZEIAACAASURBVGgrSQ+GOB5P07TebKYHtDBNtlrJ6SwLFQEzrvvzGakWCLBshGCNQ7BNtsrLogz1ZyGr6H88JhHBvkzG69yLnyb7x/L5i/XIdwXES+79hIKj/qzJ3MsJ7ccGB0I88j0HEYM1uatwsdv6/5JZ4S84Ao6AI+AIOAKOwK5DwD0sdl2XeoMcAUfAEdjRCNiPbdsdDCEKxQpBCoEDec8PfLwTeA0CFXIH8gHilx2okE38eOd1fthv185DC/MA2YDIApGJ0SbaQuF1wrggLFiyUNrFrl5i03Mc9ec9vCcQOTgvRBqEJG1GvIDsgLwAB84FifFWGUIPZOn7ZJyX5+zKhdjgPGBku7F9R7bA2MRi4pVdgu9ghHthPJ9SLy/IvlbU1bhIbV6rIjhQJFC0JFEUIoW91llPeV0ErFvJjutVUWKZqLoIAUOzQiJIr9mBiPL08jzs8Lbyh3rCOIMcgzxDFCP5s3nzbNc828Qu6//UIiQtFB3zkXmKMb+b6s8JzbZ/e+FsuXq6JdK0XszHQRTGloUTQqhEhETIRcDYzjVwEG3bqnOAIQQy9xAECvqRdZhHcCSnBOI5a7GFJuxWN2bW28tjOCeiA68xT1jr3yiDbEZGfLMMAZrrIYJwf2COmTdHt/P/Ufki5yKvyf+WkYcGwZnrbLo4361SW/3ajdMHo9m5pahaqexVBKipOI73JVl+XZ6FsWo1HJDLxVRUq96tEFFnoihMVuL4wWYrS5M0bUi4sPvfloRUKkVM+pbNCM+QsVJz/6bg/UafcX9HJPvWHljaRobvbHsfIfknZXjjIG4wTvnewPcAv59v9aD06zkCjoAj4Ag4Ao7AQBFwD4uBwukncwQcAUfAEVgvAh0eCu1kPz/iCckBIQjpDknDj3dyMUDiQtBD8JiIAckPWUes7+JHu7wELklSut569vpcl/pDUJhnBSSYxaYmlAhEL69BgLGjElKMxK1vK9uCtwShYtg9CxEFifX1smkZcevZdUn7+BziBaQVxIeRVuDEZyDFIEURMxB32FkKPuBGfSDesJ4hMtzDQuhsoJQ7axkLjF8IbMgqyCXGNP2I6DQqCvvxIrVNKLj4ihYQZAP1sI9mUFqi63JJegorFeSxsR5qC88eS/hMzgvz0GGeJfK22HXixSox6JlLkNusTQgVXyQzgpE5ulIy5tV6FaGI9Q3xkXWRc69WWBt+VYa3FWT2UnsS99U+fDm93zY/uc8gHrA+H5fx962yl8vYEb9aYX1lLUZIwKMNLyXEDfqO/mDdNa8XjmMtQFhnPYBg5nrmbYcXx/fJ8JhbrfwHHUA/cyzec+zCZ02/qOymHfYfOjETnZtdrD54Zq6h+9ONWZrub6XhQKUarlucTw4sJa2xLI/G9N6MPC6Ot1rpWIiie/Msf1hhohIlt3hQggb9hfja2gwvi1LAtPwnlqfqm8p+5978BbJby79X6+N+30cA47sA3ykYc4wvVnj3sOoXQT/OEXAEHAFHwBFwBIYGAfewGJqu8Io4Ao6AI+AIdCBggWsg1yEDIesgYyDyCYkBEcQju1Mh8fmBzm5WSCEIGwggvDMWJCaIu4i2ikS1nfSQVUUCZRmiAQQ1f/M6cashsdnN/mzqWLYDAYPPQ3DQFvJPQELRFks2jkADGUrbaR84sGOX80FOgBHHIk6wA5MQGBAz7PDlePOo4Bijq7MtxEeXvTxKSVrRP4wBxh8CBY8Q28/Vs6vV29fp8b6eYgVQDfDbWmw0OqIFvU8wNc203LJT9DdLvlqfwiBnIcYhyGhnMUeVoLsgAnejcNE2ci3JPXOTucgcZ/c0yZjp537I5s6JwM581rr3yhArmaNvkYEn6wa9hQDyHbKf6Pxw29+IYP9V9mdl/3xEY3FOpPWmC7cr1Gmo3moL0WNrM6GfMNZkZgEJtV/WZ6V/RseRV4lcQjy+W8aabnmZbMe7hZyCsGZNoNjmMbufUZ8Pyf67DIJ7tRBihJhiHv6ajDF3mwwPm13Z14gVpx+ebywtJXV5TeypVqOjrZBfH1XCASXbvj6pZnuzqCJfijxVOKj9lVq1vtRK86Bk3EprQT7uu7XssaLyPcGE1v5WvT4HQ7nuI0pxn2etZwMC6wXPuVezZmxGYcxiePG8ScY4ZB25LLxuNgNQP6cj4Ag4Ao6AI+AIbB8CA/wJvH2N8Cs7Ao6AI7AbEOjI4UCTjMhoj019yQ/rXboDnnZa+6FSCQXFDmPIepIBQ8KzM9VyNEDoHZdBAiFWQMrzPjsMzYtgoKREjzFnhBRvQzBCUkBOQDJSV8QVDM8HjuU+DJnFcwgmBArbhYu4QNgd2oD3BQQIO305JwQEXhOIN3iWfED2aRmCCAIHr0GKIV5AyhTxumUUMLqwr96FihKVAT5AhrbtaKdfMXbU/kLZLwhSX3ZhhD+yG3/lWrQHotmo14VGSvUpqtgD4WR2h8ZETeNTI67IcdGb3mLMEcbKCrlTXiNDMPx1GWP9/TIIVHaLM3d3W2GuIiTQp8wl5iTGvEW4IA796mUpnJVI9C9aAT6nkF/gTxg3duVTeE64NtaHIg9PeT3WMHAlRwXH4qWFcNErpwJeWQi5iCD0C+e87EspViAQsKbiUYHAxPxkbQXLHy6xXwkrZuAvl/0DOYzHxOtkrLuMhSKfQIdnS/s96KJZpjoRugtRmf7lHLzP+o1HzTfIEFIox2XTHRVjHv6+DILarl2Ihis1YCe+d/+p2TiKo1qa5xOKrKb7pQSLJHuiwkEdjEM2udBMR5qtdF7eFFlciUI9rtwwWq/l8qq4r5Vm5xUOqpqmOdl9kG6LcJLkwxiUl0UZ/onvKnjL8cj4Yk1gvDC2rB83E/4X0S4ZwhXjaEH1Krwt3NNqM2H3czsCjoAj4Ag4Ao7AIBFwwWKQaPq5HAFHwBHYGAIWBsnWZh6NWLbd80Z47Mrdkx3w0VZ+bJvgwNsQ8bwGqQPhBPEPKQAxyvEQ9ggDEIm8B362k3VjvdP/py0uNqQmBC7kNHWlHeyehbDgPUheSxIOoUh9Cd8yXX4OUYbQURzP59gpiUBhCZfZyYsHBcKIhX5iRyd/gwfEFTuyaT+YXRT2aSvCZPUP2e44si28TFXPmb+QYpDK7Lwmt8Azu7Y0KsbHRYWQTSnBljRq8IrIRa3l6tH4aLgrOqAx0Ar3RlMio2OR5LmIt1xxzCsF8QoxdY9e/wo9kgtjxRIfDkdk5LR4R3ZPOKHrfrIIG9UKP6D/GU/tBfGLGOmdu76Zl6+SIWggVhSeT/K0oAXNXeJpYeszj+DCekPc+S+VkSAXsXH1koYT6afCm5UA/c5oMixG42F/Pho+Ge8R2dwoCGvO2553IoNkbAtJRbg3+sDCxYH5a2W9RIsf0nsQpq/QOfgs4WEuh/vHSn3BGjot497B/ARLnn+7jLBQq5XbdcArZayvEMPMC9Zc5l4hDq+TGKbv+TxCBaIF9312y/+iDHGF+fzSFSqHFx/tYvxw77C8Rlsh1q+G2Ybfl7AQP3j6fG1ivEEIvUlt8ri22crHladiZHEpHYti9UEe4Ts2qQbX41Cpy8tipF6LlrI0xr3i5GKSjVQqWTPNivsh90rur4gWPXM+SMzoq+6lWIF4yQcI68W6yHXYcNBvQYjkfv6FMsYVY5PvCYxT7v/kq/gxGRsfECN7eeC8RO+xTrGRgfP9gYwNELtiLPQLph/nCDgCjoAj4Ag4AjsXAdu9unNb4DV3BBwBR2CHI1B6VkAqW5x7nlvsYwvfU/yoltmuTF4vym7ZId+RA+JC8/QEMh88+MEOGcDfhL4AD0gddkkiVLCbkB/okAT8QEcQKAg6lUXhtKlhEdo8ZKgr91cIJupJX0HgIlhAYENy4v1BHSEk6FtIDYyd1ISM4HO0jb8hwvgbMpNkx/yNgIEQAhaIFrSVY7ku5AZjievaLm0bR7tmvKht21JWyWUA/ohUjEH6kbBe5BZht203on+5Dan+VfRPIySlh5EvNLoJ01SEaorCQjwd/iyaEHm1KLFuJGRRQzvzpzRGKsU4a2iGQE4y3hlbXJ8xQ30IM2ZhwyDBepdcu/7nwqslXHwg/Zh2jOdqQ17MLfIyQHpDpvE3ZNxKBUHxz2X/ILtNVmbO6E2WSdTY1tKjX61O4MhcA1vmFoQ3OHyd7Of6rnga3i/h6cOyj+ZnwpweW5K1FuVh8cH4pnBS/dvqJSZ0qZ+tM6yJ1AMym8de5S/0xg/KWCcevBxFizJUD31JThE8KliXWUfxgPua8rEbfqy9rNPkisC7hXsNcwEsea/wpuCD6xQqwgrjD1Id497xVBnrCnXvJUZyn2PdJ8fM/5ThWbO403NY4AWhdsT7pkamJidHDk80anuzPL9psZncuLCQPEkOFfsrlUraStJDWZZNKQrkQiVWIKiQ1yRinJe3xUmFhJpV1u37l1rZ21ut5HPKYwFOiEynJEpsyBulFKvxsnmcjLUSEZP+Wq0gfrH5gPsGoeBoJ2PrS2SEkLpbdlzGBga+E7DOI66x7rMeMa9XK3io/qbst2TNy3HurwaQv+8IOAKOgCPgCDgCw4eAe1gMX594jRwBR+DyQ8DEYxMqLJY1JAWECD+qIcgw/oYog+hmF2Wrg+jfsSGjeoS2UvNyyCAwgYyl3U+QQcqzexvM2C3M3/yIBzN2FHI8BOPaIvMPZuzRn5Ca9BVeDvQT9YHwgtCg/yC5qCv1Rnhh9z2kGSIGAgTH05e0jePZGQlhAbnCedlNDWHB+cEAbHid8y1T3MvhZCCvCtstwpbaMmzFsIb4ZNcr4gR9RigQ+skSaTM+l0saPidh4IQEh6dnD4bZ7JNhUl4TIVcvYkVOCZPaUvVxHL5HMdr/Pj8dxvX6fHx1OJ03RW7Xir61dYNxRkG8wlOHekFosQsXgYuQMez0hbjqXqKwT6T5z1duDN+lUfsX2YnwzwoRlegqiGkQpCaIrCZYIJZ8l+yrZORR+F8yI3gtNFnPagzRG8wh5iKPiDZgQP2ZY7QNz5nOAqnITncKQg3rETuj5/NWmM0XwnF5WFyjWX9Afz+oWc46wIhpVf/9mjwfzEuCEHl/ImNN4TrfL+sWIx8xA4+A22RvEsHK8esm2Lu0e8WXlHug/f3inveka6a2bLd3m/cT8xJPCohliP/VQvS8Q8cgSuFBw/3nb2TckyzUG4+EftqswrxmzDGPGVt/L/ttGVckbwX3ufbCvYd5Txs/KuOe8dldkMOkECwWl5KRKCwdai2lByRCKE9FfrCVZ1NxnjclWow3k7SeJFmoVSr6bhTmdd8bjyL9GccNfZdYzONoQo+3xHohy9MTOoY+rUoQAeOu47HTw6KLuETdWPNZ95jPYN6PFxNCxavpHxniBJ+z3FLv0XPmM33OdwLmK4awwprCmo4nx/tkjGPzvLxoMJR/sEmC8UCOnE9RfxctusHkrzkCjoAj4Ag4Ao7AMCHggsUw9YbXxRFwBHY1Ait4EBjBDdkJ+QDhwM5PyEGMH6L8EIYQhbzgNT4DuW2eGWB3UcifXQQmP/z5kU6bLQwU5D47Ti3iPseAERhavHdwAx/+3qpiYWMgLRAnrH/oM4QJ6tme7Jp8E5Cb7IiHOGFHOmQYRIT1O8QEpAWJWDkvYwTikV2+7NqnmCeGhcbiNRsP7lUxoN7vQVTRxxDEEE6Mz+tkCAaQX5CciEgQiBfCPmWnQqbwTlcrGwt0Wa3wpBAVVUhzJlNl4Y/0HCKacf3e5B/DqWhP8bm09pOXZploq1shZJZN5jljBTKN73zkRmCcQXheEobqAkzV8EuVJ4YbK48Lr9Ee5HPZXWEhvSv8rUYUdWFcPVf2r2TfXY69XudijkKg8zmIOYg3vC8u7Ei/cM3hemIEJF5dny9j/jL3CL9CIuSViokVMPTfW7ad9r8jPxuS9ONhTI+Mkbr6l9A/zPOFNYoV7ddHtKKPRUMW+LIG9PL6+E69R1JwPH/+UHafxg1eHVsmHJQV53oD9/JewUuBeyrCBLgTKg0PCxMSe/Ulu93fJfvfMghl1moL/cQcoP4Dw20VwSNT2+w+SB0sVNRtev7lsq8tH9vbwnj9NhmJxBFd3qVznNV1NtXTsBeYA3gdvMeVP3tP1EwOV6rxvpFqZVwhnhpJM6krP4U8KQgTFY1JxeD5uHJdSKjXelmp1JXXYkoLdaRcF6l67spqFJ3Sm2f0vYy1iznIWlmIT73qusL4Mg8s1gkExJetMr4QHvCs4H6PqMl9/Hh5Xb4nsH5TD/rZhGjepn5ci0fWUDZt/JKMHCZ8B+B7A/kruhU2euBtx/eGRbUFr5uBjd8e1/SXHQFHwBFwBBwBR8ARWDcCLlisGzr/oCPgCDgCA0HAdmezHkMqmlcFP0YtFITtzObHMD9g+ZEJQcr7kBf84OYRo6z4o3sgtd7ak9De9l3ZeBVYXghwgjAGP2J22w98diqCD5/Fu6Cf3Y6DaJXRzRAOEIeQCEbOWV4N+onQVdSZPqXekJvsjGcMQHLTp/Q79aa9PPIa7YZEhaCEyIB8gvywpNp2LasHYsUg2nXZn6NHSB6ILohQPGQgDek/+op+5/XHqfffJzukUfpkiRIPZZ8Ji9lJCWvVgnBa1P/3SbB4VDFKlukjdnArFnuxc5Zd1YgMDyhkUjtxdUl/dBCeRkRZ/heSrloIoT/VhyG2iYXPGIXE7iwILD+sOn5ptD/8WmV/uC2+IdyX3h5OySOE80DK0Va8JiDN8DwgUXGvAknMOCY8zcdkhChh7A8jYUb7ED4RW+gjvGQg+BGRVxMraD87ozkHHlG0j/nJTuo7FGZrRKGgnqlXmZQQhxhi5aqlD0KbPnl3iS/rCeGfqHdn4d7xkzIEUPpkVmMj3QbyMpfXBTiYt8WG1ugeZDL9wBxlvaU/ESroT8jblQp5WJZzwSzfVzkHc4b5ZPXcrrHLmm/3BeqGxwWiWrdCCDiMsGEfoP7CaWYb+noVuPt7u1qNI4V5qlWrlYpEiKk0DweVXPuIptNkrlwVCvFUrVajtF6tJOr4WO839NpCnqVRHIfRmvwsdD+cregvhY26IloWDBkjlI0k3ua7xg3l+OC+/bIVWvQTXEvGOs+mk2IOykxIah9X3cJU2Z2Ctfu4jDYgfrA+ES4K8aLbvKdKr5X9jgzPnHtKr5udKmD1N2j8KEfAEXAEHAFHwBHYsQi4YLFju84r7gg4ArsMAX6Esibz45md+eyih/CEeIKEN28CSBTINCOmIa75sctr/PCEuLYdeBsigIYF35JwV7jq3DwGwOS4DAK/XRSA0DVyCQzMoyHSZ3Ua0RObXwqBpOwz8IdEQGCgUFcSglvibQhfI84giOlD+rcMClQQ1JARGDswIc0YCxAciBycn+MhNdoFna1o5+YjOdxXYJ5a2Cd2apNMm1309Av9O6IZCtl5Xo9PUOifUxqZH5dg0cjuD5HCOu0vqfoP6fGqNtr+H/WZ/1H2OeMAbwQ8NFYUK/qBqi0ECOLFO/UZ5hFEG/X80aLOlxYI3p+V/brCV/1p9TnFbuCF5uuLOhFehHHLPKPenOvf9agL4cu+pzTi6v9XmXkJ8flhKObBRZtIvEwIKObsV8u+so8Kkt+AnfiIBsx51gFwYv4iTCQK6QVGth6wVrHWm6jZxyVWPIT1gPoyVv5IRjgZRKRudedeQ5iul8nImkLIoPZE35dcaC0hj0ohot+QT+Be02fAKxlgmCjOyz0UrxjG8T/JCAPFOOxVEODAjbkBLuyAPy5DuLId+Ct8fMvesvsMF6R+hHn7Kxnhrn5KxnxrL1+vP2gbnhafKD0thvI+odBM3UAsRC2pDYnu40meZfNLrSRO0ny/JIhmvVaZ0T1+XtsSRsYb1YoOzNIkq+dJyj2zWq/F81GImR9nJXgc1zet+5aaEuqi6LTS2dO3G/GWMdGN9Z9E14Rn6iwICdzf/1aGoMncZ93l/l2EolptfvUQ5GgT45J1GUENAeTnZXgSIUSbt1d7fQjVx/cO1urjOu8DO1XA6jZQ/DVHwBFwBBwBR8AR2D0IuGCxe/rSW+IIOAI7EwEjDfhhDWEIIc2PWMhQiE8Ibn6UsoOb5/zQheDixy6P7LiHiODHsu28h2yBuLKYzENJTKyju0yAQaABB/CB8AMz2szOYX6wQ3xB4luc8XVcasMfAXP6lD5BfLKk29SXevM3fQyJBjENwUR9ESb4DG2hDeyCJl41BbITYgKChPZvdxs3DNIOPEFBrsognyBDIQiZh/QdfxOeRSmxw53ymmhoJH5UOQvuUlilRna35vBcuEbixeiFsE/LROoflP3Ozm+EBIhHzkd5xO9igGCJoFoSUQUzyPpheXJu1XO8RNoLXgLU6xdkzDFC5HxG3h58prn08sKLgPlHgSiFjPtj2XJehu4FLwUIszfK3irD44Jzb1tuC2FBG1hfSWjMbnTmJ0T/81ZoR/tbrNm0/W4ZhDciDHMUwem88C7aJrx4RHBkTeAzU1lUOdeqjCavfN07O12hLlq3O+Por1Av87rCMweMaQ+hYDoLdUC0eKWMZLyEnRtUH/RLANv45vhizEi42KhoYThyP8VbDQ8D2o+YtJJYARb0IZ4IiGncbyCB6UsI5WG8j9LXjCc8QhjDloy52/D4//QiY5pQYG/UmD81pG3qVndey+M4SpI003ebKNFgqdWq0bxSUTwgL4s9EjIOViRVNNM0by2muUI/1aIQ1Um8jZdFkrYQPCYUJmqSHBfKfWGhI9vHYK9r93qdsca9mjWS9eNbexz4er1+XMYcw2uOuW/5tfq6Zh8eVtwzEMwJI8icx5uN9bybBx1zAnHlz8t6XJRgpq8K+UGOgCPgCDgCjoAj4AhsMgIuWGwywH56R8ARcARWQYAfvOzWhqxhpxxEKEQ2Pz4h3/kxDCEBCcaPXAhOXsPjAgLGdgVDPvE6QgY/iCG2IcJJyr2bEi5DIkGqQRobqQvEvA55yg9vsDASeas8Kzq7GRLEwkLxHv3LPZe6s+MaEQKCm/5iFyREA8ewM5K603eQG/Q544O20jbaaYJMEfprizxHOtt3uf5NX0BmE2LGQnshJn6RDDGK2OktJdQ+mN0XFvJTSo69oHGQKxzUOYX+ycoEucuJXtl1Dxn6JhnCFeIH83ZLdnKLACM8DMQs44q1hjHI9f9NW+dCwln5dT35PdnP6XOEL2McMs4LklteF4xZdhB/h4z8FoxlsOlWSP6N0VYEvDtF5h8vz9WVGJZIMvBShsliHjIH6UPWDvqGBNWIT6sVBBcEY3ZQU38ECuY3nhVJF0KYuc06xVrQTONadak6efK+qc+zNc2849p30FOHtZDl1ieEiIKQpJ8IyfXiHo35dr3+hvIa1K1n8uHVwOB9C/MkT4l+Pfw4jrUSTFjXCRWVbsDTgnWUeyEiPt4ViFCPlv1Fj/pD9nNt+hAxHPwsF8hOCK9oY4W8OXwvoC+Zf90K3mCQ2czz/1Pi3k+3btkxPYS5XJ4X8qjIlLYilkdFvCgVYlF5LOaUu2JKXhKL8rJYaKVppNBQsSI+RZUoj2txNM/TLAuTWriVgDtIu8gPSay4Q9bUZAO79XrPMGbYXEDeCMj/b+kBEusiQhjCLOvCZubvoT0WIpLrkFcJT6Fu6/DL9XqRE03r4EdMVN2yjvYLOQKOgCPgCDgCjoAjsAoCLlj4EHEEHAFHYPsRMHIbogyCENKB3XcIDzwnJjE/dDkOUhECCsKBHbTEP2d3Ps9Z0w+VxuctcSPhlHZT4mUjSi0EFu0GGwuPwCPW7y7fzRgBXB8yGrHJdjxDdNMvEJrs/qXO9DfELiQhZLjFpbYkoJAdEA+QEBf6s/ws9V4LkbkZ7byczmnx8CG3EQ75mxAzRup/Tr14rzwojqjHblDPZOr5qyRUXKUjY/21T68hUlj4DpIkQ6wiPCJOWR6aLYspXhLqTRFW5KGAbGeMvk4G4dnNS4LdutSb8Ys3QbH7vBwEjHna8BYZ5C84/YgMIaBXYdc384HExhCtkP+sdf2S3Sucuvdbaq/t6Ad/SG3mIKFcaMsPrHBS8+BCZEHYYY1mXjI/EXEQJBAqetW/mON5FLeSqF5rVccWPnHFl7c+fvgrEU0Qqvk8x9hawFhYb4g/2gKWiEhgjDhFEvDOwq58vHqIa09cfcbjRknVWKJD3i5a6PkKsIakDAlFuy3EzlrXNj7HvYCQXuQToK38jRDIjvJuBUGHsWrjFpzo42EJU3ahzqvssM/JR1D2NeMQI5TZTV0aTX6DZ8tIwl0keN4pnhbyjEjkJREWFpNqXImq9bzycEMJtdM8PyBraQAou0WssFH5iHJU5EHPFRpqQe9V9V5T3hgn4ig/reX4zsU8vUuHWAi1VdebjpBMjFMGNKHj8Gxho0mvwtxiXLH5YKPzaoXLXHjLvk9yn0Gk+2sZ3yNZt9sLnhjkP+E7ZYM8Nnq8aM6tFqaqn8r4MY6AI+AIOAKOgCPgCKwXARcs1oucf84RcAQcgcEgYLsjIaYhq9gVS+HHIz8yLSfD0/QcwgmSkGP5AYzXhb0PyQQpww9oSAjILx45Dz+upVnk2S7ajd++8xUMLXFmO8G3VsJrMD36iHhCHS3UAgQnu3YhNyA46R/EDEviasmaOZ5+g9iwsF60rTNPBXXdrvYNCqehPQ/kVDtZo7/pH4RBiO1bZQhK7Gj+qIzd26PypDiXnw0TSqr8oISLw9lD4Zn6+wbNQMQISGPmMKLA75fjFdIfYpE5TIHQ2jKxoh18CHbi2us1RIP3yn5O9v/KuiWZJgcF5PYfyNg1XHhYyAPCQqs8JG+JItxR2TaIfWLo9yqEU/lumYVKQnwFlw3t9O91sdKrgu+/7DSH2Iaw/0YZHhUrhbLilHjC0GbGg3l08Uh7Wb8ZN13npTApvOGSuFFPKiP3nhm9dqaRzh3T39NnR6+FJEf0sNwo1I/1gzWgeK4d5iZY9mgaG70vKZyD8UfhpFxEUQAAIABJREFU3JCYhIDqLMf0wnPLNrFGfVLWLeFvj2tf9DLX4RyrksAdJzPRuQjphKdGLy+LLvH8zdOQ+TktQ0hkXEEkI2D0KuCBYEEYKLze2r32+mnrMB1jgiHr0l/KaNt/7lHBf6/X8Sz5Oxlefuvt661sf7EJoNlKpUNED8Rxhe9CR9MsVQCoCE/SVhSHRX3NCRI2tEVD413JLqRUnFMS7kYrSSv6FqSFLp9R1Cj0jAXZhXmrc+HFcUl7unh8MNZY/xFkbRPC1/QAAi8WPBwKjyuusYWAcT0EVeYij8+Q/bTsy8pxgbcc7cATiWPxttgJ42ALIfRLOQKOgCPgCDgCjsB2IuCCxXai79d2BBwBR2AZAfsRy5qMGMGPYH5IIlhYCCAIJbwpILPZEcf7FIg9fnASjuZZ5SPEmcWlhwSDGIUUXSjDQ62VSBrWfgI386IwjwrqutXEQDd8rG4Q0GBPnSwhOqQoO6ohx3jPkqZDTtKvmMXXvhD+aReJTcM6nrrWqyS48aIgDBQkPMIhuUb+RTP3mZIY7lc6+KOie8aVVHksu1c7tNPwPgkYh/UIqcX8pI8RLSAH+SzCBf0NSQ+Z1SoJ/+3EhjFLfSCuWHsIwvQlMgj9zoIXAsT0q2WsQRcRcWoL4/2MSHpCoUDGs8uXcDSv6DgR49ySfSMYQB4jDLHzF1HWBL2B4FLmqkA8ZN1AsKA+ENsreYFwbdqDFwpt5RFPEPrxQoiX1XYjv/rWfwwvf/+LFiVSzM3X9k6dG7nqWBZXD54ZOzYb4jhT6JpiHWAnuMAEzwMiVAlRZSHCqPOKibF7gMQaghBO30JmI5yx+7698N7zZVwXjwTWIIjW9RCYds8qhIc1FhO91vpZjkdEwvOJc7CuPnOFazOHPyWjH2+TcU9dD7ZrbN6WHM59hvwFCFVgQn93I9Rfo9d/QvZ7ZT6LbRFL+0VEwgGCAnVUWKfQlKPFKQkT08uuidGZqBIaSmGhsE/KXBHnR2uVSIm2ozQPeVKr8npo6fjz+vDJVpI3NbdsPhVeD5y/z7rwOUQAjkcEwIvMCnOYucSah/cYghnCCvNoO/AFHuYj6wj1+g0ZIpXNbeY59zbWMYS94l7UJw5+mCPgCDgCjoAj4Ag4ApuKgAsWmwqvn9wRcAQcgUcQ4Id0l4Lng5HbvM1BkHiPlbFb1DwwSI7LD0/Ibn5YQrbwY9hCDLxAz/Gu4EexJW+GvOGHs8WoL37bFzsRo2jHiRa98CsxwoXE8OOxX/JhYEO0S/2KOqheEGFGVvBoooQJF7xP35jQZDkrrA07IY76wHAcwhMhBkJum3gEqTOjEXa9ZmRVuSrukCfFQjQR9mQPhCcqf8XV6k12qHOchbhhJz9kMV42fPdi9zOixbD1re3qt2Ta/0F1JBlxt/J9evHdZVsKL4vOIuGCxNx4JBAKi12+eKQg4kCUUkys4Dmh735Hdlz2m+V1IV0HIlqIlAV3+hLxF5FiWgY5D6G7WvklHQAZCdFHG+hbiOG++k9Ea3TTqbfHH7z6mxp6vCqJ60fOjk/np6Zuzs6OXrM31Eb2KFTNERGsNbGt9yvm/mIchXoUsuMiWMGW+wJCi60Nl6zfqwgmSRkyiDH88zJ2fpOTxAr3F8pXydh5T84LBDXEma59uwJgRuhyyFo/a6ct7omdXhZdPCvaj6cNiGufL+uVw8GOJ/QVY5dQZIgXhEXacffEHn0AduCO4EdIoNtlfA94WZfj8bZhrXqnsMXboCcGqwlyK4yHgb9FLoqWEmdroD2s0FCno0rlXJbkSaUeGpogE3o9arVwKOVLV5SkaXqiWmVeybsiyT6T5RnCMSIe915Kv2ICYxvyn80jzJFv6GgcogDfy5hbrHvmZXlus8fXCv1TeN6of+lnxBPWYYR3y8dkYdTYLGOhJwfeZ35CR8ARcAQcAUfAEXAE1oqACxZrRcyPdwQcAUdg8AiYYMEPS8g5BAbIIsyITXbkE/aJ3doIEZDe7FhmJymvIWLwY5QkkPwghfyGjGOdh4hgpyU/tIsf0CLRtysZ9eDRK89YCgZbLlT02SBwpy/YmUlp97ow7xDbhQmRcIE4cs+KPhHehMNE8jBnEA8J+8Qu7CfIIokVd6uH6hInJtM7NBfPK7FvJXxSEdFP6HXEia+UMWchsAixhHcFgoV5SFmehmEcr9QJ4qpIyCr7cRkhorqVn9KLt8lOC6u8WzgkiRYtiRYINaxDPLIufbMMwaObZwOCBufFm+F9MtZDy+HToxoXv9yF2La5h+cIwi5r5w+ucjJ2I0P80od/VNYDPFiX+xIqOD9ihR6imcbheiOZPfrg5E17qiEZPTN1w9y5iemRpcah6ThGp4hPVSvRfu0IPybtFaFmPsviJWUMPqEwNovaHU5/IHK2tBt8zeQ6fSNcELO5j7D+vEP2nC4Y0N/gzn0EMh/sL4lvvwJ2RXtlFqavrz7rkuOin7lh12KusVOcsdNLrKAdePwgxr1e9kEZ4zzbKTkc+gJy+SDGB98B8AJizcETirBniF6dBUGSfB+IG/R332N7DfUZ5KF4R5yUR9KywJ8roXYUHsziUFOcp0mFhzqnsFFnNHgWJQAe0nedfcp7oQmWz2pe3a+/Tysr90klGDLvqGwN3hXcvxHF8EYiXxj5b9oLQiiF72NPlb1LZnlvBonBms+lMZ5q/rN2IVxwX0O8RbThNUs8bgLOms/vH3AEHAFHwBFwBBwBR2DQCLhgMWhE/XyOgCPgCKwdAQuDYTvt+QFJfgp28fEaPyxtpyrEETtJiTcOSUPsbYghXoN8IaEmuSz4UY2xk5BzQLZaTgRIi2a58x/loh9iaO2t8k8UCJT44kizHL3ikXjR5j3DYSZStL/mCLYhUHrQdGJibkvtj+1Ygv+ayd22i1joNUhOyLya6Lwz2clwXF4VjxPNs0ez7sqcx7zYtcquZsIaQWwxN9llC0kPuQZhb0nUbc4Pax8b4YlY8NZyLfm2sv54m1hBzMH74MdkMxBiPUSLXKIF65ARqITXIkwUJDNiUHsxr4s/1oskhsXb4qP6PMRfz7Wq/pJLoDQymz5kfaR/XiR7sYwcBysVyMzflzFnWYfBgf63ECurfPyit4uY9wu1vbW5+sG9I8n5WlYfrzVrew7ntcZUVhu5rlGvxo1GdY8I1QPaDq51vXJcqtiDeh4pO/dos5mwdpNjAcEilQgyv07RglwljGXuFa8tHyH5IVfbC4IOyYIhZSmM3X5DxTB2wKmyUh6KtQDIsT3yVtC3hFCclnHfW0mEIv8IniVsAiBPCrved/O9zzwtIKXB6etkzOXOwlr1WzLWKYQqBA7G+9Bh0xYWSvknslSihbJqh71xlCn0UzhbiSoTtWq0V9m2xyRqTORpPp/H0YIEi3PKW3FOosUd8rm4X587q89B0l8iVvTw4rGQY2wIIXTds2R81+pW3qIX+b6FNxY4JsMyzkovD9q9pHZSN9q1kftjDwj8ZUfAEXAEHAFHwBFwBDaOgAsWG8fQz+AIOAKOwCAQMAKTRwhXSAPEBgQKSE7IMgo7hBEcOA7yiljVEGrs7OOHKD9AIQHZFVyQW+XfEBYQfuz84zV2L/OY7EZvi0F0yCaco33nqiUHt8vspoTomwDdJac0MtoIF+aMJfu1xObFnGJ8l/NlPeIcRDEiBF4T10HtyIviSH4qvECPV+YzylvRVLij/MKcJT4418OrAmIY8h1iiDm8StLkrYBtTdcAP+pOnP/flkEMf3GXM5BQG+8RMtb+g6xIPt2jsEax9oAr6xRiBAQg4VW6FTxV2PltHh9r8W5gzWOtpO/wqoCYR7BYTax4s47BA4HP4+mAWWz39ZC4hWCRxrXKQm1P7dTkDftq1eqebGTy6rHRkVrcGNkfqpESBldGGtXqsSxXEKhc4yYPVyw2tUan6bGsEolkj88naUY98JZLJFo01yla4GnB/eWdMtYkxIpOwYK+IL8H5OstshP6jCVC79pRHSFpNluQA1N+wyB8fUH5HK+dXuUP9cb/kCFUMBdXGqMrnGbHvWXCI/3BeoRo8+QerQA/uy8hXFjIuqFqdJtogaeF1oO8lmaFt0VjqdWKJVbQ1rNa+a/Qys+aeyLNMr4P3anHeytxPLvUTNa6FrM5hA0grFl4J1C6rSOMM9Y0Qnay1i0Oi1jR2YmbHaJqqAaNV8YRcAQcAUfAEXAEdiQCLljsyG7zSjsCjsBuQsBCGbXlYIBw5Qf4h2T8+GZ38LQMsopdtpCg/HC2Xa/8+OY1diojbEDmWPJafmiTCwPiDvKCH93s/OMaEF9GLPUbw3k3Qb+lbekSsmo95OeW1nnILmYiBdVi/CLI8RpzxfKC8DpJm9nND+lsoWyKJOaaYwhDq+4oNfJVj8ux/3Odv6XPzyhMz0MhUa6KlsJB3a3XyGNBPZh3lreCfA1cgzkHSXh+CBJqb6QrWV8II/TfZXgpIJC2F2K2kxfhjbKW8CJmfnMFoo7d9+zmJo8ABZEDzwuI8We3ndg8kn5Rr7G+/ScZBDqiRbFzuUejTLhiNzTrJKIHayDrI+H0Ogvn4fswffb9ZV34m5BItsYSNmjNpQwHxeeUBzid0NjTbnCNpZGxyero+DVjY9W5OF8cW2gqh8LoxIO1WhyPjGg4abwp1v4NSZ6lSZqfGqvUopaeLiyGExItCP1HnfG0WEuy4Av1L8ND4WkAnohNCOGIOe1lWn+wIx9PEwjYt8tMRO+JhUI75fKs2GzBgv7hXvZ4GfOduuMV0lmYf4RjI/wV7YSEZ8f7qmtAzwYO6RuMzx7eAfQF5Dn9/f/LSEb+HV2aAZYkiuY4xL03yfDOGDqs2kQLhIiFVpJq5kSsCRWt8czZXK51iTwrFnSDmEnzfL4SxbPysphRPotUn+/XW8iEMdYO7i3cV1jvuoWy437zKhkCd+EtuxvH2ZAOf6+WI+AIOAKOgCPgCOxCBFyw2IWd6k1yBByBHY2AhdPgRzckq3lM8JwfwTfJ+GEOEQsxB8EHKQc5Oi3jc4ShsdBRiBIQO6z37JTmBz4hpsh7wQ9sCBx2oS+JTHPRYkcPnZ1d+RVCPlm4JxoIacS4h8BGjGNOYPwNQc17EJi8x/jGq4jd5JB2kFSEQltr/paHJU78k2jyQ+lxJS+dCftEic2KxuP8zDs8DyCpCAPCjm+uBalexAffKWLFKoQn6w/tgeAmTFDnjnzWF3IHID4gqq4Wt912ftO3RdJfGV4pN5cY6qFYszD6kvK7MrwxWMNMROkWugYBCY8zJAbWR9ZMco/0Kn+pN14joy4k1DYvDtbSDa2JEKt/8iuvCvXkvNbhaM/s2NEDY62Z/aEVH5mfuOIK5QU+URsfa+WLrYnGaPWBSqUyN1qvTMrH4upWFCbHGtUgonV+bKQ2OrfQPFCrpZ+ZmV1YkmhRkMhriL1/SdvLmPas/8wPhBpwIsRXe2Eu/ZAMMYqx/ucyBLkVcZFokSJaIF6sgPt632INgFCHeEeIYqf783qcDKEC0QUBv/ByGtYd7+sFo/1zK4hqeNUgqhKGjXULT8sXtn2WccAaiicScwXxkPHPfGe+bUY/bqjJpWjBOsBcaMnbwsYyHhC6J+QPKy13EsWBkFCtJbJ0l0Jftwt3EXu4l7CWgAuC3jHZD5TYdJ4CD7CXyrgH8RxBduiEng0B7h92BBwBR8ARcAQcAUdgixFwwWKLAffLOQKOgCPQBwL80GXHOD+U+UHO8ztl/IBmFykEE8QafxO3m5AlxOZmJzHkLcQir0Mq8cMZAg7iiV3MiBm8zw9xRAt26nI+VIummNxeu5b7qLYf4ggMDAHzpjCBwkJ4MBcg29jlihi3nHh1WYRjjPOc3bD8jYAAicVYh3BiLhREq8Z62o+nBcc2X78sQEQNkfAVJW2dL0g94pcjVFhOEnZyUx/IPUj0InzOThEr+ug11gXWGULQEWIJnInj3lnwYIAkJsHr2T7IYbAFs7fJ6L/vkpH0udtuea5FrH1IVEQRxgH1Yf1izSxCL8kQaG+Vsb6xs3wlsYJz4sHxYRkkuMXvX0+uikvAwMPipo//aF3bvY/cN/X4qYfHrj03trB0drL50KMW0mMTeW306tGRejraqEfNvHK0XqscyRTTRi1ZiOOwWKtUl6pjebVRr+gctVR5LqqLi62jed46LVHjtM7PbvF1E6OlpwUENjghOJE7qVvBgwF8yMvCvKLfVryuxIp116tHHWxNwOMQYYu5960yxmO38it68XfKPoWsP99tPLZ5wXAO2tUukF4g6oVzj8vsjJfLvkZIRCDEi4L8MCTiptgGBmvMtJ58nwxxijBaK+aP2S4ESsGO8GiMNQQp5bbIuWeUnnUKrvbIKGSu9CtAMgYYX4izjK9rZYh6CDndCp4VYMa6iCfsSh5m2wWXX9cRcAQcAUfAEXAEHIEdhYALFjuqu7yyjoAjcBkhwA9rSFpIUAq79iDTiC3NzscPyth5zE5iiFgIJ4hSiBzLU8FrkLUQFBAO/I14wa5Uzgvpy3mN8J3rN2TOTu0HkaiQGTeIvAETQmiQQJjkq4vlDktEIggxRB0KeN7BbuSd2uYdWm8II/rKBAujnegf3oM8xZuB8Qzhyu7wp8kgrdgJy/cbSOfHyPgMxCOC3fHy9UU8OvoRLRAdlPA5VWJtxgCCIKGCuL6JfUa6Q+gXu7j1mX5DjgxV96yyQ5u1gnByb5CxDrGGgHl7gUCGDIUoZr2hb4oiTHoVcH1YGHMsZN9rZAiw3yZ7VMeHWLu+p6wHIsOUaMVPxVdLIGqpz2vFmoZYxS5rcmp0E1XslJCxtIU+M3GXfhvIXFd7ogc++NJqGtVGzzcO1K88//HrR/O5m0fj5MY96bnnZAceNRpX9ypkTauZ1+qtWqW2EFcqtSRJ43q9Ukk09BdCokTc2c2zcwpqk+eNJMmuaDTif47i2szcfHMggkBJZDOWmR8IRpCv3FssVr/hRRgcPFwQy5kHJtb17Nj1vLFC0mPuZazNXyJ7jowQRr3Eiv+l935PRn9yX5z7uZP/GF75uovECBMmaIeFBLMcDrwHvtjQeResB1c+U3rVcO97ncyS0dOnFDxo2gseLISQYr59RP3C94SeWKwnZNp629H5uVK0yyRc2IYLE7cuhCZbgzeSeXUhcpOonHsLwjf3km6F9c5CboHtQh9C7aCa7udxBBwBR8ARcAQcAUdg1yLggsWu7VpvmCPgCOxgBPiRzQ9vSw4KEWo7CCHYp0sjnjixxSHl8KiARLICucjuQIyd4JCs/AAn/jzEAzvAIWogKSB0+CwEBiFz+iJyhxlfkSu0BQwRb8CMsCGQncUue70PFpBekN579bcJQxAPCELsImanOILQ0/U+OIKheahArFZFTOxIYnqY+q4td4tVi3FphJMl1kW4QJzgkfnBGKYPwZ++gLxkZz1jnWPweOCz5p1EP3Je+pdHXienRb/hofgc54UQh8Bi3CBqQXpTF0gr6jEQEnmY+qetLoY7oeVYm26TdQoWHI53BImrj5LPQnOEfuun0JesW+S2+BYZO7spnaIFc/DzSqvK8+WX4uvCQQlK1yk7SUszmboRDsqI927X/iu9SLx+xA36lsLjhslphAqdpwhbdnj2E9ckcf0LJ5f2hmrW/JGzSw88Jq2NhXq9Hsabp8N85aZTWWVE+barlUajNquLp1mI9yo01BReQLV6nLSSaLRazY5pWd5TrcQPxHF8ZyWOFh5SLpbZOat6P/D2PqYULTjZ62WMZzxZupWf1ovccyz/CCLTZq6BF7DUdfACYJ6zlrOuP6NHHd+t17mnIVx+4P7WLbO/f/oPO/vVBFFet3nNa2DAo4112kZfrupRsrEe2LpPq6+bmpfMYe6LhPoiZBZeRrSzs+CdBOZ816CvTaQdynWuTZRYzzym/Qh13FcQwhDI6P+vkLHedyuIpnx34jhEXL5frOfaWzcA/EqOgCPgCDgCjoAj4AjsEARcsNghHeXVdAQcgcsOAX70stsTYoAfwZBwiAvEyudvCDvWcBKJIlZYEm7eZ5cf5AKEBMQOSUchDSES2SkIycrrthOd9yBbOT9E7rzIsoV+dp8PS6+IgIFkQoyBsKYN7SIF4ox5nkBkQ0j8U/kaJDdEBbuxKZ8vM+Kbcz5ZBhkNvhBlEBlcpxAvdF1Ia8gKRI4TvrNyXSPCiLJOoYI5QH+COTurEZEgh0j8DLFE3xBOCDGJ3a+EgsLzAS8AQsAwfyBXCeNB3zFfOAeFPqN/8bQgEfeKJFPpZQFZh7DFnKT/GVeMDeq0qGOGksQr2xuUU6DYUT6AvAKsLawh5Jz4VdnXyhADrbADHk8L1qmK5sjfrUHYA2PODWEOec5cfL7su2WEjKLQl8slDt+k/78w+1z4t/E14SlawZ4VVbTWVYt53I2A5Zysh/Q3ax59yNqaD2LulmIFRCfrBevrUyp58uLR1swNSaW+v5othSyeCHl9bKke5w83R8ZnopGRfUmeV7M0NDL1UD2OCQml0ZkvKva+1IrKZFSJFOkmP6EwUadarbzaSpKpvZMjZwclWFzAc/m+gXcL4W/wkumG4f/U619T4oaYTrjCzRItEBOY34hWiIVfLOMe95K2Orc//Xf647hsT5I3Pnoquf7c++a+jXnJ3KfPeTTPCtYQzk+hv2grxDyvsd7glUhf8rmWdu9bvoSul95hIaMQpcDxj8u2slb+lx6YMhcR718pY11lDeV+x1zdTeQ89xXuIawzfEegnS+Q9RIraD/HcL95p4y5QKLt3YRJjyHhLzsCjoAj4Ag4Ao6AI7D5CLhgsfkY+xUcAUfAEVgvAvbDl1BQtovvs3oO2QBhAIHDj2wS3UK6QSa8Xcbn2AVOKBzIHuLtE3uc53yG3eb8KGc3KcYPcnakQs5AEPLDuyUit7Uakbvehm3C5whfQju+VwYhBRkFJmCAWMEjIs10qNQXQtrEu6LwKJFBXD6xrBPPIasgGyEtIK/Ai2N5D7ECkYLrIRQh9oD3b8gQg/rdTb4JEAz3Kbsk1badzEaK2k5nxiT9xevgiSjBLl8S5zJGGbuMf94jbAkhakxQoi/IMUGf8xn6iO86iHH0D8QnogNkJOPcdlL3QzIxViDTjaxjHg4kfNAgek6CRK/TGEFbPHLcBkULsAJLdrJD8L5J9tsyyD4rL9cTdh/jwXCPRIu7ROT1K+iAKXON/gVjkmKz7kGgX1zo2Qn1aVM7/kUnR6xuvcuH9BYhoOh/xpjN/YEkYpZYYZ47rBuILM+WPRTl+VNjVa4iNULJt0Mz2xfmRq5otfZcdWKkXouzWrWStdJKK0v3VavxovzblrI0kzNFPKbcFgItS6uKEJUm2b485PJAyZfmFpK9mk8QzoMu9C1zg+TaCBH/WkaYqM5Cn/9HGaEJWWcfVB+DY799fMkJO0JBmWcFc521GdESD4tvkLWLY+3neYv+gFgvPAFOJjeefsvM/xNOtm5mzeB+wDl5bqGuGJuMIMYBwihrDu8hQvIeaz5jkfWH42yur7uNlzR6gC+U8z/qZ26XpDqE+6xw5/sF/Un7vkz21V2qxf0S+wsZngTgDFE/GBefAeKw1lOVmx2499D35KpgswPfmRBqbO3sPC3fudj0cJuMdY65mLpYsVb0/XhHwBFwBBwBR8ARcAR6I+CChY8OR8ARcASGBAGJA91qQuxyI0gswTBrNz+QIcggCdn5CcmC2ABlx3uQZuw6tx/i/A2hT8gVfmhDNJC4FlIGIQPyFhKS4xBBIGXjfnafbyd8IhtoL+FfnieDbLBQQGBj3hG0aTaM3zIS4rGJsO+LrwqV8WaoazN+8+FWqE3eGB5+z4Ph3O3zYenu6bLtdAakFecHf8gcsDKhh3NC6NEX4P/TMohZQqW8TcQFOHu5FAEb5LbTGVwhES3UE+MZwhT8EIogqi10GcQir0Gq4UVEXyNUGAlpwgeiEoX5APENsc78gKieLs+PJwbng2wlCfeqoaHKBNqQfBCYQ1dEVF6oU3si4Sc/5qoClysPTdoO81zkppGveT8EZ4/Ggh0eCswL8G0XLPgIRDPG+6/S3ChIvV7AKbl5e6GurFGIg4wH5hiCBTHlD1nQJQSKila5SFeIoLN7lTz8pj6D4MUYQLig3muKNS9Bolux0GWMQcbUtAxxjLUW4lfXkwRR6GKkzV4II61zIUpm76lXq3c3q7Wj8p6I4yyu1KJoshLLIyXE8m4LaVWeFdU4ThebSSrRYzHJsgmpGJPSOO6TkLE0NV5JX/ZlN20GeU5lGeN470Havlj2yOB6BIX/rKcIQCTqRrj4sPqYOTmIXeYmOiNO4FHD+EKI7CZWWM4UBC6E5g98aP5FD7955kepKf2N0SeMIZ6zhvN8Lw4smvusNbSZtR6ymr7kOfdbPLR4j8/zt3kV9CNwPoLUFj7Dk2otc1r3qkT9BoYIEXfL/kz232Tc/zoL84/s45bniXlkwvMWtnLjlyqFCgsDhVjBvcSERgSLXoXx/i4Zc4PvSayDgxjzG2+Un8ERcAQcAUfAEXAEHIFdhIALFruoM70pjoAjsGsRgByBmILAg7yznaFsqeZvyAZIQWJ6E/6G1wlxxM5JSB5IBYgkjm3fUQ7BaB4bEMaQMZAyCBiIF4VnxzCJFiIZ2AULKYU9VoYoA+kAPuy0R6Sw0D9nw/jNV4V9zxFTeMWVoX6wGmLxVQt3LoXRG8ZCPJoUIkbrVBbGHh2F8cdMhJnba+H0/6mEqvipZA7iCizBbHn3dHX/6ZAtHgrZPEQ4WEFMghsiEEQYJOXzVU/IPogNCKC7Seqtx8uylJ4V7WGf6CvGG/jarmd2QEOKQvrSf4xnwp5BQyM84EnBc8gywv1QIB057htXABavI8g1CEiECwQPdlMzH+gvyErOM5D8BSvUY0veQqiQMBFPjjeih2cWKyONamVhKYmWllps5I/3TY1AzCm3c0x7i3aL4MwPz0GJAAAgAElEQVTWQnC2NYR+ZH6w/iA3sNbQf53lRXrhtTLzaOmXZF9m+ZeFJebS72m03KPRcTgaDd+HWBGJYox7BWzhw7NKJF3V/JwNt2vVvD0a0bM43Esc/wF1iJHbjLHnyhiPhNlhDbW8OIrulJPDIkSt2dNJY+8nT+979IcWJq+ptlphvFrL5uRNkUoerqFtyMtiRKGgEIubWZ61KpIw9P5kIw8z6jdFj8qXpiZG5HURx+q7WH3XL55raTLnZI1j3v6wrFdOi39VjiOSXDOXyY2wpPUPIrcQete465xzgCHjiPsT6z2i1y+tUHnCszGeIdw//onFL0WsMG8XW1d4RNDg3EIumpAodEjdwnyQ+BwtlaKl1oRcGBceGcwPRDbEG+6FrPP2uwnhbahEi1KwXG+duD9xz4J8xxPxx2S/1gNz1uMfkbEe/4qM0G+sA5sVFmyFrl/7W6VQwThjbB0o20tb2PDAPF5JrHh1+T7rEd+nwGtovOzWjoZ/whFwBBwBR8ARcAQcgeFFwAWL4e0br5kj4Ag4AgUCpecFnhb8CdEGGcSPbdv1zyPkGCEaIHdIhAtByzH8AH+WjBAOEIsQadMyE0EQJtjBynGE0jDCgx/yJnBwzfUSIQPpRZEMEFCIE7SNcD+E9oFsZkcsdUV4QRwAh/kwcv3V4cBzG2H88yQ+7NsjsSIL85+KQzRVDXuekYba4TgkDzW1tb4ZJp5yIIw86rCEiCwc/pZ6uP5nRsPiHUk4+74kRHURXMlYiEazMHLtbEhOT4bmAw+FsesP6r1rQjrfDA/ftqj0zSNh5h8OhORhSA9IcupBLP/PyD6p+hNC4uMbCZkyECA38SQ9Qj5xRfoOYwxB8EJs2Y5mxii7l3nkPb6XQEE/SYYXC6IU4xOSjONMrOC8kI+rFXIpQDj+vQxiDSKUcQMZazuuOU8Rn759F708KgI5CUrPitWus+3vI1bsmRypLrXSRmWxOVqvVbQRv5IsLLVak2ONqFKJJs7PNzMR4hIhQ4yYIdIbvBMR3wvrFC0sfBNhUUjc+/UyxCUK6xTiEDuXyTnAbnXbzX7JelLvlZVg+Vyt9FPho8pVcSY+rHB3NRGFefj+yk3FmOhZsk+HR0UHwgP5eXlm3CvPiizMpXeEWP1aUb+ul2hkLC8Ho1pefxCJIect3wpEOzkg2kp+t+o7H+dJKx3b/6bFQ4+dCY2RG6oj1Zkoj09KnpiIo3hEznQjAiaWSabIpVuEmhJwJ3EUzsvj4qwSWcyq7+6qVfHLiLrll1gJjrW+Bz7cH9hxz7Ugqae7nIT5Q+gojHWOufYn5WcJFcV9xUSVle4jiJiWWwkvKgQw7lvfvELFqRtebXgLfkBiRfLu868wMdTWE8ZIkVxdY1/iUZTqv3FV5JBwlcV5JqEoyzLutS29rqf5qPqL5wikeHMh+lMQOBBHCs+s3VLKpOsIOrQT/BB0STZNmK1uhWNeIftK2U/J3qF+Jp/DQMKrbRaupVjBeGVMcI/mewTCOHP2VhlhBHsVwj4izDHPPyFjXK93DdmsJvp5HQFHwBFwBBwBR8AR2DUIuGCxa7rSG+IIOAKXCQIQP+YlwQ9vi8HNDkFEB3aRP0FmO0IhgiEXMAQNdrEjXLDDkB/tkAx8FlIXon26PA/kLsfwoz5FLdnKfBYiFtj9Tl2oIyQW9WYHM8QTbaJuEKKECLEQQrRjIRx4wd7Q2NcIE08YDfUDe0My/+lQmzocpp40FhpXj4bKmPCrzofoSSK08krIm4uhfq3Om4q0FoUVUnlgXHdvmHjqfoWLb4SZD54MjSv3hkzH5UdntAH32kIASWYVuOVsFI5882honXti2Pv0KJx7X6rjpyRsfDrkGW0glwjeIHi/vF3tYicqZDlkx3ERRdR9N5X2uGY8h+hkDPEcog9xidcYn/QpO3vNQwYykNBe7GQmxAwC1BeVWNHXkEtrLZanBaGC8WEx6gk1xHVtV7A2wT8SFgqhQsbcquuROZeI4N7WHcQSJFZqe+FZMbfYqtUq8Xijpn37eb5fczYVD7t0dmYhtFri1nLt4o9DfXy0zhuxvC5mtdt8YaRebbaHiep2oagMOdWRa4BDwRgxAnzbPRfayTySIUN+4gUFnhCitpZ1Xs7GEOuc7bjfK3GiUXm0BA/xyrLJnnIVvaSezbiCVr3snnA4PxO+QtLkexEN9Cqk+mfUr9SbsUY9rS7dCHUbx8V4kCEGM54YyySBfraM87I2MV67lavFhr8tr9T/fPHI4z+cHZiejGpjoVobUV4KrWNZvlePOnfUStI0kRoxSoRAiRRKxp3NqsV3VuLonmo1n5Fgsai+W0gSUnRvegEX5h6JuMEK8RtholdBUEZkZP4iNN4mI+/LspC8jLX1K+c28Qds8Wp4usxy2Xy7npOzole5XW8gVhRi5Jn0miDBIjyUXMfnbc3hvNw/NBfkXZWFfXFNhHMWj2UhPyZFSLJdNKI5MpJF0b3yaPmcBI0bVMFRYa51Ote9rxCkyKGBhxD3yOL+qSTbaxbxV8ozs07BcAV41vwW7eG+ROg0E90Jt/hmGeO+WyH8Ht4vJGL/TVmm9YHvDrb5YcsEjC7rUnt9mSs2fxHE8aJAeEAUZ2PBC1dA6716D/tDGRsjGFvuWbHm4eUfcAQcAUfAEXAEHAFHYG0IuGCxNrz8aEfAEXAEhgEBiAUjfnjkxzOkEt4TPP+YDEINQghRAyGDnc28B2FeEDgyzgNxbKEyjOThEVLOwjxAKlVE6KabLVqIdOC+9BwZZBdkgnmSUN97ZAgUvAZ5Rnif4zIEgc8L1ck7wlWv2C9PiHGFeKqGpfskNByrh7HJA8pZ0QrVg2prrRlqI+winZbRLrWzDhmjXbQ1rg1WwnG0GmoHIVc/ozBSUwofdSwsnlDYluoB5cHQ5udkKcQT9ZDukQAyEoXquatDfX4qVEfOh6kvPBnOvveWMPfhxdCC97mQY4QdqwgUEGoQ9fepvfTVO4gjzoE7vEAKtRu4gjGY8kibIYrAGTGC8ck4gwSFECQkCccypjmGeOl4VEAMr7fQhxDJXAsSlfnAGGK+IIZdJFrobyMhed28PxA5GiK4EfeYRxdC8OCFsVVFBGnXS+FZceP0wUoryWpYrRaPN1vZvvGx2h7tFD9cr8ZXtJJQmZlbkpoRn280akvKi7C4uJjcn2b5+Ynx+kQ6Vm9KxIDAB/u17hoGM0S4d8kQLUh0Duad/fadeg1BFfxI3stcYP0xAptHE7hYgxg/GOsV4+CIZs5DMnbfI15d4l2RayXLkV7Vgkw0eS5ZKqdVmc6Th1eVAH6vHiHCIZ7ZPc9Yw5OAMUH/Mk6RPUwsYX2kLRDXjE+IdT5D3ambeZSsJD6+PsqzX8wqjeb47N3jNSXXXmpMKLxcfkbraivN5EkRZUfFjrckONUV+kkYyd8izxfkGSNconoc63p5kQ0D34qkUVMYqa0pXAes3i5jThD2iQQRrMndCnMarwgWPzClD7kf0bcWRsc8bWwdZ47xOcbOcRmeahReQwTrJMw5L2OJMQeJnH9s4SslWDzXxPl27ys8Va6Wb8Wj1aO1LM0fJREiF8b75Kki0jqPJAbNt9K0qtcPCu+RShQWEJIkZDBWyXPBvZAxzegqrqF5l69VtGjPM9MB3JrFj+7Qb/hV6sGMQe6z3DSIcHjX9Aq9x5zHo+hrZIRG5P76fhlC1Ud0j5vV/W2rxmo3AJjHjB/6j3WD7xZ4abKZgHGGV2qvggjzczLmPCI3YxHrJbZuuAP8BI6AI+AIOAKOgCPgCDgCywi4YOEjwRFwBByBnYmAiRbtoTYgBfgxze5GSBV+oEM8IFRAwFkSYogEEkZDtPGjHbKRz9nOQXaScn+AiOB5ES5ns2ESsUFyV0gSQk38lQxigb+pLzs5CREC0UWdIMtsN/e8xIo7w/U//9xw/iPHJVhMhvHHjivoy5kweuNSqEx9NlRqTy3bBDHGecHGcKJ9EOYQkBAbXA+CEgHoujD6KAiYPDSu+qeQpTeE9Mz9YeF4LbTO7lU2AAkYe8dDdHpPaOw/F5JDUZh4+lVh/IZmmL8nCSdf+/Ew/2lC4kCUGDlLP3BNCJCfkF2htrMTlXATO67gmaBKm9FfhcAlw4MCPMGSsQVZyWu8TxgO+oJ+xCOIXdmQwfwNuQlBTZiOjRYIUApiA2OIcQ/xzPnZoc04oI6dhBr1p9B3jDt24yKoQHAPjVdMmVw7RqiYlPCgWDYHRbreJEL8qMRF4ZnfGFfCqOjvqt6bTRLlQYha55ohnllqJbEIc4U9C+nM7JJEDFwwQn7P/eeylYhYjdNuJYeY1Bt/Wb5JgmzD0I4nXBSGiMR4oU/Ak0cK5DVjgP6hX+gvCEXqxfxk9z79wFhi/TOh40J9suNaGxY1fjTCcq0S8qroJr8Q2sUKuRkQHSzBMjkLzFONOrIG0C6O+QIZ44EwRdQDrxHWFSu9wlMx5hDLHoxq9VQeLQ/m+48dVMwuOVPkU+LOD1TSfF7+PfKtICxR2KMUFggWrTjkCzqeYIDNJElZr05XK5WlahTP1+UVM8j8FT361drWUv8iGLMuM59ZE79W9k1t7W9/+lXlHy8tHyH6ETrw1IAQZ54TTqvwXpIhZLIe3NrlfJ1ixd/pGIQKPHYYOwV5/J7z38W6Qp8Z6Y7YgTjJenuFDtpfjaMxTELQpDzgNF8qo+QFiZXtvJbnR8gPonmjmFHKYyG1QkpHU54Yp3XGUzqpeSEyHjc7HFcPWLfsZRMuwROPi/9WYv0DK9SAjQMYHhaMD75b0Nd34lk4wLwx/YBAvVl/zDuKMcDfbHLg3oP6i9djr8K9mTB3b5PxPQiBrD3h+rAITP1g4cc4Ao6AI+AIOAKOgCOwIxFwwWJHdptX2hFwBC5HBMpcFp1NL6I1lT+mLeQGNB3kELthC7JGBjlkO/sh4CAVIGAgdSDC+BuSwn6Y8xwCjnNt6u5/kRnscFz2klgmCyED2HUPuQDxATkIQWS7odkdCVEFcTkXDnzFWNj3vKeFqaePh8knH1UoKB1fuTtMXf0UCQq0A3IC4uS4jJ2SFnuatkGSQYhBxoGVhRDheDw8OAaMPlNcL658LsSH5F2xd39IHvhAWHoQQvzm0LhGBGttf9hzRN4Wo+qPbDHsuXVMYsfBMPvBT4cHXn9XWDrB+WgL54SMpY20FdLznHCANCVBN0TJUJcyX4WFpAEzntMfjDmEGdqJOMGYpB8pELfgyvsQlrz+IRmCGrHQ+QxCDrlKBl0Y81yPXd+MZ/BnVz1jgf6nnu2F9jAWEZpoHyIZY9HC2Gy6gNcvAAf2jimdQahrfdirvBRXzS+2rtcLV8u74irtzT8QxfG8+NiqduhXG/VqroqPLiw0pxQiSlx52H9ycfakBuES2/j3jDeWFFqK/lhzUuoyDj7i5x/LSEqL/wlzurMQJ56EvghA75SR74CxQn+AO2GWwJq5hXhB3yAWtBPXl4ZDSsPnoqlwe14NaXYiXC8p5kl9yKzf3Va5v9Zzxse3ySzUEOsMO8xZQwglA1n/fWX7ENnaC+O/vSAW/77sfTLW1cVk4sr5E9/0BhbihmwqjtI5pRNJWnm2pL6oVavRlNQJtTebE1l+Tow5/VLTsYt5XEnyKD9ZkZdJpVJd9hvZ2sJaiqBj9w36DjIXj5fVCnOJ0DsImoR9otCvCDmMEeb+aoW+eKMMzwo+B6nMOYw85tHuVQheiBVPkwDU1NyQ0BMfkffEFRJ8aho8jSQhPBrTIcQS8xo6ZhzsdZKWPrOkG84eZQo5qrviUQXfkp6R017GoN1vwWNg90aFizKxpSsOK3hnrIbbRt4HU9ZI8MaTBcyZH4i4vQoiH8cwH5gvfPaDur8RNg7M+B5iodhM6M5WEcz6aYOdiz5inPG9h+8NGGOUewvjhflsQnav87I2fUDGPZl5zLpguZcu+cwA6t5P+/wYR8ARcAQcAUfAEXAELisEXLC4rLrbG+sIOAK7EYEyTBPCRfuuPwgBfpxDxEMw8aMbcokf3ZD2EEi8b0IAP/Ih7BEFIHchkCAWOJYCQbYiobIWbEVeQGa8SAahgVE3yDB221MviCTIAuoBycGue4q1h13uk8o1cU+Y/tGnh7EbFHN8pB6iSYVlKkI7sSObz1N/2kb9uQaP7eFeOB87+SEjKVyb3dSEAIF8h0Tl8xAckCBc96w8NkZC5Wrlyrg6Da2Z4+JfHq9w562wdO9SiCYqYeKxk0rULep07qFw5MXTYc9Trw/3vTYLZ996t7QMcKRutJHrTcvYNcze9YeEDZ4vECRvFBFCfYex2A5W86awEEqIO4w98LQQZQg1FHAEV8hwSGli4UNIMxboX8x22w+qzYxndm/TjyTmZTwRrgRC3AQI83xpvyZ1LMJ2yRgvFpedtlnemEHVcUPnGR9Dq4hG5haaYxIpDspR4jEKe3Ok0aiOiqStkR8hrkRprVI9Pze/1FDHKU9CXlNYqCt0/Iy8Mz6rziMhcbJY017/PK/+6hs/8rASdLfWGvKmFC3A7i4ZoVR+vsS/WxsRpphPhIeiD1ijEElZxwgpBMHdb7lfq9VpJdi+XavFP2sFe5xGoUIo9cwp0e28X932IrlUMAo7zFlP2kunWMF7kLkIw5RflpGYlzGEeEPb5j/7ineZ4IUoNCcx6W75T+yp1+IRheeSKFY5LxVpj8IXaR2J8LJYIGeFiPOsGuXzWRadlD7NWJ4fpHdFvyDrONZi5jChf5ir3FtIroLHEutXp1dN56lNrOB11mbEWvNYYp61h3Kyz3INQhIh/DD3wJL52EtUYw2iH4pcRyqHNLaPS6i4RwG1rlWkrbEQx1lFq3OS5XGSZjUdk8VxnMobKSFEV61eSzWPiMk1oWCIZ9IsmdS8uU4DEyGE+oJBjIfTWufIGrAelkPpc+Ynj28GUxleii+Q9fIq4n0K8wbRDrGCzQHgh3DMd4y7yz4sPJxKwZ75YXPEvN7MS8K+f7AG22vmacW4o78ZU494Rz6yhjOXzetnJVwRFv9Ihihm85bx13RRYiXY/D1HwBFwBBwBR8ARcAQGj4ALFoPH1M/oCDgCjsB2IWAhUuyRH/X86If8hvhmzTdvC36YQ5bzAx/CAIMosN2JtnsUIprzDSxms4gJSGPyOTxfBhECUcVuWMgPdlpjvG7hQsATshnCgzZBfkyEK77+U+G6n3p+GDm2V+LAHRIRICogvCDQ2LULoQWxRVgZiEPaBFHCeSCrIQ3Z7U0x4gU8aC+kF48Q74YNeOEZgNgDOULIi48poTe78OdCltRCND4RWnfdE6pXqp7JVLjihQeDeMYwcl0jjD3qfGj90E3hnl++N5x9R1NihiWBhvziXBbnHeGIOpLA9C0iSuiroSgi8yCG6BcjjBhTvAYutMf6zwgk6s1rEFg80vf/LEMkQqzAKPQFZJYJR4NqL944FK7L2IdsxFsCMqogHWUmHl0Q/JSbIlfOCt6HrEZ4ob8ZE4wBhLVhKfHSUjKiGPxTIl6PKNn29Y1a5UrRtKPytliUF8VklkcNMa8tJXCu5K1E8fjDUr0aTaZpvGexlT2kz9KfzUq1oig4+ZzUDOUfjthVnYmQTddKyJaiBTgTsofwaggSnfksDD/EubduAExyKbBWQGKORaPh7dlCuEPeFR/Q7CW5NmOO+fQSmeWaWOvlOsWKXp9nXL1JxvrAczyKEDFYa0janoXfpToh1W56xtHd8qI4pb46pnl1gCTb6pvT6owJJX7eI+GiEDYlXkCY5kpc8WAU54sKYWTk8VrbMajjGS/MV9qHMEVuC7DFo4b192dlrIn9FMtvwbHdxApeZ65SWFOYe1zbwvO0XwO8OIeFDMPbh/Vf60qkHCZ5LERbCrqV1uJISen1ThqW9DhCBDF5WcwJ25Zwj9NEx2ZB8yYfV76QE6V3I3sCwJ71gusP1MNlu5Nur0LIE/KN+ymeB4xp1lUeEQFWC933HTrmObLXyxDmCcXE/f7XZawP3PsQvOhb+toSdnPfoy+5b7P2YvTvcRl9zZpCH9OT5g3J/Zv6cF76CS9GhLTV6qhDwi/IyCnFOGPtQJDj2gPtZy7kxRFwBBwBR8ARcAQcAUdgdQRcsFgdIz/CEXAEHIGdhICRriYw2A5ERAGILwgAiADCO0CQQ+TyIx8CjWP42whcfrhbCIcNYyDCA7aOUDzkqkBE4FoIEc+WIahAYkAEQUooB8X4uTB6w0RoHM7Cni+uh5GjSyGZxatiMozdMhka194kkYLPQSxDWEBoQEDjDcEj10OIOC6D4IBsok28xy5PniMM8Gg48di+S5i/wcwIMsvLwDEYoWK4l84oIfcp2ZFQe+wh7d0d0RmjkJ1fCNE+5bhQ0J6R68ZC9qnFcN2PXxP2fclcOPGri2HxXiO/aDvPIfAJPUIbCJP0WOFGbosTIpRo57YUEXXmSWGiFriALSIAhbEEgWQ5U9jhTFt4nePoU/qA/ub19t3ztOtdMnbB9iItN9JuBCwj2szTxjyIILy6FhHMzVK0oO20gc9y/MDCwGykUXyWcFCVaqyw/HLnqSr7u57UapWFNM2qskPatT8uJjYSEavxqGhlIaopOL92jSs+VKWS1pWZJa9EtZFG7ah2kzcXmskDEjlSCRcIe7aGdOb3WLXaJNnVuGW9gYDEywKSEo+qfgueLcwHvGN6FQhz+oId0TZPZyo3h7n0wwWpzfVN5HydnrNG3Cr7jX4rsYbj8HogXNFtZb3ZPY5okxZCRffC64W3l0ohShCKSGLFfQr9pB398Zw8Aib1Hl4ImiPKDR1HkMYIIHWJHsyVIr+QyO4199Ea2tbtUFsvaQPtfFuJL2vit8gQpH9mg9eAEEfc/D0ZnnDMPcalJT3udnoTUxCZuc/dQTgoiQ8HcjlRaMmei+O8JWFoUr1CGCiBGkak0VWEPX/PSuBTlK5sNkQKGaUwa/rQ1Xr9lPJe0FFNrYUQ6gXuaxXzNojHdn+cPgd7xDj6gfmJJwLh2hAOVyrTevM/dRyAiPgOGfOGsJBPliEuMr4RRBAP2FDA3GKTAvcSBAjuh6wPfAYxkT7Hc4e68L2CYygrrR3tVUGU/i0Za4Td69tzVnRU2/90BBwBR8ARcAQcAUfAEdgKBFyw2AqU/RqOgCPgCGw9Au0EvJH1EPaQPggUEH386G8Ps2C75S00B8fYbta0DD21rpaIvITAJgwQRDzEgxGMhIXhenOhftXR0Lji3nDohQ+F5NzBUD80EWKFGx+7ZX+IlUA7q30i7L/xSGgcgSCznBwQg+yepJ7s1rVQUrQRwgvC0nJg8D67+BE2aDfHQEZD/LUTcJ2CBbhxDGIFxxXeDyWGRrDb7k8Ij1oQi6xHEap7D4fW4qz279ZC8nAmAWaPQkIlYeJJi+FRr6oqSfjJcN8fyPPiNEQLnjB8Dkw4D3WclhEP/APC8D0igmnTlpVSqOB61MtyVUAG8tyS2iI4UFd2lrOzFRIJUQKCH1KLR+oNYYzAAZlpO7AhwMD1STJ2tXJOiKhBlTfoRCR5hgSDZGOsWf+bF1FBKDO+JVBcKCKagyzRa5BXfHbodttKsFAoGwXYr8SVhaVkSomZeb6oF+URopzaaTqjnBZyvIgntXN8f5pnoxIxWs2FRP2Sy6kirkueUJ6E/LRe1+cz+nKvyNvDCqPT0t+JvCzWRcyWnhYQ8fQB4gIJudnt/K19dC5jBRG1syB4HZcxZgj3RX0Zd6xrEJskrzfRdkF9x/izNc7G47frNWLasw4R2olzMuYYF/0Ursm1ITp5pI3MCRJKIwTbmpnhqdPjhO3rM+OLZM9F+Dphr/pCnEsljGI8jkyAZW5B3DKX8PpBIKQu/yLxAhKdtvI37bzkupuYA4Fr0Vd4W7A2so6RD4R5xboGrhDQ/cxrsOAcPy5jPaDQJuavrSW9MOVY8wjk8XphSf+e19TerxzaNyhnxf6slU8mUaY6RVrDlFxbanI5QnA1IsW5cljEWn/zs/JxC8pfoYhqxOdSou5lkZp2sRasVI+y6ut7UH/yQcYtpbjOJvbfWitJfRjj5HgAj/fK8GRBcCa3xfQaTojnBWalXdTk/JZrwjwuEY4JJditsPFhLQVvDwrzCtGE8cX9AfA3tX/XUkk/1hFwBBwBR8ARcAQcgcsVAfsyfLm239vtCDgCjsBlgUCZmJu2Wq4BnltCaYh8CHKIGIgviiXGtHAr6xYsRLRDrv2gzOK7Ez6I60BqfzhU9z45HHh+M0w+oRKWHhgPo8cOSqA4LS8EySqnK6F2bCE0riLMjcKnxJyrPW8CbaD+FiYFQcLIO65jO8V5DYKS42krhAsEFEQL5zQRopuHBdeDhDNRwsjGEqqC6OAYyI5i560MwgPyDYJ+XoLFAbHHSyLARtQO7XZfmNOG6dGw8OkkzPzDQ+He3/pImP0ImIMRCdMh94iBD0FjMd4hKn9FhCx13pJSCha2uYH6gQG7YBGzqNtyOKxl/CCZj5cYPK08hrAa9APEK6E/8LABe4hE+uI9Mo7tFTKos52QS1x/pQJeXJOE3oQj4pE+g9CG2Ma7hnrZTuGCnNqIILdKfTbt7Tf83V2xEmmPKJzNwYdnF2+uVSvX1uuV65vN9Gb13ZXakj85v9isa0COVbRlPKqEUb1Hngr5W8QLiBdpIvEijj6pL4T3NZPsjizNPi6wTui9GYkZENEFWbje3eSa/3zXtNwUYPENMnI8MJaYi/0UwsWw0x5ylLGCyMBrtqPe5l1XEplwNxIvmKOMUz5vO6m/XM8Zm5CXCAYIkOTPaCdOj+vv18hoB2sWHh2MQ8Yy10M0ZUwzphjThH9alcwWKU19OCfhxphj1I062JpmCa0haCFR/6asN14HCDaIAIgEjHFCrkEWv1/GeakL6xJ9x/xkjKebnfei7GsLzURbzIONNRqhyNYOdsFbqC3yYSBoUU88rfA2o10IQrTDPFIT38kAACAASURBVCvM40cvLZf2MEYS1uy+QN/Sp4+VYPFozYGGNL0jEiZuUadMKjTUlOb6lHJWjP1f9t4E2rLrrO/cZ7zDu2+uuVSq0lDWZFmWLRkLDzK2wdgYbDOPJkCThLWgoResdNOkF1mdJqFXQicQr84KBHDSDA2sBMgKBpvBYBvj9owsybJsSaUq1aCqV1VvuuOZ+v+7737lq6eaJ1XV26fWrnPeuWfY+9vD2fv//waZJslDVOmKIgjLSj794rCruCK5gnPHZeEOq189JxIwEnn0vHrNV3T/F9V1IKkg+7sX2ydOFeAsB2NBuIdrtZfaZZTq9kwb3wUIO7691DlxqLCW+JnzKedLcA11h9XXbiX6KZYZuKUzK8ozjiEvQV79K70ELkoCr3799zNu0DfZk8zSj3GSbVxJp/rMx37rnN+si8qIv8lLwEvAS8BLwEvgEiTgLSwuQXj+Vi8BLwEvgetFAgbGCmxh0YIGLosWQCyANkClcaAdcMnArvXg/HkXeRRY+2t1A1qSgHCAZ4BJJID8ntv+A3LEsXtKwatlhdCL3fRrF1zz9sSFTeUnPummXg8wiUsUgCsAcfLM/YB8AAymTYwVBW5DAE5sQQbJwEINcM/c+Jg7D9OyB9gyrVnuM1DMtLIpLzIwKw0AXHMzY6Q/IA3HBr6aOwneybmmiBYF6g6P600AdrIgUfmrzqrcXMlV1HdMyV3Ufe7ZX3zEnfwImu+AoYCRAHdob1udIcMfllzRPP34lQ7IPSIrkAmJMiJH5E6ijVAfgKS47gDohSQAtEIzmt8gIsg7pBGAK9dwH/XEuTcpnSsQKuAs8UhsOxtZgfb5PiUICsBe3FNRF8iTd1P3kD60GdriKU3065GsMIGstHtFo5Z2BMzuE8C6WYYT/Voa5audLC7Koi4vUYN+f9ApArmMKoICbfGiCuT+KYvVaMVx4Ld/rX+ozrcNwdmyWpVbKJsjIqczuTUaq5rTH44sLZA9/QxrCOrpf1SC7Pp5JQNW7AHUESA1hJL5kqfPAWx/elRv5GmYZUvnCoo7cs3UFnFBH6ZstAlIAAgs8sAYSPslDgVxGRh7yDdtGVKTtgs5QP9jbKHdsyEbS1jlnBb4GWnNj245dR/vpSzI34Ib0zZ5F/LC2orn4dIMlzW0a7MSM2ID//+cp49CdNLuIWUsH1gnDLXilYdnBXxz3xXZRtYtvKuvccq01S0Y8h+M8sU3BxnzDaCeIVnYsJQj7x9XYrzgOmSzRihim3P2jfea5RvPQX471Z7v0A8QZscjEd56WD8K3JJSrQwUk6cUlVxVkHjik6s0kE+oMAqLOHayPgq7xHRRX1gQ+XFcl0AWMyZfcGyXc2X+NO3D6o/9FVcwE+EznsX175P88X542o36WVB90yeQOeM79Utfwf2axYk6lwiu5O+MG/R12hV9mW8EJCXfNvKbq31d9Bh3JTPun+0lcC4JiJygHfPNMGKCPd8JlHSYy5sLU8bbNSWate8d32O+tyt6xpBsVzrt90uExrmy4X/3EvAS8BLwEvASuOwS8ITFZRepf6CXgJeAl8C1K4ERMJujYM2xNhYtBvpZnAEjL05ptF4ooCvwAvDsLUpoMJumLYslQCiAvr1u+w/vdVP3vsolOxqutjOUW6RFV5zoumjyUZfKNVQ8BZiN5rABeuSP7xYLM/LMMQsuc+1jpAKAEos1wAnAMhZnLNggPVjAmXY1e54DeA4YT3nNpQiV+AKXHKPfzVWT/c79LPLIiwFLgGPIEA1w+x3rAgD9NQuPOMlc0Ry4sqEy9RI39eCsu+NXX+P2/8sFd/QP75JLLK4b+mBXMqAfcgAwE4C1JRn/pUCW07nNIW+Xa0PWgMWUaY8SfwOGIl/Kxt/ULzJESxqtaeoBrXNAVLRYIV7MsgUZ4zoEcOt8ttPFmEAGTynRNtCO5W/eB0hJXqhzAF4Ab95L+2FPnbBxfqhxrnRdaxU+uW+h2jw34fK8itMkStI0dGmS3KRA2lIMr/Z3OoNlmVL0BMDO1eJ4nkDOeVHEcm+zIo1xeY9S/Isw7PSzolMUBbYXHZEViYBZ01a/LCDeiLSgn9CmiWsBaUGf+ZASpCF97R1KuFTCwoj3c60RS9QV9WsWUxedrxGhkIm4ID+AlRBatHGzMqONjJO4ADq0H7NUYAwbB5OHjQoXYhex8RxzNTau4c05LIUoM+/GmgNZGLj/YR0bEUCbN2sVCD2uY2NMQ17mQopxg35nFlsXkd3zv8UAYI1TjFGAZtQn4wUb4xrltfhBHIOY00cvyvUa1g4C3ZEnbYfvQlPteJ+Ihl1rHzvxdK7qy+fTjOJqhzKt6EVVVZffrTKsFHPFhYX8P3VLMRZZvyrE7Cn+S3WzLDOek1VcR8dHRqQF5TEC/PwFco4rz+Hy6WqMU/a9W78n5ybb4fHpiiJCw751q6pz6oDv/P+lhMsn2igWg8S6uBprT74bKC+w/a4SBAX9hXztU+L3oZUMdenJisvWjP2DLkECIg2Y65FKEQSMmae2kcUEf1v/5DojIoywNktfxlCICb4LzIXMio/vJvMz4s6gCIJiDLZTkHd8Z+gTNl/i/cPvLNYXvN9bYVxC5fpbvQS8BLwEvAQuSgJXXGPnonLlb/IS8BLwEvASuGoSGLmLMrNx3nsKjLtQomJ48xpY8S1KuE8BqEejEVCQhdAdLt22yU29JnWteyK39dsbLjspF0mVAlbXn3DTXzstawRIBUBM0xgD6ALsZ3EGWGha/iymcPNjFhdm/cA5Flvsb1XiOgvIbeAdADzXDBeHI2FbjIb1mq3IhgWgWV2M7+07yjPInxENgPeAhxbrges4hkwBTAPwgkBpyl3UNpf3um7l7w661Ufrrvv4E+7g+3V+AMjDMyk/AC/l5Jlo+fI3ANB/u1Jgy8jCArnhpgpZsShGCxrZUQeAPciXhTF1+xklAFEsK7ge0JfYFGiJIxfqh7JgdfOMEqTH2SwmkA/t4Gzb7+lHgDHaDItt8oh8LNA2PvQhrgCoyC95sLocEnIX08bPkaer+vO//++PxVOtWksxJ3Y1a+nmJA2/QT14vt3JvrK02ruzUYt25qXbpFDCaT/LpgcDNb0gPCHXT7lc9LfU2FdV13+veBX7B3mxrGPa1uPSKqcc9DfkN7hU9zdjLmWsz9AfaOO0ayPAIAWoJxK/jwMwRqyeVr6fv2Po99+2F2mInysGgAiMcasqjo28XD8enBawvUjC4lSGRy6ATrn+GQXVfpcueK8S7finlP6GNnuWBmaatsgOYMqs5Wy/IDlcdrD9fBr8OpdC42Mot5+PBcU5XyPCwsZZyBo2AmnfraDzbxTZMBxLxFzcJhuKCbmJqonQ2Cz3T5niW7TlEopxQUGTNOjK/EJEXiai4lCe5U8pd4/nZYllzUG5STuhvvACMPGcGbvGLxjJzSydxvtBWK/BaQZlEkWlxpMhyXuusWDkGsxcRfH9oD74Hj+kBIHBuM/YTXt9pxJjMecZB861kQeshvac4cL36fyvKPGN+kdKkH7UHXvywDeY71V/LN7Nud7pf/cSuGISGJEREGxm7WvzSeYtNj/lO8k8mLbL+A7hwNyaYwhtUwjg+8D8kz4HSU16j8ayXB2b0EgoldA3bGNuRgwXzv8/Sri8G8ZVUkLpxtzE0lcZ92w+zP2nvkXeAmNMov7QS8BLwEvAS+CySeBqaLlctsz6B3kJeAl4CXgJXH4JjADbNbf2Y9slALnfrceg/Q6QDUjE4ohFj+I3JE23+Zu7Ii3abvqh3a7oH3HpzpsVYPuES+YB8lkgoWUL2MbiCKANEBxiATCaRRsawrZQ4x1cz2KKBRqoJYs6i73BYo9nAFaQFwsYDejBfZQZ8Bzg3SwkTgdQAnJY0FUdvsASwywzzNJj3L88zza/7YCOgOnkcY8S4MwBgceJS5pTbvrhW1xjx5LLHtrhgmblnnvfFxQT1ggDvtfIkHs4ZnHKbwC+v0OGLuc2FmzbyoacyTflMa0+CALqiDyRH/YAQsgBUoKNuoM8oP6IV8FvbABIbD+uRBkgElgoU//UF5p/e0bXsKPsaN5DgLHAxlUQ2uM801x78AzaB/ez4OYe8ksZzLUWzzLg+7onKyjMa+/bVXx53/Feox6frNViRdTOn5PFxIwA2Mk4CZYHWbUjk+lEkVcyp1DDVQhhaZqn2g3yTBYVhRzjVJXcR5Ux9S5Ncv0+JKXoQ/SrYXsj+PZIdqeqRcDlWBWd96H1L3MZxI20G6sX3mmufU499FwugT4HhLm2Gfk6Pp5VIgCqs8UBWOfKySwf1hfqimm6j+dtRF6Y+zvAKNryG5XG+9AL8jYiZJCbgemQTdfMtq7+XmShcjkyOrKyYCyi7LQjtmW1LFn1yP2TC46r05+IwkpjbLBL50UMOxEW8gsl9kLERl/kxCCowkI371c07qerMHpOnhQfU4tUHIuSMccstS5Hlq+VZ9BXzJIvF/lZE2HZkqXWShxFkVzMJfq7bDVTxoSBxoLsbKTFiAjIRVzQr/le881gbEabG9dutGms4viNbwS/ERuGusMCjrb+JiW+148oYVHHdxUynLHfrGhu0TEkHt+Y71GCuMYVFc/me/SflRj7+f6Td7MeJf7JFevLeo/fvAQuRAKQerRHxm++t/QX2jjWrLRb/sY14cNK9AfaPXNWs2hljs38jPmlhq1A8XuCN2t/b6DAVa4qFDItcVGcuHzQk47M8FP+hPbMs5gvMWdnI7bYnypBVvBOlFCYQ9Fv+Nss5fbpmL7NXOyirR1H7/Q7LwEvAS8BLwEvgTNKwBMWvnF4CXgJeAl4CQwlcAkExSkJCqB4m/5A8wvyAcDAQBCCcH5Grp46rrZtq4u31l3jtik3OHbINfYuujACfGfh9J7R3hZDPIfFnPlkB5QGTGUzgsG00gD4AL8N3GdxBdDHIg6ywLTVDHjlOkB3fuMZFtODvHDMvQBU5MHcmnDMtZTL8sDetFJ5P/miLCz+0G4DnAdsMYsOyBgWoSwwKRubXGHFLZfuLV10fKfb8aN1l26qu5XPL7kTf7ni8pNcj696nkvekC2LxXuRucCXD46eczl35uaKxSsLYot3YlYplBmLlc8rmaUERBVufd6khKwoq8WOQIZY2uDWBuuJ1yshL9Pawz0PYBXl3LOuINTD+0e/IwvqlEU0VhzIZJ8S4JbFEQH4soDRlt8bwqJinVyGGvkKvp13u/mqAmqnWVEeFRDRy7PeTJX3M3mLkmZlGqaSUhhEXTm7qct1/3Je5EddUDQU54LINh1pkOPHf6CWLD5j2L4BTGhjRgCsf/UF/X0GwuF0wPXFAiCWTwN7bHywcjgLZPxSBzA+D8EZeUO/hqhlPGTcC5V3I/0oj4HyZ7U+OY/33TCXjJEWQ/cqatOJyDjGrxU5hsrES+yvoqiXxuFEIUZYvqCmZeGn75++QniKUh8QvVcEZXAiD4LDIimW1TUWxfmZe7KLbZ/XnIxHlhXkyyyKRE7ENYXt2CKrCoKTL/UHeUtu5NJGLVmRFdZx3GPNTNV7uncIVp4HcTF0vzeKaWLB6YkPw4YsaePUj1lBQi4AkuIuDpkz9kNsMAfAnZy5quH8HiWexfcALXHICe6lP/B9xRUU7yjORXiO8uN3XgJXVQKyrjC3eOaikrkihJ652rSYRQSzf536H3OqWxmwpGlwrxq6hq0Id3cNnblPAXhuDTERU5eO9NFPavps6NooSRSsp3DdxQXth7o6YjDUUcp8SGBoCKTb0A+Zg9sGQfgRJXPDypiKUsn7R/ljTm0x2zwBeFVbjn+Zl4CXgJfAxpCAJyw2Rj37UnoJeAl4CVxRCQiMADj+X5VY0KD1hUk6IBtgmwW6nnAv+9fbXPPOSCukRVlZ9F3zZQDMLNhYpAFWAzawcAN8BqAzCwUACf7mPYDk5kLGYhGYVhrlBKwGLAcAAfwgT387eiZAOdppACE8C6CdhRZ5AJg3cJvnAngDlJhmJs8E2OH5aIWi8cZmYCHPsI1zBvriBoN8oBnHs8i/ucpCLxxrEVaQuUiLL7po670ubJ1wW75TJXgwdLNv3uSe/52dbvFjFiiRdwDSIDviWgSSP+D/vxAoY/7rx7JySYcAosiCPe8jr8gNUoI626MEgIQFhmn7saClrpAXe2QMkEQdkj9AJ0gis8JgkYw8sYDZrUTdAjJBhFh8EeSH1uzfjd7DdbwXOVNvBlazgDaNXnMnxLNuSLJC5bKtVHDgbl4Eq2lcPDLIu4Miy9+QhP1bItedK6JWLpcu8u0SnBwMhMZWxYpiVRzs9wtknwmuEOgQQCadEMCLXGnjyP5UXIVzuYEZy8sVOzxNYGJ7F3VtWuIAPeSbv21coI2wDWOZ6DnD9nAdEBe05Q8o/YgSffwx5f3j5Ft7yvluJYDZT+hv+tALQKNzucG6YhX1Ej9YbbUYgfFDKyuIODWGhoC7IQgoAkIgvCA+WVfg7khmRz1dEwmYV4yL4IR+EffnVgUILsqw4DkJlXoAbM+vhX5wmcVrZHsqWWxK4iiMoyAIg/C4/pvtD7JZIaKz6k2ZrLLqklMuK6wTaRIvDLK8i+XVecpknJy0MZtzfPsYa5gvGAFnygZm6US/ZX7w56M2bm5qICT4PvE73x3KctFxUC6zXP3jvATORwJ8g2m/zJdQHGJ+9RpZ3m7X8d9Jm+BBjer8pu9zNRtE8avjtP5l7btFNni5+ukr41pd1su4sYtWwiimP8T5oO/SiUmX1Nf0ezTm6S2D4bk40eVRdJvud0XWF4GRu0KWF/w9vG6NvWCDOHm7Etavf63EvIu53uuUGA/JN65JD4p44ftjpMuLyu1dRp1PU/DXeAl4CXgJeAmsl4AnLHyb8BLwEvAS8BK4JAkILEfj6yeUAJwBHljtAGyzoAGohrQ45Pb83E0uWyVmReCmXv9RqXwBgLM4e6USQAXm6XyXACs+rcRKCxcPaHBBBqDlBeDN4g3Agvst8OC4Fri5lKFcAJMQBIDlLAwBMvcpAX6/VQmwjzzzHKwdeL9pMJM33s3vaP9DdLAog2yAUOGZkCIAJGb1YYCLAagA6IBkgPAEOgRUwaUFz+YZgPnk0YJnQ0BELp7ouPDW1HWfmnNBHLjN75lz+fKyW33EtK2RuZE2yIHzP6O6+HciLcjzJW1aKOPr2EgK5I2lCPI3CxfyCYjHOSN1IHAgFiCrLDg3cgNopb4oKwte8o71Ce0D2ZFf/Jmbmy8WwJQHUOu/KyH3fUqQV9ShOf+hTdAeDKSintjMx/PoT2nXSrXa/rgR99/5+lvKX//gE0Mf1nFYhjW3eCgKB08lwWBLEvae7xbtvBaUOyqFF24XDQG2taIKGkUYupMK2J0oXAWxK44rITv6rJF0FvPjWpbfuAsojhvSipehSdVVIPJJubIRvloV+iFSIVL93eVUPY0HAvmLa5G0gGgYkTPmzoxxhnHyx5Sw2KLfMFbRT7BqI2D5vxr1k1N1xTM2KmkhWdi4Sps4KaF8SUDczRoLtgiPE0GhMT0IWgLpD4mkeK7XzxMRFXXpKyNb+U2pntXI8qSsChjn6RO4QbphrCvGxsEhYS/3T00Fq2ilaZTNTrbo983Flc7tRRHek8RhX2PDpMDR2+Qu6rD+Ptyspz1ZZcmdVgU5VJyLtDiNhcMLxhR9u4ycIGvI2ay7+NuupS7smHo9E0F/LY9XN+InyJfpAiUggJ/5FXNDlDf6GoteFoROSgWRjqNvjOL0ZllLbBKJ8DaZfjXCKPk9kQlJGCd3pPVWu8wHDyW1xu36W9xDouFKXSYIJvU3lpSu1lL3CKM1TQ596CEiYllchOHU8O8obUhvSDZmShAWvZWTLkwyl/e78iBlVhdDXRxcrKJcwtyXvPItwmUb8zTmHIyNuGTDUurLw7Hz7HGWLlBS/nIvAS8BLwEvgY0sAU9YbOTa92X3EvAS8BK4RAmMyAp8R9viC5DBrCbQzgLYfsyFzZtd6+UNN3HPAde6FzCEYMxodENysGgD0Gbhw97850IcsN5iD8DPdQaam/a8mapTErN04DdzCwPwAagBIE7wZ/IDgfF1o/dBiACC8z3kWgB3AHVAq31KkAIW/wJyA1KFfNr15I8FHIs0c0dEPkxrFW00riWf5InFH+QGYL0FgTaXALyLZ6+5xwijo27+GwcuO77Ntb+4yy1/qufK/nOu8yXyQBnJD+8kIRvOfY/q5HcvB2mhZ1GX5BHNV4sPwruoD2REPeKPHFlxzfePfsPfOAtbyggxhK9lyCCAVSxcSJALWEtwzLWQFciG+sCyYp8SRMnDSsiTtsJvFsAdOZnbLmsD5McII/I0bA83OlmhMg63H3nbnYVIC2lPTiw1yqeOCrN/QrY3tWawsDd1S1NhlfWXs1ZY5VtOzsYHpnrVXFZUtUEt7MfiLFbLMigHrtEpqoR6Z0OGHJuVhb3qWtzT32gH8npRltKeb3V7g7yq0mCQFVFXauITjVR++V1DwGsmwNWttPtDV1EC9YfluxaJi7F6oH8zbnyrEpZsEIH0L/rAe0fXYW0BkIT10ylgfaOSFpALAtKpY+qXdnxUJIUR0oeIWSELih0KSJ/IkuAgftB0qlEV5YwOZV3gnhMGaIQ14yDA/Gnb/kXGcnlJ+9HIAsVIaYgvCPRt7c7gfrmIOVmvJ/quBTeLxLhDA2lfrF8m3neTCAu1LZziu82pTDEGedHevnmS7/YpV2UXU7DzjHEyTkR4UuJiBO3veckkMCIp6HPM8ZhD3SHDiJfFtWBR+2/Q+PNgGFVTcSPZ5cpQZILbGiXNlsgKV+TZD4T6oIlcdSIrXi5LCvEasUiImoiGVN0RL1D6XwPXcOqj4yGJoWFNxEcgcmOt3LbnOFozCoa0GE5YlQGOs37f9dsnh1YXxPcZWVx8ky6xWGC8ZJ8Sc1BctTF+8H1ifshYe0ljwUtWQf7FXgJeAl4CXgLXnAQ8YXHNVYnPkJeAl4CXwHUlAdwdARygRc9CBfCehRirI1ZDz4qs6LttPzhwM2/e4WpbzCc117DIQePefFRzPQA2ABMLHoBsng1wzd9cx0KPBIDHxnlzxWQAhrkwYg3GO9D6+iElvnlYOEAiYCUBIAtJYC6meI69iwDPlOVLo+fjgonfyB/AKPmmvAD1WA6wUON9BhQaYQHQb77PjVDBEgFtNYJF8xzM63k2i0AsMsgfz+HejykYecel2yfdrh/f4o78/oSrsiOu+zTyI39GknAvdfBflKgTAidejo26gIyhDBAG1IFZjVB+gFPKBTlFmZA3ebHg2/xtcT+oMwgOyk2Zrb74nfdASpDQ3IO0sgDp1IvFELF5i5FG5IFrqXNzA2Ry3nCAFqTFo3/9U7IucCekO5n1y8lOMzzWO5lt2dQITqRZvj1ul9XhTe4Lm2tRZ+r55NYn8sId75WTR2eT/YF0MGvSxQyToJMomEp2PN+T7R+86pza05ejoV3kM8y6IsryMh0Mcmmohk259tkqomLLoOilZVFG4i62Z1kVJHEgJdNY3rLKDhrjIrNWllZ67enJejGKb3FGDfqrbakwZmUBKERA4u9VYlz9BuX1N0b9B//itkH+MtZBHP6BkhFPFynaG+I2xgBzOcTxpOp9QlieLG8YN4au0CYFBO7QaITbqLYwu4PaP6O/D8p6AMKiLULiRpWlEfsTAjin5fo+FiB68yAv7yk7mbw+hV0lzO0SnS8VfxtS+R6xwHMiKqaqovpskkQHllf7/QtwDXVDNCxfCC+B9RIQIXE6ofCNYmPeyHyTeR1zwFTj0N2aNX5TnAb3NqaDHV3NagKFn9i8u5IFRJl3FqPmyoKGLQ1KsrhIg7QuPZa18GlxQ11WewiKMFwLNyZiYvibxjgUNfht3PL4jBXGfUmToVHuIMtCUWyakVgRV4gIGXTbchU11P8gmPcw3s/wZc69RekZJcZI5uTM6cgAc2fmi8zH/OYl4CXgJeAl4CVwSRLwhMUlic/f7CXgJeAlsHElIE1+zMTRmse9D6soADNAazStZl3zrsJNP/QJ17z1Hjf3Tc+7eI5vDgsZLB3YWLgBwEECADizKgL8hxzAigDAGjDbLBYA6Dk2LXoWYyyQbEFo19nvvAMwm8Uh53g/C0Y28kteAOMtUDagFNehLcpz36+EFjOEBhYCEAFmTUFeLa4G7+A+nsl5IxGMwDCf+kakIB+egyslXF8hByvv7Tpm8QcwRN5eobToajeXWiw+7bZ82x6XTH3CPf+7L3edpygPeQZkRcsNkuDblB5T3SxJY/XjOr7obeQWaujrf/Qeykh9mQwpH+QKpAQyRrP7cSUsLCCEKAPuoSgP13AfQc6xuoCM4ln8TX1zDvlwD6QIi2DIImTHvciCa8kPC2HqiPwYUcEC/UZ016Iint+mOl9zm5b/26gIJ+PlcE//6GDnYr1cWZwMo1lBHsdr8UI8GRxyE8HxlUaw3GklB9xqOB3Vg5Vb5uLn1NcqRe5c+qta2K4CedKqBZ2yHi7Xfu4vXkAKGaH4AkJovcsX5ce2Yf/U71eKQKIdpMo67n3k1qecEEFRW1rtJ/VUcGrs5gaDclqxR9WuROJkedqqJ8elWS8Cpzgq11Cxru9ob2PQtdaOyBdEH37EGQ++Uem3RWh0RVwQD4ZzH1Ua+kDX9ltKjA2QHEPQaCNYWZzB+oE2Z/FYzH1QV5ibXNxVjMPPC9d7Wi7R+HaxaUyujujvw2qt5rLuRtYWpm8qZkWo+OKBxvJgUhYUJxXkZpvAyxS8U2xFU/9PwQQSu1e/rUh+ZSJ/c/JFM61z7UY96bcVNsfa26me7w+8BDa2BPg2MS4zJ7T5LueY7+2JkvCfNvVlnt1RKbZEdEzeoOaSWtmttaq832nM5P1g6KIpTmRJoTAVsdw44fIJ0oA9FhSyfBruRU4wzg1xHVlJrMj6gvddyMYcSr6i4kwZDMJaLVT8niFBIuuOxR2ONgAAIABJREFUkb3q0E2obSjbMG4yxyNhgfHNSn+shPUsc8Flxa64Ut/9Cymbv9ZLwEvAS8BL4DqVgCcsrtOK89n2EvAS8BJ4KSUgMPJdej9ulW5RgqRggUJMiIGLZ55wjVv3utr2rpt6ZSw3UAcVaHtOCyGAQOI4WNwCAH4SCytAa75JLIC4ho3zaNID7lvwXJ5hQL25JwKIAgw3qwYWSGjkmwUCC0aAdbT3ed8eJYJwQ7iYOybAdsBxrjGi4Q06xiLjtUoWrwHLhQeVALMs/gQLRVvIkTfebW6x7Fm8ZxgMUckAX8qHixeL3UDZeI65t+G6tRgRUbLTJduOurJ7QKTFba6hteIz/+Kg6z7DQhHLB7SwgYghVaiT71QdbRZIzOLxUjbyQHkgFMgLMjL3NMjSrBkgKdgIjAoQSHlJkBUQD/tG5yF/kBuEgwVWp+6xqqDukQ/tg9+QBfWBSy7OWxBoIyq4zgiVG35RPEYAjER9KtA4soH8sfZVj8qVZLJ6suqGUadTTH9KoOL+yPVfW6tOTK+UM09OxEdXam610wjLKCtjxXYI21mVuqno6NZmcHK2Hq50QlfcIw4IAg1CzjQmIZJoE5CMkEinNuWvUHs7BfZDYOgceRv6qNAxv1l9QWBc8LbeymEsCLfA1KDWH+RTq91MVkhuqtPLtsjKoiavNfX+oKhLBpvkKqoni4uJYLZJUIvuoJdvkwupoF5LunpAopgXxLS41ggL5MQ4+B+U/tFInvT5Z8irZPCojnGxB3kx8vsxJFsZ//79qF1csKxvoBsYG4zoZAzh+JQVHmrF+pvz5i4KCzLa9tAdGgG8byBZnK4oCrEddElR6LbVkrhWROUmxYCZyzLRE65KJKGUGB/iLyqZXbRlwbQljuUlX3iqPLA9ouDbuWJa4DJrdQPI6wZvDr54FysBAkvLysKsGhhPmMdgidBX/8o01DBPxdr3rfLS5Ka2pW7r7YWb2ppVMmiYFTkQTcx2W/1Oz6WNXB6bYn04Q9fRVzfr5UodV5+cGVpSyPehyATFqDD74hFZQd4Vo4Jv9oVu5h5OX2zxFmGikFeDIG22hoRILvdQY8G4154dBCgK4GYVhRnWASgj4Zbwr5SwAmT+yVzZb14CXgJeAl4CXgIXJQHTSr2om/1NXgJeAl4CXgIbTwICHt+uUmNZAeB+rxJLJsDjSTfxip6bf0vNte4pXO32FTd5J8qZz8l+HY17rmMBx2IKF0LsDRjiewRwDVh0nxLguFlQAHqzAcaZFYWRE+YGiMWhgaFGavBs7mEP6A7IumeUD64HCAeIhVzgHkB3NPw5j3aYxZzYp2MWYuQD8AqNf0gGc1kEMDjuCoq8kk9AxnELEc6Tb7Pk4N2A/uSNcuDmCUAf6wOTDXnn2YD+s67oL7ve08+7zhOzcgs15/b9YsdlC5TFLBN4Hnn8ghIkxgcFDF+Se6hR8G0Ws5QTeSIvLCrMgoJzLFr5HQKFtoDWNyAgbQSC4nOj/HAvhAYgK/eNk1UmKyOHyD9WI2wGJhoxYUSJ1swbYyqzjrCg0MiSRFtkTzsygoA21ssUQ/hovrc8lN0jpxGDnXHQ2/657nsO3lH7sOovWJiKjuxthou3HMzu/ctWuFDcnH7uzc3w5PMiK74cBdnL5C0b2Vs94m4IogmwHFdg1CN/s1EfABPUlwXdtH5Insgf19CuyTvt3Yi74QMuhsAYuXEKpd09ITLipm4vu0WxKaZqSeja3ezlHREYjSRGIbxWlUGkDOUCYTvTrfRgHMdHpE/abTXS/brgQL0W59Iu78rSgjwS0+KaIi5UVvrRDyjRt6jff6w8DkmjkRwIyo0lxvhGv6TeNnLw7aE8RjEbGNON4GOsZEw3t0i0R9qoxRbqC3y/Yd2ajMWwaIiom5aVxS2yR7pf6bWKYXG/BFETaTHIs6opS6RMAT+critrkbyv6UdhmgMRGM9q/P24aI1PyUrpCfW/BcmM8d9vXgIbTgIjsoJxhbkR37ydmqC8VcZJO8QivFqmDw/Qj5jSzWyr3OZbU5c2FThneiB9nkQkROQ237Li+p2gvfx80l56Pt7CuaKfuKWjE4onMS0ri9aQqFAfLUVMjFs8rMm7qh7RnG1Ov8mK7OI3WWkM8l43yLN+VOSDMJNrqKzLJ35tCk6gbuJoDAN3V4pps/aDKcJiOcx35/eVPsSY6i0tLr4u/J1eAl4CXgIbWQLewmIj174vu5eAl4CXwAVKQKDpa3TLP1DCYgGAdC1GQ33XM27Lux9wm7+r5bpfVuzevaGLZz/rkq2YvgPwo5m9VwntfLSxWNwAdpIAPgHe0OYG7AAMRduexZhpw/IMgE60uAD2AewgNfiO4ZoJ0InnADBxzB4wyqwU2EOSsLDimTyL6wHHIRbMXH+fjlmVAcpiXcF7WXzyHs5DXEBmYA4PoI7GnGnw6vCUpQXH5BOwl41FrOWFfLNRBs7zDAN3eS95MoCX+wHQIHE+46JazU3cVXPpXMPly7GbvDdwJz5s1g+4jOE6yoULKywttqvOjgsM/uTonZeyIx8WoJyyG6mC7Hgf70WuyJM6MHda5A8glfOUD2KDOuYaiA8jvMzlk62KT5ESusZAsBvekuI8KggZQ/YgSyPp6ANG7PGI4fkk6FXz0b6+CIvuZ7vvWbopeWS/lKTr7XLeTUbHFmRJMTETHbptPt7/qqKK+rWgvRIHgzR0OfVpxAL9kLqnfqhr+hEkiQVkpy1Qp+SHhJWNWWSYFZTleY9+o70/M/ZM+n4wZoExFMH5EBgEysbKIlf8CrmvUSiCqq84FlUcJ7snGjFj1JY8RxZVXw5t5Ja72KzyDxTj49agLNpZv/pU4EKNKSXXLjXkwl/AqxNpQTDuay0QN2Mo8sTii779+8rjB4bCWhuDCFaPfP8XpX88Ov8Ptf+fla4p8mWUt6u6E5BeCaS38d+s2fiGmZXd0FG70vCaG91SAHlQVsmkjwWFLCWCNIhWi7xI81J2SArVK2y1KbcwqWBRuYwSPCln+XJCI93woCiLqiviYnecBCcV++JQLYkOykrpBETI6NlXtX6vtZeNCKHxbI2iIbvKy+daq61Lz88ooDbzROaMb1IaWp2q32xRTIiHoqT2CpEMOrH6bBgWu3e+vO9mb+rI5VPkahOVm5jryYohHiSNIJNLqJUgKJYPPtZoN2e7u2Zv6sVJo3InD8t4sJJphWwv1DvNSgyS4m/0IhRdbtH+FSMlDlPuuajCqbu3Nd38dOXyKYW1ui2op40gaEzk+j5CVpzyxIrCSFWtjaFBMNAx33PIcyylydMnlAaSTynSYsN/hy6qMvxNXgJeAl4CG1gCnrDYwJXvi+4l4CXgJXAhEhCgCBj5Y0pYFljw6add47Y9bv6b73dTr8lcf/+kSxVYu3XXomJWAKoBSKN1zTFAtGlisZgyF0OAl4DftykByAH0s7g3Y/dxtz+8m2dAfJirDoAmiAyex7UskiBCAHVZWY0HprZg4ACq3A8x8mElQFizsEDTn/vfpGSkAouwW5WMxMCSYM/od/Jumrs80yw7KAP5JE+AurwbgGwtauKaHM1lFPnhm2x7SAueC3AMUAzICyD9cqV9IoIOu83fus1NPbDDPflT8+7EXzyi88iYdz49eg4EAYvnH1Pd7RcADJB8wdsolgX3WewI8mwxOwCqKc+B0YORj1miYBUC4UJ9Wn3RFpCtxfXAmsVceNli9gWa9/p9KKMNaklh9WVmJOxpJxAGtFOICtoHMqP+kT19wVxrrYqUyD60/NPIODyS3ZnLoiJVkO1lBdXOH2j+wRda4fGuYlrMp2H7eOTyY8ImARvM2oW+A1BOPzBijf5KHWINRf8x8o92QL2SByyFLJ4LfcL6JmQllgLkl35Ce+Z5XMt1tFGeXajNjlvTnJbAGFkWEHC76vQGmYIky/VTIJKiujMrq939vGwKJJKrm2g1jqO6iI0ZXbqqJ/d7vXy6089uEvJ6cKrZqMvtBaYYx2WBsSTC4loEVhg7cLXBWPP9Su9WQnvVrACQF0Tgzyv9D0q0gZ8ZXcN9N7prIxXx7NsIKIa4oL2Ztdu4idaw3jcKoPxVK4tK3EQYy1JCjvFdTf1pRsrbPUlInmsCIaTSoFYHUd+pDWNbuEquoAJ5kNLVcTgnsuNmkYBP6j7GIiN+zlUdN+TvI5lam4qa9QSXW9VUSzywNrmfc3/8yf35RCOtji/SpV35XW+49Vocb27I+rnUQp0hsDZ1y3yO+dZdSu9QnT+qOBJv0P4dSb3p4lpDwavl6qke7d6kL3WtFcnTZy7XT2V/YrYMJjfncVVmURBVsTiAemMqn2/O5iurx1w7rlXxxFyeR0n1zMpCuiPrJ5tk2HBC/fCoSAJZbyheWVVt0vFaO6oqcYkVbt70DSBxqsIaiu/wnnPIwMjcA1EcL0fxRD+aKcVFRlUYd+5bOtKs5bL46K8uY+WhAUD/GCFkwqi/eb4p5PCa+5Sntw0JlbVv+wvcSF5qXfj7vQS8BLwEvARufAl4wuLGr2NfQi8BLwEvgcslAYK9AkgDXgJUbnJzbwld6+VzbvbNSwoCXXOzX7fswrqAjgmAagB6QHeAVBbwgJXj3x0AUABrLCsMxAZsteCdAB9odGPhwP3mrsP8tHMOYBTyANAT91S8j3sA9Ti297E3Swjyb+50AHwBaFlMAdKa9jgEgxEqAP8QCBABkCFYEnC9AYAAuhAL5BfQlvyZNqUBzKb9Tt4MzGBhaO5I1ixVvmpVwv1D1zRKmPbzNxprPB95LWgd+ogbHJt3u36ypcDm97nnfhUNa/LBtUYUIRdkTN29X+mitlFA61KLXkgnFp3mJsjikSAb01SmfMiH9yJrC5ANsEqZzAqGe80Ni8nS6vmUJQVgz0Vl+jq76SwxKig/sqWNYAlgwZVpw7RXZG/EkMmTNgsaNpTrz217EMAfbeqyU84USsP2+WfL/6T3QPP3PyNXUOFddUKgDK8H9KYN09ZpR9YP6UMQEjyXvgFZRf2y8V6eaYAl/QUAx9o9z6Lt0uYpB20aQou+zTMhsjjH77QdrHIsdgn964xAh9zQhPKhX1PDqYuUmE7TciKJQiE3QS8RgxFHcRdgRY23XlSVQNlicrU7qBTwVN6ipKgaBrHiiqo/hQd02yfjKCLPvM9kOSriS74zQoI6Qb7fofRvlIj/YhvXMIb+rNK/Gp2E1LiXAN1YpLzkpbgGMmDExTWQlWshC9KMDrsym0j1ZRJGGYh3CDqyeVK/l21F4OTMnn5e1WVVIWxSVEUYCIRXzJowzELZNclh1A59G3bpHuYHfY0zG9KKYMztWKRYHzJIcank1JQrrVAyjEXqJGHdFXJhxzexm6ZRMRiUpQiM7ObtM2cdb9bH77kWGs5Gy8NpyApT3uBbzNzr1Uq7NGf5vjBOXdKQG6eh66REhEVT5ERTREXsGjMLbuXYfBXF7fb0ts5SfbKYln2grAS/KlHCXzemyiypuadEWOT1pUCEelFMzC0eO/5seKK9OME8lLFe36vgXeqnuP9bewLERFnJcqo8qYDZfGdlHpWoT0cExj7XNtQNCaPiLkWz2aw+faQ1XyrkU9Gpt7IPNqeTNx4/UJuJ4nnXW1kaxrbghqoa531PvSLR2Z/VBcTv+CPJj3mMKSCduojYH37zEvAS8BLwEvASOJ0EPGHh24WXgJeAl4CXwDklIDD1J3XRw0qAkACYK27bd7Xd1u+b0TomcVErc9Ov3aJF08dcfc8OuS6CnCBuAa6TzK8+9wG2AQZCVgBeA2KyyAKEBXQ1ywreAzjOeVvkcD9gohERZiWBtjnPZAGHFQT3AYICCgDQWUBiAFY2A05ZYVksCu4xDXGuARjmmbyP5wLkYkVgbqZMu53zgMaAqtxvZWVRZuA7e8rAotaWpEONdyXTrKRM9jt54TmQQuPEgFlmcN3DWs4uuqnXHnWDAydVB3tcd3/pjv8ZMsLaAmsYZABZxEL2HtXhtEDrX6ZwF7uNrC1Mo9tcP41bwJBvQGy079nzmwXHtvJyfj1wWo25MbjY7N0I941brxjJxh4wnz5FmwfkR/aAFbRf+hTyhrxjD6HwIlAA4Yy5gRnXJB/W5zrChDrCxdg+JdoR+TKXZrRl2iVt3wg3+gbapfxN3izQJnVPvbPnOcSpgdSgf0MK0lbpnxAg9C2eA6GB6zWLeUO5DhDUmzxAvJBf29RuArSV5We/LndOdbmrSaT+jZaq8hFMKRD3NllNTEpFtJ9leSuMwlT++uUwHKXTqiF0tiXS48moESy0e64QtphPSyl69P5rTfMZQBiC4kdG5f+n2v+DkXxNJMjnPyn9tBLjABvExruUhirdfvMSGJOAvD6VWRVGPewlBKzLFCBoy7RCXESgQC7yLCcAVP0HXWqhr8S3V0xeuaQRCZhkWRmLF5QPqTLVvfRxc8m4oYQ8RlaIBw01plVpLUm2SI6Mi0WchF2nsWalk01oADoeVHlboHS/UY9XGrWEcX318LGV4h2v2rnhLaGuk4Yz/q3GivSNSt+jb84b1wiKhuJN1GSFoLjUw+mOeMGoJux+xg3ayXKRp8cbM1m9Nd9xUapva6VvO11s7TvJ1lUHXFD7+T3F2L69MV0mjSV3tLMY72pM9xf6ndrb5EKKecEmERP0Xe5X5wyZrxJ4e6LIBsfEVOxVzAvNGYLzCsStvi1jirIXaiSQrkg3Tou4OT2I5VDx+Yn58HOiTdLaxPLXnDwUzx5/tj4MyO1EVlSDrgsTlRXlgKHLqOGGRdYdeuL7QsXo0MDxAeVp2cezuE5auM+ml4CXgJfANSABT1hcA5Xgs+Al4CXgJXAtS0BA4VuVv4eUANAB5ve7ze/a7bZ+782uLsXp/PgJF81PuWQmc7Wdfa3KADNNix7NanP/ZID1eLBeQHiIARbsLNTQHMY1E8f8ZhrctjgEDOHYEoH9IA/MGsKc6wI0ci8WBvxmmtxjOmwvcDlDPiE0LI88B0DViJSDozxizWFAKtfgxgptcOJzmNsbyjtu0WFkxdqq1aIWfpXQ4JxpdbMHwLV4HGYJYs+z+/m75aL6wNVvK13/yEm3+TvvUiDuR13nSZMZ4CSa65SNuntIdfmYAN+hKv3FbiPSgneYVj2PMosSjs2SxUgJU70bdwd26vUbxdWTFfg0lhT8ZO3ZXCqZtq0FdAcQoQ0D9kMIQF6YNQJ1AdBP37G6P2v1ns7lzbqYEdQdzyLRDyA0rB4NzCevRkZxHSSFuXHjFurb4pxAXtKujVCBEKTvYOHEOayceBbX0wdwG8XGOfoVBCfvW1U+kAFxWYbtDwsJaXzXu70iEIAqrDBIO/18Vtrgc3Jxkw6KfEIYSmNiIlmWn/26IB1xFuFgtTPoiNhYjeUCp9fPZ2SJ8bxePCPCYkXkR0eoI3Esimss+DYy/TWlb1X6WiU0eiGFv4IGNvE8Rhv9Hm3az4z+Zgz/cf3+S7rOA6ImpQ2+H8X1gCzOZDmxqDi+/VoaLwkknVIsi6YCV8TS1BboqHi/IeM69m76Q/6jdG2qwyLLginFsejoWIHtK76XfCuNrL/hJCxi4nRlsvmJzLXCumQ4J+B3TmDtZuG528XslCJOO1EUbi2ycnuUxs/mVdXpd7JOu5vtn591J0SalnIfNfi9jz49eNmeTYw73hrq2m091DfzU77PfK/eoURsoTfo4yLnauo2eSbgPhVp0RhaWkQC80UcVPkgCgbdstWcIX6FPk9Zshq4wbLojLZgf6xn+a6TGmHstqZx9S06XpAFRm9mR3tPe2kyWzw8tTuMKlxPjbagX+b9ZbmgSvR966mXDt1y6s+b1GW5hm8l52hTpzWFGF4WVMthJDOgWv4RXTURp/n8/K6T/eZMN2qfbDbFT96iyz43d3Nv75bb+6vPfjqZXtgfTXWXZdBRMEAodJ3CrGF1QflPbVU1K0rz3wRRUojI+UOdP695yrVb/T5nXgJeAl4CXgJXSwKesLhakvbv8RLwEvASuA4lIHDwHmUbV0SPKmGxcJ+bvP8uN/O6gesdwnA8dQ0ZNVR5T+TF3+t3tL73jYqK9jcEB4s6QEcDsol/AYDO3wZImlYZ1gpoJHLeXD+Z9QSPNcsF3oPrGBY+kB38jUso7gOsAzwF9Afw/xul1ykBkK4HAWzhCSBMXi3mBOe534IZ79ExBAAyYKHKuwFdeTfl5HqAGsBDWxAC4vOdNTBah6fyb36C+Y1jQET2gM4cm+soi7/BvfZcs7TgXEuqdMtu5g2SkeoCi5dnfh7tdPMlDFkBgUTdQN48oDo9LLD3MW6+2G1EMtjC+qyPEWjD72ZBcbGvvFHvo05pI5b26Jg2Rp3Rb16hRBu3tglwD0FmcVtAqKkH2uYYQnBFxGV9x/qxBZQffxlt3tr0uIszc39GOc1tGlYW9G1zH3W/jumHEDL0PY6H7iyUsBKiTdMfcH22qHYc7Vv5o/xI7Z2FgNKVWhoOyiqayOU1Q7YUhXLR0Z0D9aZmTPjgomqEaSSF0LKXDXJxFaXyUm0WOCuyQhSGqBZpPE/U0qimvyCAGFOuRWCFse19ShAWdygBaGFBMT62cfwFpX+u9L+NKuj/1B7fGxA+fvMSGEqA4OIE3hbRx3fzWXWdJ+UpbVLkXxZUwfSIIc/UxyAu5B5K0bmDQNrfAkld2ZP2eFLJu7186rfU3yY1GtFHz0ub+wargkAu6ZqJYnoo7ZD8Xja0WJF1o5TWZ6IgPikZTmiwmpELu5Y+iIq5U+wTyHtCMXcgW5N6LV6Yn2kuL630gmuQLL3BquvCi4ProlFwbcB/LBuZH2MByPzyB2Xd4NKmdHeGrqD0CZJPMMiLOK3nItX1HRPtoAbRWWyEso4Q0e5OyoKhEEmQps1sIW0OmEvyLee7x3yWsZ6+dFQfVd55R63Z396ab+8Sy+GyfiyLBkwigpqCes8T4XvNbacsoWRpqL/pvnyn/0rptO6gdAe5+nxtol+rNbO2nvd80hg8VpsY3COXUJNJmiVxPdsma4+kMdXft23v8svlIEqWH0VaawUL+Z+n96WNiVCxLVy/3XVFPlib8KpwQ+uL0aZxY0vpsu9Pkubfvu7tP3H4b//033ni/MKboL/DS8BLwEtgw0nAExYbrsp9gb0EvAS8BC5IAoCIAKeQB7e5eHrFTX/tZtd4mYJrb5V36znZvk8KGJwG2AdYBGgEqARs3DdaLL1Fe0BYwD9zYWOaXhagz1zYmGYmzwHM5HfezXkjNyxOBdYVbCzkXqOEFhl+73k/izTyZMF8KcO4hri9f1zjDA12I1F4FsncGrEHNAUghqhgUWlWESy8AF3NX7+Bs+MWFfae9ZqnnLfYDxzzLL7NlJFyG0Fje8pr5QAYAvwF+G27iQdrrr5LeRwcc8/8AoQKZUaGgN2QNQDByIY6vSTCgkyc77ZRYlCcSx6nsaygv1CHuHWAoILI49jqHXKCY9oc7pmoU9oYbc2CWtNGh31nnYXEubJzwb+f5vmnc5d0RhdKKr+5B6MvESeDtgjBR3uHhLhFycg4yDVcHz2tRPumzyEva9OMC1t3Pf+TR2u1D0otdG+yUHt7Kg8Zspqo+r1BEQoAlDK4Uonap9xhBK4vECkSVZF3ev0pATMNgYa9Ki+PD1zeFmCrC5NlaY8/r3vbcotjgZkvWFYXc8OYdcTpbj+lFYvFh679gC76DaX3Kr1H6TeVTq6zsiD/v69khAXP/RXd+326biMCyhdTLRvlHhF41ar6QE+dZlGjyTGFYMDN2kAAa6SvohzVhzJfEhIqAyUhkQMFsu8Ah2Zyv6Zo3LNlFTyjP2lX15obtatRh4FcO0FONEXktERcTCnUx55GPe3IYitZ7Q1mhFvXRaM2B1m5WXYp9bQWI/NccSxWRGR0F1d7wVSz9tzURO1pkUZdxblYVV8deEuLq1F95/eOEVmBUgvfIcjitythDfhOLBlweyRywiV1WVTIHdQQtC/L5bUYYIHFnhrGexh0kubJgzO78378zMRs53m1nekozY9G8TBwNWO3zWP13QqXiyyK+u308KCT7tDxoCqGZMRQ0UfWC6t6z0Dvl2VPwLxheHqUmGMwPx5XdBkaXgzJiqBa1X6f/uyIMKnNbFteTBrZk93leihLi7q+k3G/XZPlRHZQJAsxWXamjfyQvqcLrfnq1lseHPxVv13sOfD3zduXn5dvqzx2WVcOpPJS5IWsTIaWJqdcRD0smXyb7v11ybLtXUOdX7vzV3kJeAl4CWxkCXjCYiPXvi+7l4CXgJfAWSQggBETd7S87lRC27jhZt6oEJJ3Kjzn1p7cEU27wZHDLplfdHETkILFE4A7YOp/VAJofb3S25QgKgDm+d0sDkwjeNwCgWNbcI27QSKn5nIJMgPNM0B4iANA3Y8o4VYGEgPgk7wAhj6u9M2jc+utK6z0RiaYxhcLO/JusRY4xvKD/OMT3rTi2fM35AjPsFXZeMBtc0Fl54x4GD9v+WCBShmRH4QPhAsxOcyVEmW2OByWZ3NP1XJJuuwCiXnbD9/sjv7XgWt/EVKC+uN+7uOZyCymbgVAf8Je7PdXTQLW1mmzgPC0H6yNcPH0aSXaM20DN0nUN2ADRAbJ3CWRWYio6woYHCM8aI+4dqIMlBcgh7LSh43M4DxEBUCLuYSC1EELHDCH/nhrVJxsbe7/WSdNjt4s5e/NC8XDzaw/P6dotwORFpJx0JUP/hNywp/IT3ycZVkSVINcjjmqMJFiOMiR/H9nCimqwBdNKaXKHb9ojBePUVetgax70SmiQueHbUcgJvXOmPN+pftG7eUOnf8kZMZ4cF6dY/zDXcl/GMns27R/n85/5BpzdfVSyde/d0wCavsdBYZeUUv7SlEW9RFxVyVJWMg5flvuZmAo5gW0Cy2VSyhcs4ks13UDWVosityw+DkBMR1O53ruehe4yvSiIlDWbi8P5qYbSRJF8i4XtAYB8w/nrVorAAAgAElEQVSBz0E4LRltFYGB4oAicQeplOKbIimCJIpfHkjzXOTEkTQJkd+UjkWuBgflHorxPqe/e9LipW81I7KCuSdzKL7XEBWvUlKDkJWDeLwoUWikMh9aVkBWaGsXWf/JoRPCKJS7p4Bv2HDj05P1Yrd4eHpw9KlNvzq9ffm7RUQksp7I5e4pE5HwqIgEWeUEg85SY/fSkcltqwutXERH2j7RbPRWFT9CDYlNz2/x/q8+GwsL1xF5wTzD5p4Wc2p4mbwziYTInciS47KuqOqT/cNzuH+a7j6g9z145MnNx5J63p+Y6+yJw2K1u1qfF9/fmN2+VOre3cpfXfzM7Jbbi74IkwNzN+cLz36m9tp+u+FWT6ROgcFFVpyKc2X5rCmGxT1lv/gancBNJMoXfvMS8BLwEvAS8BI4owQ8YeEbh5eAl4CXgJfAiyQgMJGFzrcrAaayyFoLgr3jR1/m6ttbbnByRfigqIL5rouGimPmLumzOsacnVgPgI3/bHT/enLCgLhxSwdbUI27SzKLBLPAGI8NYcGAuQ+wn2ehoW7ECODn14/yZv57razj5IWByEYicB/PNjc9WF7wDogUA4optFljWKBtC5ptmm28y8qyvvwsKLnPysW7KQNWEBybdQfkBc8l/7wfsBZCZfx55v5qSlEPV11604S7+z/d7h5594rrHzILE67BPzLlQEbfrjr+e4HIvNNvl1ECZ4lRQZ3RryCPINVwKYHlkQWgp50BztOXsCygHfMbQBfHFtD8vFxxXcYiXalHmUUUZCgbAbmRkREU9DWLk2KyQ260X+LcII+9UbksP1BfmpL1REMERFElr1mox9ueWe3Gt/bkVzsTaCJAdUoxK1p5npVRUDTqSZbHSSXH/RE6pkUYxicExh7UheovFX2ffmhE4ZUq/wue+yd/86VTxO3e3fNOrmGGLuXkJqZSUPHx2DtW/4y1/7cS7kgYs8bJjeGzR9YYf6tDwCFIHrZfVGJcPJ1Lr6tSVv+Sa04CtClZU1RHZGFUrxT8RY2pKTc2wtnL+agKckGyrSLL60NCQ9fIkknn3BEsM/T3IXXQA7qfsetF7fCaK+1lztD0ZD2UoGAr5FIunlH8HGmm50F3UO2WfHA9V+9nlcb3MtM1fHNbEvh0LO32flEKtnbtJIkP445ukAWTdTmlw82PrrN5wJmULS5zSfzjREycTgi0aeoDokIKMMHbxWo/JKZAxMLQJZML4lRWFQ25hJockhfaVkVaHJJ7qJZ+1fwrwM0gLjpN6WT4HrlX2nnw8W13HD8w+0zayGZ23nP40aSePSMLh81xUnwmnRh0Dz+x9YdkXbGls9icVAwMtS2RASLZz7QpO/qOBaYAw3zRXI4aq5HpHaXIiai1abUn0mJm7qbFbTq3jdgrfIXndi3e21up7Zb7qpbcQc30OjXIDeajR2Xx0YrCYugSNYpcraicLEOqcHJTVp/Zkd0221UbbibuuUdrkdw0KjRGuUbgKAK5YuP8qNga5qK/KVn/N+QkSwvvHsp3PS8BLwEvAS+B00rAExa+YXgJeAl4CXgJnE4CBHUlkDTAPEDiTW77P9wp90/SGKwFrnV34aoic8mOWJEE/1q/s3rC3z6uXDj+EyULnD0O2o9bUxhZMW51YO6UyNO4RpgF27a8AvxyjgUU8TV4l1lC8AzcN7HYN/dR9i4jQNav9gwQwO0OCz3AY0B+yBqAUxLfTN5ppvVowSMfCz7MgnbcddOZykIZXmCePyoU+UXLHHASUBaSCCsLjtHsQxsNjfz1ZSGva/kLY+Wn6Ljm3gl3169F7vPfxLXmcoryPDeSDUA4dfzbo3f73ZWRgFnj0EYAlbFyoU1RJ1gd0WYA7AHpcTHBMaAI7RaAA4sC2rVZ79wwwNXI4uKUZdIY0UNbpvzIgvaKvCAoAEiQGeQdLqW4RgRG2U3KxWLSPZEV+eRsUOXTU+GmE0fjO9Pn+9MTWZbOhS6Ku8OAwUWsQKZhkiarCo4b5VVdsq16LqyEy1ZJV9rN8uFyWDEtlhXW4rISFmcI1kurG45FIigiaVcnCgAOFBWudAbyKCN9bPEptVQBN+BWvhrvBhnx9wdHbQgiBxlBtKzfICZ+QekblWhnaLd+jzS3f81rbp9GWhvzlJHvS+oHXxZo2RFkviqN/0XphreKvNpRBMXdukgRLKplERP69lX6TlYLumYYT0fnTJN76KbuRrSuOFPT2DI/EXS6KMW7VC7ndhASR/11Ffd0ZVHWWo00F2na7/alox66nkihSHIUECxLs6xaESA81esPpgd5qpghQzkSomBfnpdNmWTgAi7zffUl65iMz4yb7DN9RrBreAj3T3L9lISRAmwrXgW/xklNlgu1w2GUNPS1WZalhcVd4jvPt8titY0XpiUC4Lu7S/WvKFUrCxNc84CsLO5QbIt6EJYH1B+jQTdJdd2crCpO94zR80QYVppnrJFdzBnNTSlECdtw/qCGmivqDPPZfbLqONia68R67o7usuwQa5kcPxU3T25andJ1rYVn51bktkpuy8Ll/mr6KQX87k1tXbm7Hpdb9bv8XrkoStwrmzNVe8fdxUDenw7027Ibytz88tFw+4mDqZYKxLMY6fFop0Ost59V+qTS4ZF7KE9avGRN3L/YS8BLwEvg2pWAJyyu3brxOfMS8BLwEnhJJCDgkEUWWru4FEIT6hWusSdwW75lh1ZmpYsmFUlQ66FodllkBb71ccUEQfGnSrgfeacS5vIs8MY1gw1sXW9BMVxDKdl5Fi7cZ/fab1xnYD2/AdoBZrKAs+DX40F/eR6gJgCwPWM8T+PWHZxHkx1QHy1RtOAA9VnwQS7wDMsPADLnbDFoFg+mvTZelvUuoE5XFiNRkBmy/IwSIKMBt3yrIYKIPUFAcvNxbN9w8kUeeM5AdSJfARMH3OQrdrlN37TgFv7EghxzH6QSYC8WMK9TXf+BgONrMbCwsnd9bessK4yYM2sK2ih9BdAC8MAsZvid3wD5LBYK7Q/XZrQzwMCh66crHaPipZb2uvJVI3nSfyFtIOtot8gVkhDCEnk1RELISELHYVoLonSyFqzslKf9cCZsVJ10z82B7BOqsF5kZagYt9lKPSm7Gr9WquxkloSV3KgFvbysZ3ESdqQd3ZfP+UBEwVDmlxMkPJMrGco03apHnV7WTJOoKc9VoYDOej2UN3xXyYtVEa+0+1USKzKr/M0IDO0pi4w1ZpX1KR1DbiKTFxEWlEGAJ+7G3qXEGM2GiyiOIcX8tsElALkgQs0sFfGVdlKg+oTa36ziQfPdKAQySmNcPU3BuNVnGJsgFA+rQ8od1LB/8s3CYmzDAY+popTjIEtBKdCtr81NNWdXOv22YleIIQ27YSQtjyoM6zXRj0Uxq8FoUrfUJdtMIt2eySRjaTVbaTWzo5It5E8m6Fiob6VA3uNTqA3eUF+a4jPP2qqENcUDqp+3EqOi1prWVCtROJL+0BUUeHyUplkUp5NhFLV0gj5hVsBrLlXX5mmQCeu3E3IRhVXlgyIQHtI+ljrQjHrbW0fX63lDV1Tn2GTGIO+Guoj5hcVfswZk8wvyslNGD5XcUIUiQSLFphDRoEl9FWzF5RTEiAiSTERFUzEzMv2u+UgVyH3VNygwd29y8+qhtXjew/koB2rZKlyjWopy97hiWHykfTxoN2ay/6M6UG0vCQzO0MGlw9tEdKzNRVHgYM4diLTwlhbnql7/u5eAl4CXwAaUgCcsNmCl+yJ7CXgJeAmcQwK/pN/R5Cd+AguSBbfp3btcNDHQIix2nScPu6nXfkmrNX4HQGShhbUBgBhWGWj8j4P39rpxAmKkbjVcvti3aNziYjwQ9Xrig+etgfNr5AJxGiwIMcCdPRughQWR/W2uooxE4LzF1CBvAKP7lCBBDilh2WBum3in5Y/fTdsZQJWys0gEXGZha5qm5BEg2giNcbLFymAkjhEmaJFDWoy7guId9yixyBv6/x/lEXDIXF1Z3IO1BXKUSK1tS+7m3hyJsCAPlI1rkRf1Rhk4pq5/gsz47bJKgDqnLdAf2BODgvZnQDPAssVvoO6w7AHgYA+gYC7OLmumrqeHjREY1k+HQKiIDNoy/ZL+DUg6qbgUSVKeCJPs0IJLb15sBCs7yqTfnKm1lmp9dySIi0ZPIUnzPI+i7ESjk802XDix0qjFS64crOZV//mk3vpyEoZLcoMzEEFQTk7UrpY1S9jtK/ZuEk6WpZuRtvWEgh3Paqwtl9sZsQGmJ119s/iLk9LeJtjpioxDaF8QmmxoqkLmLIuYCE5HsoxcQ+EWanz7Tl3/b/XbhgOYr6d+cLXyuo60qAksHwiExMKJ7wwEBd85+kTdlXKbpqC7AtYP6nOTaX90dN2GDObebCSuniap4n40l1cHrW4/u32QFS3FqWhlZZ52e1VLRGMqonEgnQ9ZqYqILBWfOMtiWa80IpGl9aBsyXzlYOXC5U6eTw4GRRNLl/4g1wBQN6WGq9UcNuR7TuMOim8z8y5iBR2Tq6cfjOvNNzWm5ofBtQP5Q0rqTZf35Rk1qRWadmWyvFiLwRYEWL3xHec7z3cfhQWsKCEumJeOb9QvpDKkhLkjnVJvYx7OfI95+PlszPXoqzyDvA9dvY3ej6U0c/OviBzJsl66SaTE6vTWlafk+ok5ymtFurSIrdE+2XRpPTsw6CV1XTNfDKLXiayRNUm1EETlV9KmWu/aHJxvMGWjTItqr4dkcFLVWlVvz4P5TbK0eKwcuIMHvxg/UGQv+JySN+J/EEftfUp/rvQRyZ/v+Yu+R3IZdT5l99d4CXgJeAl4CdyAEvCExQ1Yqb5IXgJeAl4CFysBgYG7dS8ABYuczyu92s1KyWvyVfPSYD7h8uWGi2cXRF6wGPvCaHEB+P2DowXMq7Vf7xrJFtvs2Sxug5EVtqAyQmP9t2l8pcO9AHUCSoagO1YRL1diwWUBPwGDWbBhEs8xe57BYs5cSxmJQX54L2Axz9ujBPFAHiy2AMfknYUUvwH8kwcWaRxTXkBUFqHseZ/FHDhbWXi35cM08rHkYHFK7BDKRjnRtsfFFYtNIygoF/kzmVFnlk/yNidHys+5+W+ecbN/vN+d/AjBdx9WYtEMqIQVx91Kbepc4DCgp98ujwSoE+oK66S7lGgfJAAD2gZWFoAKnKPe0HLHmsmCUG94suJs1aC2Sp/J1G7pi2wrYdWrFUHSnCienC7yVn8lfNnB1aLWDeKlxXrVW86KTXuzPGhkg3KyVS1OzEadTtpoHperfmmOV0eLoLaw2ps6JjrjRF6WbblzKa40YSGN9qEVmaw6UsWpiGU9MStQ6NZMbmCkqa3YxmUk4mJOf2+rp7nMK6Kn+6Xr6G854qhkiBG1ZYNB+2EsYGwjEZT7TEQLRNj3Kv3OSG7/RHtiYPg4Npen398IT6Ht8D3meygigjZVYdEEkd7EU78u2Kw+s0PHS/pd37uKNsh3D2B1aBG2kdxBUemKMeNEKLpuL1vuD8rjGFyob2oYEYRbuob8ZzYJSiFCUgGVgxWZqPbUt1P14Uoen+T2KXLNujTzw6iRpuGsyI5pXd+XlUUmgyvqpIdbKO1f1LdFON4I7e6aKMM4MD4Ksg0xzLi6VwTET4uUeLg+OSvPm8kwEatCYZMUvLr+6TBObxMpJeujNbdP6htmTWtWks/oNFa0zGGZO1KX9DNiWTHfQ5Fkn9KdSswlUb7hWrPyPZeMmJ/yLWDeznP3KJkbUN7LOeYjWEGHioXhjj0zv33lWOtOWVJE09uWZWkRObmFciIoZEHSP9hbre3KutJ9qYb5OBFl0TONqd7norigjDQ8vh3MdZnXcG4adZnaRPWutFEtF1nw7H3fkn2q1w5+4+hT0Y/pd5SL1m8/Psoz44iRLFdLWeBcMvW/ewl4CXgJeAm8xBLwhMVLXAH+9V4CXgJeAteYBL5H+QEIx21NexgToX7zNnkmEcgdzLjGrVrJ3CIlwAiXQixQAGYBM1hgnU5rbDx+hWlOmbsnCx5r1hiIwhYq6/dGdpj7IxZxAPos7iwwLwAwYDwLPbPKMKsGIwRYFJlmGN9AFngANGiPkj+ewe+UyVwl8XwjBygzwJ8tJo1A4Xe0w4yAYM9ibjzYt/027uPB8kXZISrIPwtckxGafWjlISO0WCGU2FgsDk3pR++wgODkmUX2qtz2z7v6nsxt+/4tbukTd6JJrvNo/PN8nkMdAzRR5wTi9dulScBinLAHkEDrHXKCYMfUJ6QaMqefoJlI+0WD+YtKtD8L6H5pudggd6+zwOhVf7HSX5l861J/kB7Ow9mkm080a2F7cxIvL/ai1snVQSRQpbdptrY0v9l9djYuA5mMtcTYzRe9vPb8crj1hIunloQyZu941c6rZXWQEFxXoGRDI8dWaWjfIzB4UgF6g6Xl7vEgCuervNwhLetFERU7BYDOEoBb1ysGR0T7In4Pbc2C8/bOAmDmAj0/NOrzjDWMcW9T+qMN0mR8Mc8hgTErC75rfC/YGKsYm+YVh4HvEN+MRbVTvp1cxx4w1BQdrlbfuSbqE6smMiIrqZ7cPy1Lw/yw/LodqIKgvbJSbatENeo4k2unUO7d1IXDPJE7KAgOxbPIulkRxnFQNmrRCVlTZSIquhP12kDK+6UA8LrGI+S/IS1XXuIKtrkmc9wHlR7GqiJWYG0RFPL9Zb661CWi5E4XlMtpq/+JOK0ellul+bw/NKztyWKBeSFtxGJYoFjDPA13kJAVbMwJmBswnqMMRJ1b3CrmmuezkV8UXlCUYA7Ce5hjkBHmh5Th1NxTMSvcoF2TdUgsp1BlpqDfhY6n5JJq+K7OUgMlFqx9mbf+qVxA1UVU5HIXxXOZ11Imc0EIqQlpASGCAkYh51T9KK32TW+twtf9YL/zZ7/U+PnucvBfX0y5DV/39Up/pcTclGcy9pwiLbB88VYW59ME/DVeAl4CXgI3ngQ8YXHj1akvkZeAl4CXwEVJQBrLaPEDqhrJsMfVFLti09u3uHSrAtMmDSlYPqrFmVkTAMSysVBhwWIaZQa2s+AwjamhT3ht5uqJY7O84BoWKhaHYVy7CvBj/FtlJu6AvK9RYuHH/YB2ZmUwbrVA3iyWBe9g4c9ikHcZ4ELgP4gKFqYErsUs36xEzDrDysIzjKxgQUneWGyadry5XiJP3GvlshgFp/NfPE7qmAsC7iM/5Jd3Uy/8zeKXsrKxCKX8vJvr+RsZQKpQxlJ1lrvJrzniZr5uhzvxQaw1ACpxN7VHyepmK3UvABgLAL+dpwTWxawwF1CAwNQn7YJ6w8UTrsVoxyzyWYjjQo1FP3tcjw0tg270GBXnKdaLvmzN8uIPkXMh64X+q+7e0ZcdQjfvfXlF1mFfroW9iTBt3zQdHry1me27OyyymSSYfDyLJz60NftQZzW5d3U5n+i/46HdNlZddF4u4Maa3Dxt6g6CutxR1QRWhgK4tsq/+E71zuNyvUMwjc39QXFzGJYLzUYqC4tidbXjHs8Ld7yWRrmSueVgbM0EoBZnib0BgPXPlX55lMc/1PU1Xe/j2FxApd3Il45IC4rIt4dvNNZgbLQRAylNEYD+ZiQ7+xvaukJ95UxVXxH7RtE+0igIT7R7g2eyQuROEBxVEOJC7p1qInjSwIUKqu1a/aKUEUagUDWCudWRszKKe3mxVX9mIj4en27VBtLh74nMXNGMie/72fr0jdwcX5KyCSCnnTOnBbB/nerxuyGYxCzhAqpSMO1xpRNZWgQteYT6ytTmzgncLNWag7nFI1MEbWjpP9Wj62tkPyqS4EuK57CsPWM2hMX4xrzNzkFG4w7K5thnkoMB+xbPjTkGCi7MEyERITDG46+94DmynKhEUHxACQUW5oUEw+Z6NpSBUM45rrx/NG1kd++85/CRuZvk+SmsmIMyl7VysGcj/xAdX1J6pcq9SyNGQwG55+9+S/bRL/9t/Mudk+FPKj7HMObHaNun/R6lf63EHBULQNxjGWHzgjz7P7wEvAS8BLwENpYEPGGxserbl9ZLwEvAS+BsEniDfmThgVb/MNCm2/7eLXL/VLqyl2mFcdA17wW0QIvKzNoByA2wZ7FkCzkA9HHLCc7bEsVICPZ2jcV5MIsDu5bfzV+uaX2yGAO8Z7FGPllYmh9dixNgLpywcuDd3AOZwN+8C3dIACwsyNBswyQftzwgEsQbQMvNiAHuZTN3UEZUDAHC0bMN/Iek4HfeY8QIlhHkd41EWAN9zGKE5xpxY/EuOMfi1RaFdj35Xm+VYu6DTBsQywvyxHkIjGdc886m2/4DSyIskDfgOPmwhB/hv1ei7j1hMaroC9wZyYS8SbQzNtolG32ERDsySwrTSN5Q2sgXKNeLvnzkkmbwgc8eLBYWN3flAz4pg9XWdHzs5HzxSBG5lX5cLd8SuOMHGq57Yip6bMtE9c/c/Bs/fjXJCvq1/IoELdFV2zSCbZf7cIWyUFzeskwHWXmr3EQVimkxDL6riOFz7U7QHMRh21X9erOZ3jwfN+KqCjsCNiEiGA8Zn+n7p21XxKsQ6PqX6wR7r859jjgXFy1wf+N1LwGRfONlGFcaoE1B7vNtHFdAALA0yx6uv6HJirNU8LDssqAg5sfyVKsed3qDlaR0TcWrGCjItgIUu52yrEiED+vaQF7+tSlwuYJaVK6WFApwviJ7Cp10iQiMCfXnkzo+2e4OFtOkgfyrkSWHdwl1hXvaiKwAHwH4/xGl++Sqy6XNSZEVEyInwvG521puFIC6rMJ+lBTVrtuPPd+Y7pa9lfrhg49vW62K8Am5W2o0pnv7V49PHDn53PSE3C7tFXFRirhg3GaeR0JhCJKCuR/1vDYHXzs+HV6DJQNzN64zV1Ncy7wUSw3azVtG4jK3gUZG/LbOM58k8PWblP5OiTnq0J2VrClWNSt9RI20H0XliYm5dm33/c8d2HLbQkvWGMz3mdMyl+QZWI5gvcFm83y+RSjZoMBxXOLr3/61ebppd3n0qf8v/tDBR6PX9FaDGRHzbFyDUsfXKCGPP1ZCKYh5lHcNNRKs33kJeAl4CWxUCXjCYqPWvC+3l4CXgJfAmASkLf6w/nxAyeI8dF19V0Ng97xWLwLIBouKY3FM3mlZGA0XNdoAxs2kHbLCYj+wYDICwgAOc1XEIse+PS/QUhs90wB9y9040QGgziLIrBpYYFncBsgHABQjQHgO+fmwEm5PDCzmHIQLGmws3kxLDCB5z+h5kBVcZ2b5vAPAGTLCwGcWbaYxD0hNuSyAN1r15irDnsH1JhPKZpYX4y6rTC6UhWvtbyMpeMd43AqeY66oAMdtYQtgSV7Jz14XpZ92Mw992cW6NF9FPpQPjTzzP8zzH1Ab+Iq01P+Gh/rtvCWwBjqvkV8strFggQQzv9O0BbQGqct9SvQvq8/zfom/8OIkMHLtVPzeR58u5mfmBneu/JfudPFFud/vfimqlu+PqsGt4eCJrw8VnKdWHntEfcDc4LirYPEytAQTO5H2q2yrPL8kzUZ0XFrWchATKuh2OeWKMlBAXkXoVQBf+QZvxE5gZrVbEbpTuYohKGtDwFcuUuOIQE6IVtqhBeM+k9CIY/Ofld47ugACA1dxxy5Oyv6uG1QCBhayNwscvsdGsNPWcpGDnnQdjenEMGjUExGI7lmRELcI2haE7RQaJ5zUuZpMKo7X4rDe7lXMC5alqB/U5RzKVcEJBdzeX0vTlbSZdOIw6KSy1Wg1U4uh4GV89TsZ7Z55Y6L4FAtxrbEpqTfkDbUUaSHqSS6VSPSGpJ4RpNrtefWBudZcewds1NTWlb2t+fZnu0uNz09vX3pTFJdfo7G601uuP/f0p3YfW1mYuKe/Wp8ri1P8x57RGAwZYO4+mSugTHO6jfkrcwvIDmJDMOegXaEMYcoy9Ft+Zx7C/NEIi+/T8W8q3ayyNPX9uF/l6sW1/ABxaRRc+/jEXOfTZR4emrvp5PT2O49Opo1BTdcyz4RUwRqD+Y5ZZvyujomNQWFYExBXjuu4nms/ldar1qZbil2N6aozv6v88JMfi9++eCis6322nqCMzJN/Wun/VcJVIXLwRDqS8ZuXgJeAl8AGlYAnLDZoxftiewl4CXgJrJPAt+pvFjz4vwW42uMm7iyHsSviuVUXzyQumuGbweKCBRHEBWA/izoWQgDkLJLMGoAFtpEVkAEE6GZRBZjLAsxcQ/FMc4m0/l4DRozEuFXXYm7O+8waAc0sA1HsnRTN7oGIQVPLXFewyGLxBmj/iBKLKkB/noeFBSAMpAjAM++HWDC3UxwDCpJ/TN+5hz0AIeXnmIUWCzYWaiQ03cxN0FATc/RcgAg2K/u4tQn1YASJgUaU0TTvTC7cTx54D/fzLORKeVjoISvyut2luw+6yQcPuZMfRnbkh+u5b58Sbg+ISUIb8ITFqGIuYGfEGzKl3qgzC/pOXdFmrP15jcELEOzluvS73nDrkCRqf+x+Red+/lhYdWRdkTGeUHcQd9SR9cUrDpBIm93GuuF4oNgAiZyDbymrpBAhobGkmgijaE6NJioGJRraq9JGne33MmlkR7iKmRnkZUtBfJ+dmnRLjTSuoihgLBiOwWhjn8kt1MjK4n/XdUZYMA58g+4BdBqW3QfyvVwt7/p5joiH02X2FGkxssAYVygYguhmmXGG+68fAVxaTpHTUB6KL5OUa9YSTyk8TaAA2nmZhPVc7t0SdOp1Mk3KeZEYLknDXD0u0okVxakB2JWbt/hYVihwdxkyLp361p/Fzdul5dzffUoCI+sK5lDUJfPB4XxT4+/eMh9I9yN09VbfNWe6rn2y6Yo8dBOzHVef7O+f3LzaE0HxgMbvm0Rl8D2Z0d8P6feDOifFH3cH0S7i+fardt9/wC3sm1898uSWpLdSU3B7WdmtfYuYDzNHhligr52NfGaOwdyNdsJ81eaUzPmYw39WaY8Sc2SsRZibUCZcnlLGvbIIOas9ZNcAACAASURBVKbyhLL+eHrTnuOfFZnSjNKiNrtjKVdLnY/S/LHJTe1pkRkoM2GlAZlyjxJzSObSEAyQJlj2MncmL/zOedy20n5512EdvVKWFpOt+XJl823ueNqsfv0Tv5O+NusHr9bv49vb9QdEEa5av7zuN/+nl4CXgJeAl8AGk4AnLDZYhfviegl4CXgJrJeAtIrv1zkWaJAQLJxYZEy4iVeELm7KlXJ9TjEsjkm1zGIk4EIJssIWSOxZbI0TBixeOAcATmDhPUp/qoQLIgB5FjHmo9ZUzAwoNKLDiAgLQs17ANe4/8+U3qTEe8ZdUZnbKBZXBtyzUMPfBUQLBAaLKrTOAPcgLHg+C0POmdUFwD5lpEz8TmIBxsIQMgCTdbPuMNdRFgQc8OIppaeVWCxSPjPvx7IDrbTxMgJU8Dem9QZQWOwNk824JYYue4FLKf420ohjnsUCErdX5P+k6u5Ot+29j4uwIO6HuabiHVipsKfuT9IWpFn+OR7it/OSgAF6ZlEBuUW7oI09M5T9GuGVr8VY8NtLKYFm73OMOfR1+gDtHl/ZgCPm7o0+fMW3UZwA2oOsI4KOrCWOCeG8pdsbbEnkDF/+7bNQPIaAMhEZ5WQcRx1ZW4SdQZ4M8mJGLWk6k5so3SM3IsEnq4nKKRh3pWfR9w1wO1t7o23+S6WfHRX2F7T/wKi9Onz1e9LiijeD6+oFY4TEhh3HztIncNlk7iHLJI62VFUpYjHMJidqNfXhE3lefUWkhHq3m1G85p6sKlaaaZw7uYCbbKX7s36pQN3lCcYDRTfuidBgLjN0BzVK11V7uU4zy/jJfA7lk+9Q+qf8XVWFS5qhm9y8LMJCBjEyd5vcvOKyXuK23/n8yuR8+xGB/k+KmHhoVG6zikhklfBOnWMeDIkwob+3TG1e7fdXa4cU2HqHglhXg05qMR2Yf75JibqHXGDuyjnmc6fbsIzDYm7cnShlgMggjW/MZ/n2Pa60C2J8Zvvy78pd1eTkptUt09tW7pJFRZQ0slkRGciA+etRXccclDk/c95PjPa0SxLzG7PcwEUVhAZ5JT9mWUocDtw9MSda1Bcqn9xcHhm0g6w26QqpRK0nLMgzc2K+0ZAyLwjAva5M/k8vAS8BLwEvgRtcAp6wuMEr2BfPS8BLwEvgPCTwLaNFiMU+WNM4rrLUxZunXTzbdWELsgBwH5CPxYxZSBjwzms4NhdOLDT2jRYdLN7Q3sVMnM1AeNNMt78tXoXFvzBghPN8r0yDmOOvUzLg355jbqfII0SGESj43uZZLIDIOyQCC0KsSXgW17GYA3QeurkYXWuECdpinGdxiByw0OAeI2xGxRpqlaHJxkKPxSKLLhZxb1VisQo5gGaaychICEgYgFL7e9yqgmfb30ZmoIEHccJ5C+INOWMb541A4p49wzxt/ba6++IPYVWCBQhWJ+bvnmuROQtS2oInLMaEeR6HFhiddgP4bUQcMjUf1OfxGH/JVZIA4wNjEvXDmEb/AMihT9C3hxtB1a+CWyhZVARLSidETtB2tspSgvCulZSxe/L7VHX6ZdHPS2GbYVMMhVzcV3Vd0ZYjfCK/1nX9ZllazAoUPZiGkbnGo2xn3IhXIYD1V3SBERaMpd+u9B8p+lWqB/8aL4EbRgKjPkXfaYt00Pc+agdBmU00050KUnGkLFzYrxWb0lo4r4A06UC+oqoi2C8wvFAIhOUoDvaJgxRhIduqMOjqP8Dq4bfFW1dctWbCXIhvAjG9/ielBhRwUhsMLSnmb15yZTHdXTw415jZuVjWW4MVWVfIjZdcC0b4hxoC9swvxzeRV8Eriiz8LbmFulWExZvDuJxR8OqVsgwz3TS78OysywcvgGSYm+ECle8S7eCNZ5AA81jIFZsDn0lQ+/QD8zvmvMSneFT5eGpu18nHN99yfJdcQTXl0upunc9lHfKs9jbnhkxgfso7+GYyP2Tee2j4nLX5p80lmZMyt4TEYJ6NDPkOoShE4fi+QWY04sTtbcxUH918SzFYPR4/qy8O35/x7Sf0B23/g0ofUzqXm8Mzlduf9xLwEvAS8BK4ziXgCYvrvAJ99r0EvAS8BC5FAgLlIBZY7OCu6TNKLDamXe2m/W7Tu9/psgVpANYPKZ4FYD+ukgD1x9098XojL8zlEUA9oC3m3B9WQkPsd5R+ZnTerjeigmeMP3OcCOCZfKuMjDC3SORj/DfyZwAxz+MZXMO7+Q0TfUgE09oyU3UD9sgTliBcwzGLRN5lJAHnOGYRxaKM/JgLLItdYXEpLBApZMWbRvlkUceC0SwnxheYPJdF8rjVhT1z3MLCgMT/n733gLLkOu87b1W93K9f5+kZzAymZwaJBEEIIAGKFEiCSaRysC0qUZQla22t5FXyyiuvJMtaOcn2ofasvPZqrXB4JJFKXEuUKFGiCAbQDAJAAARIEGEwOXfufrHC/n817xvUNHo6DAYTq+bcea/rVd2697uh7v3/vwAxQvk4yI+D67IWKpyj/OYqatwFgzyDNkGebEAhL9B+o73Ij83pQfqEgFq05vJjYxJA7vQLawc+L7pWbOcfnS3MWTch2eKVgZrzY00JYOWi/s3cwNiAmGVMAqSgpXo2fsUlFGMUhlGkUhG0d1EAZyRg0yuV3clemIyEUTwoa4uk3Qub5WJwulCUkw4xFop70dL1JQGhDQXmxT/+kXI5YN7ZDNkAkAQgRIwfjt9Qwm94Gssit7K4hL0gf9S1IgGbm1OFCZEPXxX1eBpLKb/oFcuxl2qOdxOvodA0ZefHR5qdpNns9FylVJitFgvLpWJKOjI3dSFBrhXBXOn16LuDApzHmoA2GFO7uWojceNTZ3QRylVvtjYyuySCuT1ygzimSi8p17p+sSLLmWLE+ok1IO41AeZRTuHQ7O6Ni7T43l6nMCTSIvIL0aIch0kpyHma0acGJ5bL88cHy/qFNSUHSjas7d7Rz+t84qO/QRSY4sr5rpviB5Eqi+V65wO1Rvu56nCrODE13VOA8FnVU+7LEhRysIrAAoNg3JR/jxJ9EfdMWBiznuaZPI/fWdfuVuJ9Sp0pM+9T1o/IEEtnyA3u5RMyp6Yc9kuuX7z568KdJ58LfmF5xnv/KgVnxcOehPd1TlisIqD8VC6BXAK5BK4HCeSExfXQynkdcwnkEsglcH4J3K+f2GixMWazwcaj64bu2eN6Rxdc4/UVV90DOM9Ghc0cRzagthENbGIA3M1CAQCQ6wEE0TqDEJH7ktRNkwXnJi/zG2/Bss36wIB6+7SNnG3MOG9kg5XH3C6RJ5snNlrsNKmTBegmf3NhxSdAPfkAVlJHyson5IyBzrwrzfqDe5CTbaDMKoK6cB1lQFuM8pEHJAjaZmaOz7O4P+viCWKFg3PZWBbkgezNNZXJF6CRMpqsVsosC1qSB+XimW90b0sedX/rfVzfsXahfORvQQ+RG33hfiXcw+THGhJYoX1vMt8MYHxO7hlCgvM2nuh3RmTRlzlPH+M59CUj3jzdb5ZB3MM1tK1Zf8QiNCJdkyUJnc5dcHmv4s6BXBhDZi1Gv2cMQAQevFT1koudWP7/abOOAvQu+Z53XH7vp+Q2Znuc+D25gepJ03qpWPTDXuj3RGUcV0DfkY7n6svtXqtS8mdkZBGqRSu6Dlis3mr35nUNc9O6QKfA0K5ICUhkIyyo+v+khKuode+/VHLKn5NL4GqRQN/KguLavOvJ3RvgcyWOEyl/aEESMrSShULBq5aKpdOVUnG501OYC7l9E1lh65GcrLj0jc57lvcm8dY46rwtFWvBje1SoJFCnAxti3u14bY3uGX5oH5qFErRpCwVqgL7AeZpO9Z+NDCg/7KsJk615iuDyqfeaxe26NpAMSOSSj1WqPV4ecve05XhG+a9+RODinSyM1k8WS/hbkoHZAAEwvlcQZl0mOvT2CkrDhSPWHufPRRI2ymmRjyyff4Nsu5o6bldz487vpfI+2D6HMrPOxBLOyx+WQuzXn9e6VNKuCy9TyuGG8WzyDDIe7TbLn60VO39kM7L6i8uifjguayRkSHx23Cf9TcibB6SjG5R/SEzqNdE8UwQ7qmv/Z7OoQf+n8oJEfWTK1YjlIV4GzlWtUoD56dyCeQSyCVwvUggfwlcLy2d1zOXQC6BXAKrS+CbdBptKKwBiGURuJH7nnFj3zjl6q8pu6AO4I5FgblLQjPfwHY2ZlnLA64B+EebynzQcv1nlADGIBDOxFR4IV6DAahmUWBumNJdvRK/Z8kLC/ppZAJ/s9GiHNQDMNKIFwN70QIjRgNls/gCXJMlSXDjRLkIGAjRQjnMioJNFn9zDyAxm1Oeb7ErrMxWTjaRECRcwyaP60yr2967BkLrp7P1o3xcx6f9bgC1yYE8KQd1ZkNKeczSIws+Z9vI3F6dMdm//f1N9+QPYHHCZhAXOMS1QP6QTHzSJ3LCgpa59IeRDbQZIDp9EdCAPkQ/NJcTtD2gO2OK84wDwJKp/nn6IH0e4CSNFyOygnFgrsdSF2t9kqN7nREXyIaxjqwg/nCxBnGABRJjwKxlLkXrM94WCoEnOMmNCtQ87ReSUqnol0VCLKtRx3W+JN9PisObDEmz15UKhWIvlOPzxJPLmaSpiaEYyU3UUrPrRHJ0RVgwb230+Kou/CMl/LVz/IrSrymlFlxXmpVFhnA7a2VE39V55kv6NImxQEqty6xv96+BpMvJmI32jvy6TUvArCI0dhiH9NNUuSFOEoHDnoaor5g1aciCQf097xe8VuICX4SFxQXABVTeRzct+Zd8A+solENI30duuIMqKz7QoGbhSj05VhmMZwS0a90U3aTV3Zn1o5fOM5BSrKUA/nlv/3Uce/Nzxxrk9U29VnGPF8Tl7nLZLZ6qN7fecjIOinFDrqEa5YFuosDWbZEXfmu+qrgYZ6EZ1mfrHaawsPK6c8gKEQWuVO12qg2FRilGO5tzlUTuoKoiTSphryBiIdkmQuakiIV26hbKS3gHfg4ypi8Pc4l6o9473SgMBpemByoHHtkxccMrjz9dGei+UnXpFSu9J5RYl5wUUXOg0yzvPblvfHD64MhtO+84euPkzSd3iODgPcs6RM90d27ZG79yeFv872YP++9boT3BOwg3VKx3WXPnY2K93pD/nksgl0AugWtQAjlhcQ02al6lXAK5BHIJrCUBuUQpSDs81CcbLjYOX6cE8HnEVXYsuht+bI8rjgauffgpN3AbQB7aXrwvzOXTSusH/gZo51qIDzboxHJgAw7Yipsl02bGLy+WFgCFHFnXSPbd9i1mOWDkhZEj5GubF8rNptDICSMssmSHkRXU1YgNNlUQLJAclBs3KNQTF0mct0DfXG9ul7JAoFlJrCwzz4Wkod5sZNl08d2sKCg3ZAFlQm5GwFisA8pCOSE82CSy+QVc5VryID9cDrCR5Nl8cg/3G3GRbR/Kb3Uhr9e4re+RD+PysHvi3RAj1J+YFbQHxBT5PUPfUB+JrK/oXH5cJAmsYklh7WWkGBqIWL/QNwicfpsSYAibdohArGBo108rAbZ/jxLaiPSBtynRBz+s9Np+Hn+nT8Yv7Y22JKQH/cgsjZ5UmfgtO65eVNtryOUUckJuZpmFqwrmESMgL1JLbzibsNuLWlJPPSH/4V/ynL9PsbMnBXAuFeQMv1AsjEsre0EkhYwvQrWRAnIHvoiJwoxOzHQ6UXkp6Hj6fT4oBNLU9j0F4D4L6K9VCgGjPQGrEBRGWHD5bqVUO/ZSHuexMLIiMLcZwcx8f/bd0CcxmBshZBkHgIdcQ5vO63famu/87uvv1N1OPxlRnuRExqVs7eviWeYqkD7WEVFBn9W73OO8PLvFFjOsJ7LC1lbp2geicOWxRsDv60KYL2cl++6geEeiIGAWti5RS7WXPDd3zHfbbo2KhVLC2pZ5CKsJ1rq0F2tG7mFd91x/7okVVH00KET3KbD29pPPjZcjxagoVruuvVCt1YZbkWJitEQehLrOKeh2IeoFyj+UFoGiE23M7tGsLFkrrnmIjHBy/VQWLV4SaaHA18k2Bdh+yCslg7NHhhIFAF8a3jY/M3N45EAceafHbpytRaF/QPE5DolQEa+WsGZ4iwiNeVmNHGstVKaOPLHt7rljQ2+UG6sPje2aaasO1WK5t2fsxrnjMsCYe/6hXRMnnx97r+Kz3Kr6LO77wq7f0efD2249MSIXWrieYi2TBMVkaM+94dNfPF56IOqlsens4H2M9R9KF7+nxPonP3IJ5BLIJZBL4DqTQE5YXGcNnlc3l0AugetbAgKgTSMLkPs7lfApC6AJMLrgxr/lDS7p9lyhUXLV3YDyAPtsjLgerS3bSpkrKBOoxUoAKAIM5TrAcMAvNnPmKorNngGDfLf8KJe5vMm6OFppYcH1BjTybLOEAJQCwL2/nz95WywMygOJQBl47wFuYflgZvOQKHf2K8KG1dwyWZ24B8AYkMv89FJWzluQWwMI+SQPNleAbDzHCBezxDCygrpk3ToZwIGFCpplgNZsiskDkM0CMKJJz3nahnreqATCwf08055DlThHOZEF7QEp84zatuV2/tRd7tD7kAsbbgBK2pu+QJ/4TvUVNK8DfaZkyiUIQEx5r/nDgP++xjdjYUKtSF8I1Fp7NEKn9BdtTjvyy7069+r+SHlI5+7u/8ZmnjaDaFp54ILNLITu13cjzAAeIC3+UIl+SD/7MyWAFgs6DZBmgcOvxfagbkZYQA4+qgToA7FoY/qS1FtuoWj3SK6hmt1ueEqgpoJZRNt7Pc+LYjccF10z8F1T4CaReEsC0IpyJaOx7HU9hboQ0DlAwO5yKViQO5nI873V3IOsVxf6FBFQLErKJ/V9SgnLnYtmZbGCkLAyZed3+rtpOJslGQQEbWQxlOjT9Nub+hkwpxGXB5/rnLM4JLzP6OsQ0bgnARyjTvaewXKQ35AXRO6Mysecam4Gz1pmrCe8/PdcAqtJoB8oOxL5kBIU/b7HpfTzSGOdd3rWYpTfNgZVX2SR999FPPtFz7+GiOq1pMa8z1r1u5SYb3ZhXVGq6kW8O3Y77ghPNCaTpl9IrRiZV1g7Ml/8rRIKA6yhmEcA4lm33ShwX3kk4wsnBxu9dtHJIoEYEukMNHNwJBBhMC5CIFTA7rhQ7omEjhNZJ3TbS+USJMYGDsqJtcJ68SvS5xI0XO6o5MvJ+cVSSF1Pq7X9YjmcOvLktmDhVH2nyvkmESf10wdGT3aWy8099xxwW246dVRU26gsK56T9Ud5eWZgQp+d5bnqHYrJMTZ/ovHe5kJ1R3mg42RpMdltlw7rfHNpuvYW5X+nCA2qUul1vB88+ezEh+qjzT0KWD7m+wlr1nnJY2jy5uhVlcHkseas95YMWcONzOnp+lWkkv/wg7+bW1lsoGPkl+QSyCWQS+BakkBOWFxLrZnXJZdALoFcAutLAIB6sA9CsxkAGGV3tOCK49td/VW+KwzLFdTgggtGAa/vY7OhBLADOGTxDoxsyAJkAOqAXFhQAIDiaogNHO8aQNKvVWJzBUhrWv/ZnZnlaSB+FtA391PU0EAunm2a42x+2Cia5QPXmfUDz+Me6ktdzMoCEIx8AW0p557+30ZGcB2EBPmQADTZJJrbJuoAgWFls9gCPIvzZ0DoF2JhGKmRrYvVh2cCtgFikP8nlNg883yeyQaZ+lFn5GzWHpBBViZIEgA+K4eVm2dwjvZDFmrnuwPXeHbRjX3ThJv+C86TNzKErKDcyIrNMOVfFFnxYpVPcs2PC5KAACLkStsNqAd/rVdS34olbz/tY++Wt/OaAJMj+qyrxXekvfxMb34tgUA5tLG/+WxI9fREmj6n/yHf6ENYDkDW0a/tgHS0YJr0Q9oV4MXcvgHe4yYIMJd+Ye51LqieV+hNSAqJflaJ+QCihnlj5bi8qMUXKbFWfqlllciHrpd4SS9KXBy7o54X1rsqlYJstwM/WJLLqIasLdoK5rvQ7oSLCsQ9XakU9ils94FWpxdDbCw3u9G737hnw8BOP5bFr+v5RlhA3tBHUsLiZTiy8xL9lHnG+iVjgncUVl8H+t9tjrN5CjKOe+i7P6D0iNKUEhYUvGf4jTFg7vsgm7mXdqZf36PEvEpiNO1XgrBlTn1Sies7GqPMpzbXkpcRz/r64uM6AXZXrXt+8vwSyBAXWaUGbjByIP28VBYUGbdqRhDS75kPKd+1Tlafr6FYF7HmYS2IIsB2P3DhwEhSaEzErj6eLCoGxLxaDFl9QZJi3cyaiXUVijJvUmLexDoyAtwX8fC8CItJkRABcSkA7kUGON7fIgSczjtZKxQqXekkxL7c/sX8nugZtv5cb1id4/ZplYvJhzmsIYuHIlYWhUrYFmmxVKr12iIxhkQsLBx9ajKSy6auynVSFh+75MpqOYn8p2Rh8eavfOJm4ms8u/u1h0ZEUoRLpwcKpw+Ojulzdnm29hGRMu/R+R1YhXQWyy4aXR5RZ35TU+HjVf+GES8pCZF4EyJF3q267x+cWCr7lR7yhmzeXyi5YyLjh87D1vE+QM700c24O1xPfvnvuQRyCeQSyCVwFUggJyyugkbKi5hLIJdALoGLKAEW/oBRgOMEXuYTl01fdaVtIyItluQWqqwNWckFxTfqPNr7ADtmdg4Aai6SDJCneGwkAJAgNACh0AJnQwVIxDOJi8A7J3XL0f9uBAj5GHFhGrDm/sM0EFOtRCXO2zmL9YC2bKqp3C+rBei2fE0DzYJM8zfm+/Y75SJPKxsgpv3Gdwt8/ef9+r2DCvfrxWb19UoWHNFIFn7Purvi/Gp1sT0acmJjxj3Img3xwf5zAJNN85vfkD/EAvLjHjal5h7K8suCIzzXCBeyvFUqdx9x4dykm/rZhlv47Jdcb2ZK5yE+cOUFaE3fMNdWl9Knf7/K1+ZHX5OVtih5Gm3qzQMKQ/kNgs2/QS007o9oHPpuV6we7Y26CV+9L5Y+p0eLC37ARYVXdstJ0w0EExqXwkD0e42eIFDgcY2AQ0poTn6z7qBNAX6zro7M6oj+xcGY+NmMtCHG/lelv1Si31hgbwJ2A4CcVwP4KgJsmUMYr/R3NO+ZNxjjfJp8LnoHlDXFWnkmIjR6cuu0NFArHJH1xFLsYo07f06xLHD1pNAV/v5eN7xBISzGZWVxUgN8vxpjfmm5Oy9CY6bZ7i3JCqM1PFjZMFmRKRBWZj+m9J/757C4eJdSOvZfaiyLPkhKP2Q+ZV4xqzsIAQhum8t536D9a+Qr33++316P6xP3hSsPs47jPGSGHczzEIC8h2hfnkV/X6m+DNiItRr9mxgmH1RizuVdB5kHccL9yIhPxoB9ktdVbY2hfmcKAMnNu8a8mfmWPz3XPEvO9K2AVhF7fmozEugTF9xyuaworJ1tPcQn6zXGuFmB8GnuKTdTvav2WjT3VXiLEcV31q4iGDQpTXsiF3w3eatXqTXc4dpwsluzB4o3rB+5ljUyoDtrTpvfFgXk/7XcLE0GpfCegeFWcebQC00OeC83Ue7Y05OyeGi7LXumnYgDN3N42MnVkiwgNmRdsZ68mT9ZFzOndaJusK21WAnkikpWep6T66ZlPfOE4ksMnHxuYkJkCmv3hkgKLNOoR6qcIwLlTllffE7urA53mqXTneXSZ1XGumJYvEq9mHmxfyRaqyZVETATIi48xcs4LRLjxqDUlkutsotF1IgI0frFe6w5Vz0hkmOr3F+VReiMiig5XRuOG3d+U/fYQ39S+mSv7b15ReV+UX+jXAAxnRMW67V8/nsugVwCuQSuMQnkhMU11qB5dXIJ5BLIJbCOBNiQ4Nse0gILCN4DaJ3ucAO3Rq61X9pYpZYbuN0sD/jEBJ6NrcVjMAAcAMisF0w7mY0S5vFm+bBf3wGZzHzdrCe411w7Gbhu7pWyQP9ZMEXX23WWh222DdyCUEBDzggRIzn4tF2gWUyYzjqWINxj7hlMfFlQgWv/RImA3GzmuQfAjU0dRAMbN4B+0xw+o+t+Lglj9cgSCVkNS4A0yoZcAPXw2wuwt0uJTRrtBZgM2GqEShrMU4fVhc0p7WHyWPlMwGe0jz+p9HrnV+Zd69m2Aqzf7o7/rgVzpp1AVsnrh5U4D4Hx8f6z8o8LlIBA24I35BreoKyMIghBASOh+8ciJt7pAZ8L8vDG3LjICZGGru4LqvXU0imU0IdHRXLQ2gN9u4eSLDC6SVcEhvqEX3Nbk2XFu4j0T6Mx9bYdK6dE4zY5SzJmS08/ASjGxY4dPIE4GIwJAq/T1/cqUQr6Alr3lwVwu0Cxr3Yb44KxRb0hbgCi7ftFQYsupKx9YDgUgLxYq5Y6cRJHim0xU6sUw6Ln1ST1aVlYeGEYLsSxPydriv1h2KE9uvq+oGshPKJTM3SHzR0CU1siJT6gu4ywuF/feT9AyG7qWBEYG3la4FZIUOZPZD2lBOHKfARJYXF4cK/CvP4jqzx0NbJivbJZHCCzpjtf+xohzydWavR5rv2MEuAk44F50yyQbH5H/pB5jA9zJ2XPIC4GAcG9KzWovfqaPzpU9TvdKKiUA292vlWWa7JKrVpsKeSCeLAk/M2PPhXe/cob4gzgvp7M898vkwTWcLtmayDGosU2Ys3D2o/1BL+bW0n68abnkMtU5YvxWFtTMe5RBEmPVDnAc0d33RUljYnEL5STWzQjMD/YXAGAzvsDF6Csm0IB/20sKRZPDbwt7AYlAfNzs0eHOgL4q1mJQhooKLVTMG7XbZVS6wsRHFha8GjWc9n1oxWJZ1DGjRxkhKUY9Tmh53dnDw/PiyRo1xQ7QwGylxTguzx9YDRQOYmRxTqTNTz3QBJj/YDCjK+yVY99dct9qvsulWpOhIosAbW68N0WTXTP+sXopkIpIhi3k5sr114uPafI3odKA93XNiaW3MLJelrHQjFyfiF6bX1s+WOqv6/rI1EYPFfEhlO8jOQRWbLMzYmuXxHDg7mbeTYm1ojcQl1PBfQLUQAAIABJREFUfXMjbZ1fk0sgl0AugWtaAjlhcU03b165XAK5BHIJvEgCWBGw4EcrFbASDVI0XAUT3Zy4oXsCVxgvucoeC1DNZoxNGWAlGzU2s1kNPXOrgU94QB00VAHWLQgh2mpssgD3eS73s2mG/CBv25gZuA7MSp5cYybg5oYqS2RQYn4HTOJaSAMAWOrDJsg2NVmXTNxjZQewZMMOMEUQa0z5gYUphxEA1NnKTB0A1SAOONjkI7939+/LarGTh5Eq3A9IR33J3+RPHmeBrf5zKBsy4fx7lQCLAfTYsNEegMnUE6IHmZAXGznuQ66mtQz8bVYhZpVifpdpB64/7Sa/+6A79aGdandPMUvaLlygfakHPt8hnegjf61kG3TKnB8XIIHuz6gNE5ERI26rv0NBKJcUODt23yVriTT+hKf/vTM9KA1GH7zihYekZMbK4ww15nkFVy7c2+/TiWuIsGjLccWseupictqV4tMpKPyXet7fX2EfQX9grNA/s4QFT6KPf4vSP1P6JSUL0P0JfQfEMFdRFyCJK+IWgBnGL+OJMcTcRR0B7C67NRHEhYBkxu+M4lKEaaTtnmvIRZRicbugG8a1wPPm5DukIxdSRZEVnSRJigTlfonSZS75KyUsKziwtMHFWArEnwcMtUfa/G3ayvRa7qOvMLdStm9VAgyjbsxrKzVpX0rxabusFZnlZSQ4c7q9R9Z6DtdB6tv+CHCXdxLvNizrqM8vKP2Pfh0YD4wX3jNfMFnpMw36LZmlbvj0iSyo93mtXy61hVLfsqIgUqKg/jPQ7kQ1P/C2FIpBTf5ppn3PLUZhEonAaO8/Mrv4B5/e19uMq7GX0pj5vZuXwBpkBesHW7vxfoH4Y95DA/9PlXgX8PYxq6HNP/zqvoP1FKA9ID1rx/QIdHb3veH0tldEZZEVAyIwPqpRjjIHVlzYPKJkwrxAWlDMh8ejnv96uXq6sVzvTsnaYEYWC0/KSuEj3WZR84h3Nm/yh6SQYyalF4z61gm2vR5ZYcQq62/mwj1KuHekbedkUfHni6fqpxpblkYULHtPe7G8PHe8MSPygPnOlF9wjccczcG6gH7zgyIXjmql0BBRUS2UQ09WIweGti4crgy2PcW0+EeeH1ewGpFVRbM21GoPb5+/VbEqlonbsTxbdfGSf9orh/S5Abmd6iiPGbnAgqhGdqy/y1HoPT12Y3xo8aQvV1nWCmc/36NvxFRjjn2p77kXZZ6fyCWQSyCXQC6BK1cCOWFx5bZNXrJcArkEcglcVAkobgUAHZsZzNgBpNkpAaDwecpV92xz3blFV9nLZofNEe8IABfAcgB+s6wwkgEQxrRKAaA4b+6VAAABqtgIkQdbEPI0F0vm8snqyO8QAmwEAXvMfZLFY7BnZrWruB7AF0KFvHHtAWnxoBJumsgj6+fX6kr9kAMA1n4liAtcw5CPkRWUm2vY9P2+EptT07qlfJSTupCnkSAG2lmdsnXjGjZaWeuLLFnDc5ElGm6UC/nwN25QCCjLeWRMeSwf0x7muWatwnPQmjSSgbqSD/EM2BzivoBris4r3uBqt4auMFR2tVvqbuEh2tmChFMG+gibykfpO4pjgTzyYxMS6GubeyIjiqIsGrKweIu+vVZ/T3nDAgQ8gdCrERKbeMbZSz1X8eppSnNMxt0X/GWNvcBtSWbdR+Vm6rTCXH46aam/J+7rdcnf7/eFlU/DwsKO92W+/5a+k9AsNTciF1LSy32PWWAB8AA2o4W6Twkyz/3r46mLHHc5XeEYaSGrCWm0uo7IiRO+55XiMDmh74PiquarleJ8FMeFXi9yIi2Ybxnn0UsoN/Ppv1AywgJwE/kQ3+d8h815gGLMiRCur+t/f1ifzCkQFbgdhARbOe9frL5wvlGUPW+B59d7ZnZvRF8xcpr+wbz400qQLW9QAhDcr8R7CIKZufd5JeZNSBQIX/Lj/cR1uJ7ifWNz+HpleVl+h6wYGqwUFA8F+dTlSmwLpIXvBdsUDNrJDdmItMuXBFDGURgtzy91jhUVL0WkRSsnLV6WJrnYmZpyB+MSoBhQmv4JaE6bY+0ELU5gHdZnjHUIDIvVcrHLcyXnxzqMdQ9jmjVeeihmhcB2f8fCCf/AyI6orpgWyHS/EuQGMmMdzZx5CgtGERpHipVQcYb84yIDblCMB2JXLMmV0m65VDqHrLBnrEFQbNbSjznaFA9szctcwxz8/UqsU2cWT9cfePrBPRrr3p1aeyy42Nuvz1jlZ/5ivvr/lCgra07mauY8+omtTwcVvPvQzW94vi1iYkoGf82l063HNE9sU71bsrCIR3fMsb4cExFyWNYbX9Y8MlobbsYEGFdsi6dkW3FIzx9OZD+Kkyjy1jW7dr46vLlQSp468mTw+bDr8Q7JHlj7Qp6zHs4JixXCyf/MJZBLIJfAtSyBnLC4lls3r1sugVwCuQTOlQCbq29TQkMMIgDte4CVMyTDwqNdN/6ugouaZe3WAPPYxLE5mFLiXjYwXGtujdgMm9slADMsDrDWSAM1KwH0AHKbVYZp8AHYAG6Z1QGbP/Ix6wLbbBsYthpZQc0M/KJsHG9VAri3DQ0kixEcZilhoJVZOqRBEpX4JB/z2c+zAfjRPuST67nX3AfgCopr+NvkYmRN1rqDa5A1dSIPc53VL/LZ8ll8gKn+c5AJm0jy5l4IE+TGwW+cp34cRu7wnefRbuRn2rzUD/IBEga5o1E+Kfv80PkDO1zSa7uh142KsKCu1IE+wb2Um40reT7Uf1b+sUEJhL/m/ETxJUQQDMsN1I1qrbeqZ/6wLCDa/oTrirxYaTF0bs6J2kskxAYf96LL5FrqXnMEJcuOh+ViajHpuF70kDuquBe/ox4CWMV4ReM2GwfgfI/8If0AGAKJQX+4WkkLIywZQxB7u3tJ9bgAlMMnw73htolBv14rJXKF4x87tZgSjC+BBLjQ5oMwYQx2BS4zfm2uYV6djjRoe8sd5lNz9cI1XI91xqrPXCeGht1D0Gn8hUP4QpD+lNI/VyJ/O2xeNqKW3wBBiVPEfQBeEKyUj371ExcshNVvRAv4j5GD0g8oMU8BuEIW0F7MlQbeQUSjwQthYtYfmykO8yXzbkpm9Q/ytvyZ081V1Vv6v1MG5l/mae7DGoPrKedXlLgHgDElmJTOa3WxmYJu9FrIioFqqdTthVVZ6AzJzdhOAac3FhUnpVj0huQKqihfUPVeFAX6DRDzaKvdG+12e1+t18onctJio5K+bNfRz+lr9F0UHOiLjGWsQZm/LTYN6wdAbdw9sp6BXGR+uW6OfvwK5jHmL2R09pDGvwgL71PdplsKClIw8KVs8ILFGfK1tV9Js3NBQPzNCl79KZEV7xRJUTn57MROTQTvFlkh1s9f6eZoIzLOrnvXIzBWWkmSP+vrKSXmGw7c7X2byiISIZmQpcOWIIifl3uov1NsiorOs9Zg7lxJrrAeZE3Ji6UlUqYm105SeNHKJvY+pnxuE3lxh85Pypqkq7+DoBB1JZOjo5XefhEcz8iioiHrC+bnaQX7npR7qEMqA+sH8saypeyr147tih8YHI8/0JoPWHdmrZYhgenPVbXZQu4WaiPdJ78ml0AugVwC14YEcsLi2mjHvBa5BHIJ5BJYVwLSkF+UpjwaswDTaE0B7rOpiV1xZMSN3Fdy4eKM3ANxDZsDCAg+TfN/Kr32DMjC+wNrBgMtjWwAkDGf5QDkbLTMasJIAzaI5qfX3kNmtUA9DIDPbtKy7pOsrmbdQR5stMgDkIjnsJkEMKOs5grErDW430A3rmNTjwUCmyeu5z427lzPpp4gi5yjXlzPvQBRFr/Dnke5zQolW14DFXlu9nvWWoTn8jyTB2WmDLQPG05AM8Aj5MxhPtlXWr3wGzJAFlYG2ghwD//ruOgy643E+WXlG7Rc4+u0Yf8v0gKW45kzIK61O31lC32n/9z8YwMSgKyQlMdEFNymlppSnIm3eIvuG0U/TAa71ccIt73ecYasOKnefEotSfyUCz98uaBCk7HmBgpf5z6TzLkPRU+6x0RcbBGc9Rf6DeICVxD3KwEWmHuJlc/8Dp14u9I3KD2mRL/MgtkXXsZLdycAHoD6ltgFcqfkz7e98cGFZPeph/2fqClotS/rBXlYigN9JtL+TP7Lnz8Z/eg3327E6MtS0vMRDX35GknM+LR5j3IY2B2/VFJFMQoIrk3eP65E0HXmxZ9R+vVX/qsGruiYu+i3zHuAewBbgJzcM6XEOwUCweaw73uJggLgAkzFOoG5jzLwfuE8lmLUnbmNuZh5ivIxp9o8zBzKfcQDgpBmHqX8aFHzvqDMAJUQNMz971TinUh9yA9wl/l3s3sls3hjrv5FpQf65UZWb1JizPBMNNr5zrun27fGyr4TdPqF4yK6jPLUuYsK4j5aKvj1XphMKH7FuKwsKt1evLtSlIOX2NWiMB6V1cV0pVLSPJQIUPSjdjeKB6r+8Y88cqT3jXdvv9rG/TnyvEb/YAwwHrAaY3wyp2NZAZn49zJ1Zv3AgbUAFnNorzMnZucWdxH73JUqbsY2azzWTC9YY2kEA6BP3R3+0cSe+N7UCuGMXG0OSV059o8tmnWO+wogffzpLfcL+L9JgaWdSAsNm3QJpkDam64+a2/Gl1kbb8SdXfYh3AvJgBIPazk72iIKBgqVcK9IBm9gpHVnodw7qlganz7x7MT9sop4m6wfVistcz5WDycURPvo9MHRqDGxGOn+18g11JKIDxEYbkTkxwG9LlG0YD6dDArxDQr0TX6RCI1lPbuGdYWusTU0axzI5mXds7856z0vWe7Q93Nifuh31j8QRrwDPqmUW1lsukvlN+QSyCWQS+DqlMBmF+FXZy3zUucSyCWQSyCXgEkAwOcblQBT0KpjA7bkxt7VcMFQxzWf6jlvGCAFkIiEhiobOq4zgoPNBhsiNnB8ssnd38+TTS8bm9TUW8niQkBeAAKRTza+AhtnNmNsXFJt5n5BDWzn0wAoIwvsGiM9DLw3SwfKyTMA6dk4WRwLsrb82Niz6QEw4jo2+OYii/wBqygXgBVlt7qahYkRApA2Fp+D/LOERJZ4MWKBayyuhIGQnOPZnDfQjU820CYT2ooymosSLFcoo8nEgEuuR5ZGyJh/asqLJpv5UQck67ni8KOusv31rjujfGPqZm4AkAltNaVE8OXLfgg8W1kGk99a2ofZawQ+r7oZv6h1S8mKrjbhvrSqA8k8cd/rldye4A7J8wxMtB5Z0dY9H1b6E7XiISXceTBmAVkhndAupy0ZZyTce2zkQNv9Tj39DgX3rhfe6P5Q1h7PR4+6w4p18bCIC/oQQZfRkr9PCY1cs+LJ5s+5X1H6D0qAXfSxS6olvpHKrnGNjRFZHXk7Y6/s9YItJw4UfrDdc7cPycXShGJHdKWF7mRt0VtYbMv4wjXf/7dPLx48No/LpZelrutYQGA5sZo2/uahsDUEQ2BlkRb7dYnF6nFeHP77hdu/80cbT36IfktfBGBivoLkok/h15159qUc/0k307ftvXRI3w3Q51lmscDcZvMkz8PlEvM4gKORvrQPc7bNlciI+e4FZ/Fn5kdAOCPn+SR2D/l/Wom5jzoxxwL4Af5iSWFAL89eSerxzNUsogDaSByQfFNK1OfPlagnvtmxGrH3WNY6rn/bxfnox63w5GosLhQCWVL6N4qHeKU808nzUzyueCk7e2GsEClyE+V5YbHoL0o13NdvxaDoT8RJsiRLjI7IjRn1kzwQ98VplouVC+9vlA0Ad1m7AHoTvB7rIg7GB6RZGiep3wexPmLc8XkOWXGxCnWl5tO3rmC8Um+zJD6tmWG8oJliYCxebGyJb2sveo8qhsUdXpDKlXcta6iV70XcPxUUUPq2mcPDCjJdlLOjtZYl60qFNaWtnVdmhPLIau/lbKb2XjA3nqxzIaAnNbYXK/WOpxgTi5VGW7YQwQ24a6o22h9RcG5ZYHgfkDXEvSJeUHLIHlpDejcqHsfk8kxtsVjuVXV9Uo+8P6mNtMoiISItr+hfKMUwZ7J3YM7Fao9A3cS3261P1jHInPmXmBSsTSGAZuV+a1+nJTWP5KziT/b5yJ55mnkyJyzW7UL5BbkEcgnkErg2JJATFtdGO+a1yCWQSyCXwEYlAAjOBsjcA/EeqLjBe4ounJ13Y++8wQUlNhMARwA+gORsEADuAbFxITDV/41zRl5wDZqvZpoOuAXIzqZrvxIbLMAfNk78xobDLBQMSDJLBXOpYXEZqBtlMQLA6moumAyc55PnGSDMJpznnqnjC249Uo2v/rXUk829lYFr+W4kBxsv/s4+C0CJZ1EHAALyM6LByrbyHPkZ0GmkSXYjau6B+ET+lp/VzTT6TAYWo4K/VxI9di/5WOwRNoXUGfmz4eVzzHmlR1zn6K3Or4y6G//ZkDv4H6kbdaXeZiFzsaIsmGxW/TwPIbHy2iwBYX2Ca7IEF38bYWbXpJrX/Wek8no5yIvUDVRTskvcqxVQ+73ehLvVm3S3+8Pqf6VViIpILtMCEYPdFDR6Qj2Nz4dVm2klwAb6LZqSv60EGEA9GVcAnACdAMgAKfcqAUwRJHi9gzH948rpM4qjERTuT/vDoe4H0/4MAcdz0Mr9M6UfVsKN3Mrjfp1gXOAe6jNKgBMXFTxfrxIX8rsszOgPqY/t2JW8nqstJ15xIiqM7fSCSjcWAKOjsrDcKQmU7Qic7UkTXSfdaYG2R+QqahniQOTCJdcu7xMaL7uMt/35Tywef9ev/s9Jofx/I+PEL3xXsHwKKwXmU/oXc/1dShBbF3pAun1e6dZ+f/sTfUJQAGbRD3m30A+NYDWSwmI/2LzH+ygrE+7LHjaHrZSbEcsQGczN1AmrB+ZZxgPnIeIMNMQtINYeZlECAXF/5kGMF8gIrExwv5d1IZUtD/OuWcm9t58fz+N+7sFdI8/l+dTF6ntR213xKBi7E3L9tFvWFBPtbm9UE0tR/bwidfCCHhZESdKN5LhO2tMTBQ0GucQZltZ5od2Ni3HS+Wq702M9cMWA3GtYKCH/9P3wUq2Qsg15qb+vEfSeumXXD7wH6IdvUwKktoN+bmQF5/6pEmOQ98kln88utfxWeR5jAEsx+jCy8iAr1M9dUJbxacHtq40kw4qysJwqEJxZE5EgM5lXmDMYyzDaBcVrWFQMh/HOUtnJNdLFqJ6Ro7Yepo1J65EVPJt5C1d0rCF437E+cHJb5bwgvqlYDh0BsTvN4qEte6aboztnX7Praw4fnD06tKTA3PeefG78Nc352hk3VkoiY9L68LeChJdnDw9PK+D2sOJWvHLu6NBDW/aefnx42/x+5Y88IHrZC3xW922VTL4oq4wHStXuoKwsWFtSHosRx3z6vBLvk1qlIe9ZXY+58G+UsHjLHrRVakknssnL3UJdjC6W55FLIJdALoErXwI5YXHlt1FewlwCuQSuEQlsUEOcLcI5GlUXGVhFKxTiwAAgAT/ekitvH3L12xuuMLgsCBPghDLgToNNE6AQf/PO4DcAFvLgb7Ow4PwBJQAnNhUA31zDBgb3HWjjUje0/tCGZZPI5s/Ig+ymG5DGymeyMBCf3rDS0oJzBtKzCeUeyswmyEgQA+v5zSwxICrYOJmLK8uHT9sk2rM4B0jG32amz7OoTxacWllu7qO+RoRkgfXstQZI8WnvZrs2S+TwnU0ess2CWEaCGNFi8rTNIWUgQCz3AqhhaVNxhfr9rv7qAdebLzq/iowByWyjTPl4Dn3mUhwrNQkNVKROZpVi1jNmDYIMKK8RUNZG1MWsd/hOO/Mb5+ibwuOSczTWX8o4g6iID4n46sgqputuFlHxzf64fIXX3ZAqFahHropgyAv0B9Ta+1Six/T5NNqP/bJa21JmwEsOc0lEXiYTCI6DSgSjNOsYxty3K9EvAa+wlOK3rGsIfvtlpQ8pIcsPlr471fZui7gAwAKMRNZoQAIo/GS/DNkPNM4BnAnezVxBH7tiD5EVNocNRK5SlTuonVESjLW8rYOtZHyy1QuGwjiuVCuVZQWzTlrtsDdULxwbblS95Wa3IrJiQVYXyVKz2xE42nm5LC0uhwD77ojOjKmHf3uiNPPcgQPv+bMFIVwpWdnZ8sp3Dxx4cFCIFWTXhR6Ao/RX5vcHlcibOelpJd4dzKXM2xbPh/F5loyVe5oLAVWzZG623Nm8eqo/ZeL5zHX2LjFrOvoNY4Exw28Q7YyPTygxt+xSgrSzgOP8DrGD5cnKY6VrN8bmv1fCdQsEEfftVkIr+SElLBZ5ny6ojEberJKtXkr/bdXT55zsB3MXJuuV1MdrYiFSpQEdFcWuaCRJfFo/jsRxLMiWMZ2Me7G3p+fiitjejsDbQqsTisjzpxWDGHldMYRF1kJJ1h/e0/tPe4MDZU9xaFIZ6NPrWymlf1/N5AVtpmTvR97REGqMJ9rk3yllLYFW6xgAwow13vcIKFT/uaik2Pq98bJfwTuRdSmkDsS8BoImQI36QjFxQeCeLw8kt1Ubrub53kH1/SfCbmG/4jfcInUHZP01itUwEPaC9uyR4ccF8u/Qp+ssW2ifC6of72DmhCwpwRiztjEFlvUyZ17l2mFZNLB+GJc1RbtYitqKMXFyaHLBk1XFTLneCUdumN8WlKKtum58dOdcu1CKRpvz1VavW6iWtCQUEeN6rZKLQsXhkNUISRYk7WNPbS2ItJhobFl6u/7eIXJin0o5o3xwMblHf48qNsZjIiyacjn1XZLVYFCMRxTDgj7HfDmlxHy4V0mBPjy/tVAP20vJqMz6JlYJ+oHixtuVeF+w3siPXAK5BHIJ5BK4DiSQExbXQSPnVcwlkEvg8kqgT1RkNcOtQAbQmuYU5wFS7Fr+9nW/aZOurEi6iRHYsJkKAszwPMB6tD1nXXGo5k79KXEsWq60A+ATEJLNAZsmNgZcb+A8zzKrAnNjBEkBwII2OMFEAcS5hw0xABCm3JQV7W1AHTZgbMqMnDGQnbwNgLYg33ZN1p2HuVcykN7qb5s5A7w+pR8sWDaaq2adQL2pG8AsZV95GMhlILO9KzlvYBabLgAsK5flvbIu2Trx/Zy27T/Y6mif1t5GvBg5YeXJkhVZUsNcZNk5/jYNYWSO+xY0pU2DGbdCz7rCWMF1T2rjGAWuvGvQdQ6glWdgv8UpWUVMmzt1HsLO2sxkm7VUMddWfBqJZZY/1IsEUIO8APUA5M1CBdcB1J924jzXAMzQZnynXqaNncorU75NjSsBiX58XM8ouLfIe/Nbvbq71Z90r/eqriqNROJV4FLoBcKCc4lbVsjJzwua/S1ZYpzWNW1dAeBvMSFWA4+s79CW2fkEQAJgk3oZsIp7G2JRAMicz10PhB6JAyDg/1J6UMRFahmluCVt6qbvH1TCzcOb+tdmPxhf/xC56lrG29IVDnwh17oaZDT2KsW2m1w+nrwuacV7G2033JCffupbKQQ+BFej3YsmGwPlr6pvjMtVTk9A7eFquTi3e8fIwrVAWvTbl7HOGGHMAN6NDOz/zHc3vvyn8wu3f0dKWMzd/d5XDH/x/c7v0T3XPADyTYsbsgswnvcAgDz9lDHI/AKJzSfj2mINGUGx3jMu+u/0WcmCvmHzON9XgvHMGfauhmBhrPE37zv6C+9M6seY4D36O0qMv/9Fyebk82lHo00MAciBdrIRksxRyAoLJuSHLF+ySzJZDXV83zsil09bZUVUkxu07WGcbNG5Yuziluf7PVG6DbmzF4eXjHlxPKCX6lNCK0f9yNtTKVdO18qlY4pl0brSYln85kefCh758pFAq6ayyk77BN1u6FdKxahWK7bUEOH0XBMXay857stF74jrZ0g/om/wTkTjnHUcczh9Z6VFxWq5/aZO/oGSKSLw3lxU/3/JfWr9ol9xVzDGWRMRlykdoVhXKOJEGr9CLqGq5ZrrRWFhaO54faeA90SxKe4fHF/eqigvYXuxslAdarnF0/WFo09uDWRdUOkqbsVm41XIfk8PTc6QAc6b03/MJ9kjSz6ZBexawmTugbBg3S2CIPnw4MRSe/Lmkz2V/Usq3ykRLnFtpLm9WOlhQVVQ3ZnLioViONyYXJjX+cOq24gsMY6KvLh36XQd66vHVOdY5MTNKusEde11CpHk8ojk8gqREx/bdsvJo7r37cpvRK6lIpE3X+/78Q3zJwaLh750w4HhG+a/PLZz9rFyvfsxERj0wf30P+UX6NrS4S/tHS4PzMnKZfmzYad5d5KGVDvnyLrKut4ItituAOUFyiWQSyCXwKWQQE5YXAop58/IJZBL4LqQQAbwzBIR1N0AdgOkzW8uv3EtwAibULQdATxME9isCthMmM9WAz5tJY8Lk3THs0HigsCL5uYIMGTQDbyi48a+oeSKY3JaU8eVABsJc0VBmQwcNssE004FpDGwCSAZ0BRABtceaPDzjgEUp76UF3KAupGn1b3/9ZwP06Y34N5iXnCvBdVmo57VNssSATwX8A2QlQ36tyqh2QvRQp67+/dSHmRnm8CV2muWZxZMN6sIs6pYzWd5tjKm8Z/Ny4gWI2XYJltdDTCzPkSZs4xUFqi252RJC8vbSBdzb4VMLNaAgfiQSWMuqElWYr3G3inY/LmWO36ANgSZ5F76Cn2G2AYX41hZfiPDeBbyQD2R7+aWjL/NMgCAE5dj/A2RxvWANgCk1I160T4AfoA4AIgA9xy0F5YIaKACwhrZRh7mE/nsmNK582lmnyMDNNP97SpP2b1CxMN3yv3TfV7RDXhDZwJ4elEafLug0dTTNWfq1XW/qhZ92FOLCE47pLPUKxRBsN4GPPu7fbdyxrIg4GDcIjuzZPpZff8hJSwu1joAvMyHPxqMEJALArKaquMX9f3XlABCfnyVTN6rcwCzWO98SddDWlyJAJjNsVHiCr3QG6ouBHdMn/LuL7fCUqUZjA/HiVdqd0OBOL7qkgS9Xji8tCz18DW4AAAgAElEQVR//gW/5XnxgLTQB4IgOSjioqP4FpFAz95VrqnN+GIehKjYpcS4UdyV+BvGPvfrToTFmU41cZvrjt/iKsfVRVL+/OzB+IGkIA/GHjFNANeZF3FbBsjP34CkzDf0Ta4zAvJsRhuxEFil7120U5nnrzoO+4QGZTerQt5LHIwX+hZEH2Ocd6FZgv2lvn9SiSD1xISBcIBkXU0N294pfPKO+h4lxtRvKTHfMX99QslcVRkxv1kZSJfZi0VUxMJmlwXqd0VWdHzPtUVW1NW8FQUQTmJfPtMSAbaxqwrATfR7NQiCksi8pXKxMCi3UoOLzQ7rlQuxfNlsmde9XlYV/qHj86WZuVZFdRoMAm9Y49WL4iTu9CJ9TVpLy515ubdqVcqFXrsThhq/qdXalTCG13D5RBHNmoL3OO81yOg3KqEgApH8D9YV0Bkrpr9T4j1pbsfmr3CCeQPV2vwluBTqy5S1RBrvQyfqpaqCJ6g399reoW7Te6Q5Xyq25ofviiLvDrl5qsgdUlVuk+aWZ2ulxZP13sBYE6uCQAB8orgOstqUVykvOaJPc426WuGYX5j/KrI2cKVaTwGpe4FcSZ2OY6+r+BFrVWhd3EZ5Tog8eaXKsVPlGKoNtb9jYHR5XJYVh/Sccnmge0pkwWkvSLbrGtY+EKGsowa1LpmQFcRjA6PN5W2Fk0cV3yLZesvJZ0RUFHT/CREUM08/uPeI6r5ded+XhH68OK0oFtPJXXPHGt+oMfa+7bcf2698b5c8hyoDndtlkVIdGGl2jj01eePCycFg3xd2HVAwbu+Od37lgM4fk1y7X31wb6M5W9veWa7eXhn0hyuDo4/PH98vi5b2qzIMEO8R+nt2Pbz5xs/vyCWQSyCXQC6Bq0oC6774rqra5IXNJZBLIJfA5ZXASqKCzYAREuaqiM0KACvAOwlwAnARgIfzbKDZQAF6AARBCmQBfnNRZNqf5GfAyXqAJ9LhWeY/FlC17aq3F10kl0BxV0E4AyMdeCZABIAJ5aT8AMGYbxuwDOgCkMJ1gNyAMWh2Abagsc2mGAKE5/C+MeLGSJcsycCGnMNInTPWH2cIHMA06kh++Bhns5cFvrPgsoH/yAfShOtwrQEgS1kpy3P98kLMcJ0RGVybLZuRB5anWU+YJjB/W7mNKDDSI0tQkI8RHfZp2vD9aqflyPoszloa2DUmm6zc7LfsOb5bn7Iy0laAh4BqbFBNptKu859z7ee3sPF2wSjX0760J/Knr5DXxThSbdd+RtTV5Ml3tJKNJAH8tL5CWSCfGBsAg4A1U5my0R8gxSjn80o8A2CU/kt8B/ou58mfcYVfZz7JD3nSv8xtFn0cMCdVI4cHXMtNFGSFrCkaeuLrvAERFiOuJ0cRJfW448mC3Dwl6qee3EMNiWTxXEfWFwelwUl8isMaDc/qvn1qKPr1RsgKirTRA9kxRiAOGTNoaP+t0g8qrQykmc3zn+gPEuDy+0WAfEokCuRDV3X9RD8v4hhAXqw8iGfwLsSm9LSun74CgbB0foz9atj1JqttN+adLr6t5weTdUVJVx8ojw1Uy1Iud6XADwaKgddUC0sTXZRUkhyNnXdc7Sfg01WWW92BcimIb96lUBgvuOraaPu8bNet4+ee55prOptrAOxwGwaYDjvRB9IVzOD4E27yr//F8omv/zcDimPhTr71F93OD36vSDjjztNqMH5wZcR7gnfWx5Vs7uFZgEyMR8Ynh83VG3lXvWxyupCMVyFUjLmx9286b6gNmGNtnmM+AmQjODikr1lA/Ya+37yBcmCJ+C1KzGHMWbQPRBDvYt5nyJ0G2QxB6HU6vUIcxZqrPL9UkIMoWX2FUTItPe/R1CrM+W3pezc1A9YLfhKBw8olVFmw5YwIgF6nE5ZEbIi08H2IAgVr38zzN1DtzV0iS4/g5PRSOQzjIQ3Q0TAOh0WwjIptkYZ8nIh0ScoKFi5AVa6tNL8nXlOEzWIvjGi73hVubWHu/Gh/xhRrGN5tJNZjKBSsdTDW6G+sMbCwhJhO630FztGba/gLv9rWS8St+bk0G50py/auqBFWHUo+WxkMvGNPjdWXZ0caivtQk0rHDsVr0HIp7ogU2KF4DN32Qln/FRflOmlG5yAeol67cFDhp7OEBfPfNoH4xJCQy7WE9UciywQtt4mVESUKgj0nd0375X6p0Fooy3Iha1B83kryLsZ6EjdSrIsaGFuLBIjq48tBqdKbnj85WFM56wqovaRntUu1bknBsu9QXelHWB3Tt5hLGL/M0fMq53aRGYMDw81FkRLML6NyE9VUeUtyITW89eaTT7Xmqqp4EOp37EffqJqVRTzsPvrU5NSEYmKUBzrb/EK8l+eJhEmGb1gIdr76qDv42PZbeu3Kt3VjL/7CH9313yWvkwrcPaG8WeOpLLivSkoSqlxUea9CCSujCGbrQuJXXNb55sK7XX5nLoFcArkEcglsVgI5YbFZieXX5xLIJZBLYIUEMi6fDKxmbjXtR4BfIzIAGyAoAIvYkbABtUDUnAM4t+DQbGpIAB6cB5wAmOA+QEgDKQx0xdDCfPKfAwatsLwwl0wAVWeQp2im4IKG3NS0AajRtGITk25e+uUlP7P+AADmPjYYPI86mYsnykrZ2OSQPxsMNtfUyYCqLNFgm44s2G/atzyD+829iBE6lJjrzUrA/k6r0j8AjiApkNsPKAH2oAHO8wDTyBM5IlMrgwFMRgrYp+VpRAPPNu381erC9SZ/A44NwOO3LJCVfUbW7J/zRpZwj1lpnNWmz+Rj5eM32sF2uhYfxH6nH7KJBrj/dSXamb8BPPa5yp6OW35SMYj3Wt2QP3mYGy/L57yfq7h8svpa+RkX1JN+Qr8wcgHZ8hvlsWCW/M1Gn99oO3wdI0fGFdcZoYLbA2RKffgNAJVy8xwsbKaUHlYyTXKuszpC3FAGQEFznUX/PRuoF3dsq5EWqWXFFuVZcHfo89UaqV+jVh9XS4n4c8PJkiuIvKjqr0HVoB2flrukloJkb1Gdiu4pAd8AuTwz2YBlhS67oMNACEhE6oWFBOeIOfETa+QIeE37L4i0eBTSQt9T6wkl5qTfV/reVe7/eZ1DSx9bjz+SjNqXGhDrW5msLJq58SnF/kC17W2Z7HhjjRn/rsXTnfEtsRfuFmo06gfFthSyS8XAb4VhVK9VS12Buh2ZY+iUX5dLqKE4StrSMBfqE6REk851BNhGAmwvOwC/joY2/d9IQtqQcTClBGj+S0ov0vj3wrZrfOXDAyIsUnku3fQO1xva4RTfgj8ByQj6Tn9inDLfMg4hyXiPnNW6Vx+w2CurdJlr71S/z6+sM6QfRIMpH+ACihgXjLXvXEcKtBHp65UgXP+TEgAlfRAyknchigYbtXSIcW9WKhWwlJgOPG9ERMV03O2VZGHU0/eCLBTU9eOmXnCR3EeV4zDpidXQczzB/7G/3Oo1FLBbnv6LzNPnMFiXukUhTA4cnauKgBgRYSGSItqtcu9UrI3JZrtbF0ExUwgEvCpOh/TnpxW3Y6lU8p9vdZLjGsvNMEp96huhdqmLf77nsbawPfqUvqNgALFIP+AdjkJINiYR+axcs3COd9zvKf2hEuuptL9coRZwl1L2yJc58Nx5TxKsi4Me2pZsE8U115yv15Zma3LW5BqyMEglLJB+B0RDfbRZas5XxkVWeNXBdlOBpT9VKXbSteUK11AHdL0AfEVOqneqhWIUKu5FQ66V0pgZUVfWfp3gRKEczbSXSq8s1uSNLQxk6WG6MC8Si1kEm3tM3rm8ox8TaXJDY3KxNrpjbr+edVAWDU+LPBhpTCwVCpXeolw8TWr1jJKHubdjDqGf8TDWwygbsW4+petOibzg3GjgRQuqf2rls+OOo7XWQuU3jjwpEUUecxiu/zSNJNOyDnmFyAezZKyJrFhIIr+ue4PacMsT4TEmOW1VLJARyXKbLFYgXVBqOrPfkMVXUKqyR5qVOygFO0+yffyPdT61I82Dbl/KoZI/K5dALoFcApdXAjlhcXnlnz89l0AugWtLAqYVb9YJbCDZVADqmGslQOXblNjkW5BaAFM2IZxjXkZrio2PaaYC0AI6AlKw2QB4xPoC4Mk087kfoN6CSJ9PA8k2tebWQq6ghlXuKHT+AOUA3Oc5bBQoM5sPQGDyZfPC32yQzI0VmwvqwcYHEPp1SmxCkAWbHzaElA2QOAvC68+z8SD4zsEm0kAXysJ37uU8WquUi3KgEWaugwzoN/IAKw/IDZ4NSItMCGRKeThPWQFf7W+IF3O9ZcRSlrSgXPxtli1ZS4msGtxKiwjyMs1bAAbbfXI/v5mLB2RiRAN1ow8AxuP+Y4qH95+ftergOtonS6JQxuw73axCrC48E5mCNpLvTqX9SgAgWNhUXbQkUKpAm3OvAfgm135Rzv9hxJhAfpOFydiICuRl44C+SxsCblJfykn5jERA+w/XKfQpNrTIEE1liz/CmDD3KxAS9Ek0xBkXuL2wYI636jsyRp48j76A3OhPjDP6L/2JvkKZjGA0N2jmguxsxfH7L5Ki5I0KRPLdPd64gKSye7NaLlLqqJcN+RPpOAXme1o04uNq4Y8lofus13VH4gOuU/jJTWlEn332BX5Btsj5c0qMAeqGpi3ywipitcOIvkAkAPJdUjBuQBGAafor/fQfrnLje3SONgPQfqjvHuqSgPmrkBX0XcYtc8SQ4gXLRYZ89btyoeOGRhOvXK0XFrcvuKHJQmnYr5fLUSdMKkvNzrBAWhe249JyKxwuFf2gVinOVstBRyBoo9ONBiuloKBKtURwNBXMNxRoaqQcn6vOvSI1LrD5Lvg26k+fZ/wBVjKGmE8hFXAp8//25XOeB8hx1uIxVzn2mOuNTLmoMiQri1/4mx1//IPMIcyhWO0wXhg/jFvOnSXNLzVZdcFSunQ3IhuLm8O8whz0lBKB73lf/bQSCgxrHW/QjyTuZR3wi0rM5Vh20A6076r9zyxE+oG3OyIcZiMvHpJr/iTwAqwtSpq7K74+pddcEJg6ISsKaVG7Nh72sbBQn5dNhteWzQV+pPykHRb/4pMsTS7fMb/YDjrdsNbq9CZUp3GRjTuUbhSzMpjEAjw9b0DExFYRF41CUDgpDvqo3lVxpRy0ej2pmheCqN3pMSdulPB5OStrRAXjaocS70tcWvI+ZO5+xxoP36ffUECwY7++APL+lRL9DItTSORcO/3Me4F3P+vzFw518Dj0FGTaLbYXg4f9YuUuxXioQzBETS03ZCUhywUnt0q9ke1zxcZWf0Buj4g/QRyIWHEcFk/tG/+CyIhXSxWB9QtWFdVKozVXKMTDIg0GaoPtBQW07pZqhVJnqdRSQOvZ9lLl+VLcPaS4EqPFanis1yzOibA4X1vbOo/1sB2snZ5QxLtnVJYbRUz0FEi7M7hl8bMiVm4fGFueErGi4OEJ6yfuZy3F/fQ3ZMA51kbmDpT3N+tM+twEddNnqqgkd061PfccfGDm0MgnFLtCcbq8j+s87rAe7zRL9ePPTrR3333wad0zqmuHZWDhSR6eLDC0cEoOqRx7RGyYhRCuWnk3US6Zr3iy8HBzUdhbkqnjwIqFA/um+5SwioGgva6I8HP6af5HLoFcArkEriMJ5ITFddTYeVVzCeQSeNkkYAC0ubgBGAIkAzxnkc9mmA0FGl1sAFisG+Bj7p9YsAOgsmngOyAEpAWLcw6ADEAhzvOdDQUbWoBIwA/yNTCS600bf2WlARuNUOHZ2p3NyXnNcW0v3kX5AVSmlPhOAgAGHKZMaFhTL/IwggIyg00OGxoAavJk04wMsmD5yu/ZMiI/IyvYSAGykR/143k829xrsYliowJ4yjsM4J5P8qf+oIJs3CkjwBx5USdc4aTaYv1y8jzb8JhFCdcasZDdK9l37jEXXeRFXU1j1uSdrQsAEuWjfcxSRF9f9AzqhpwBFSgT8vuwEprwtC8ujwBTTPbkYVYJK60x6G/Ug/MrSRLaiX5n5BGyooyqk7/gqrfe4FqILv3dNGepn7kf47c1DwFeNhYoA/dSf0Nqeb7JgX5DP6aN2dgjI57Jd0gvCAj6OAfXUF/GBpqB5MdY4iCPb1NifAFAkD99iL4KGQXZQV9ig8t4tHUPz8evPJttCDYO+gabd8BAyMJUDlguCeBKwSwsK3R2RJKdEhHxCi8W8CsEXDXtJdO6r+ym5R5qp2CBkqwsviwri096Fc0Bo+5JWVUc1m+dwrvXjVXRL87mPmQJsdZBf0hJGAH7aHozl6CtiLuZ1Vw8kde/VHqL0n9U+mj/fvoPhBBjBvBgNbc2tAft8x+U/kLpkmgvZ+uvOtIPGS+krbELdotHu0VNtTVMhNoEQ34vKU/5heJgr+ONCNdcKsj8YqnZHdegKQ/Wy3PdXlQKw7Aa+Di+8U/KJ37Si5LqwlJnXJk/J1IjHKgW/S1jdeZH+i19HSKIZ9Jf6KtGDBvhuGYjXYQfjaRh7DP+AHkYPwSXRUv7jUq8ZzZ2JMlvleb2v7G97c60nRXT4v7uA7/ya6XpZ9HUZs7iecyvzBFxTlKsK1Z7l/DJHESsGCZd5jusJ3BdyDzJ3PXeNXLj/frWfns+pk/izDCeGZvMf+clLvp5xorh0FUhurIeCl0gOiLxatJoxsWdznsFEReaqOK24t5KZ9rryoHNiFwsJbIuUqeOiwrUTTwLT7Fc/MvpUmlhuaNSuIFmKxyPkninrEe2yb3VhAaAHxQCgaDJmGLOdEVm1NqdqBpFUVEkRZE4NeVSIeyGkS9CskUdJJtVyVWRPOs27HoXbMBdm4HotD+J9x3vLeYV5tr1yCzWDf9VifHNeISoYN42xY0kH5/ntBIy5p1/9ujKEdqyVlzygDc5vjveEUfLisEQb5VVhFs4VZdFge9Gdsz1asPNoqwWEsgIEQQdWUT4AuFvEmFRlTXBvbJ0EFcWpOEXdM2dA0PtQ4Vqr0BU7cGti9OyQggVB2KbLA1Cl4SlYq27Q9+Xq6X2TNzzW3Ec8A7d7HGHyJUn5L7pIblimi3Xusne1+3fpeePiCgY1ifvKNatrKtYb/GeYj1ksXPseYwD1lN84oaTdxd9k3tZi9eL1d5tE7un98nF01Gtjni/pOsq1WHXgUd2xOM3znxYbqmeU33fEPUKY7KkGMbV3NiumUTkxTMydrpR8w1lsH2OPXtUpMVcoVxJCqWy8utKhmd5CaxpaTPGRE66bbZ35NfnEsglkEvgKpVATlhcpQ2XFzuXQC6BK04CLOhNmxXQ0wB2QHQW2ZjzA0IALLDoZ7HOdab9byA/GyizoGCDAVBkVheAhdwLCMWngVI8y9zgWLwB7lkNaOY6ykpelMt3cw8X3OjbCy5qmWsngFqAb/IFHN7f/45rHlzZcB2bHJ5v4DefBpLbb7apMMsFXXJeKwvuBeCjzgCrpvnGeXYslIONEyAZZUcjlWdCGpgmGOUyQoH7kT1gmmnLcz3XmOYx5aeeyIPv/GZBtLPAklkrWPmRMWCgXct5DrMs4F7KigYb+dOmWdLDrEa4h7JRZtoTTTPqZoQMQDp9BjlyHe3BtdSZMpuVC9/NesUsTsyqxQBMnoUs6G/kZbKgnwy7cEEWNqpOvEg5KQv5AagZ6cD9ax59ywqeh1yMtKM81kcoNxthZEI96SfIiE0xz7tXifpyjvJDGjCmzL2V/U1foA2m+nmQL3XCEgCwhk0wz6Q9qINppwLkQWiQHwnQlbJQjjMuCV7od7ZLpvwdXEN1f0SO3KuSh+/2ipCYkLLlTrUY/XVQZEQlqbuRZMZ1vTHVX3EqFIT7OEkt9ZBKczQlLvAoAay4yrEO4bD6TRd2lvaFlKHsEBf/XQkgO0uqWc5v0hf61zOl73ZPq4yxgDfuBxj9MSU0vAHT7EDdGqsWSCfmvH26HhC/e6nAsj5ZQZti5UI/2SXo9b2KQaF+4g2GrvZsOx7xltzY9qW4Vmn1yl67271BmuOJ3MPUBGR6xWXF5PaSSN9jP/Db8nU/2unJF47nlkRcdHRdUS51uoMDZV3tQer8YyUsD+hT1J0+SX+DJEOz+YSsMOi/WPrQz5DhORrd61lgrOPyyTSz6fP0bZ7PHPk2Jdr1xzNttN5X3k2MuwclgkcKC0cp70+duckrHvn2/9rd/ZtvhwxO+/Olatf1Cn2V/m5WF5DV9B3GlcWq4DvjckqJeQjALmvVR5X5mzmdxDz3f/TbhfmQvnc+YI95vq230rSXJIfUeeTSxcklVLInVj8XRRfJXdS8/m7LN9Sc3KKVNHMFslyQTYI7KcsLuWtxBZF6/qnZ5UtiQXW+9tXYVJG8ShjHY7KAmsDNjtw+jWvKnhBRsSjEuCjOOZaJiC/SYlJAaVljeEAkZKjP0OuF0yJikBdzYu8SB+Bm3NKGtC/vWtre1gPMJygrQKyvR1YgHpRbcNPGO5T6mNVTaiV4uYPan6/9LtN5xh3vBuYwCB1ieJ0JuK0zcuFUHJxoec253pOyeCiXa51CoRwONbYshoq7IO+BcSiXS5FIiuej0D81c1jLGrmKUlyHLUoyDkiWNGbSdaksMk5VhlptxY44pGtOJWGgdk4ain0xq3VCS/cPBGHwql6rOLk0PXBYlgh3iQS5ELF0dd92kSWs0WdFUAyIvOBdxBzAnoL3Au8dlGCYS+gXrAlZK9NneD89r4QSC+dYR/HJe4y1wtf2r3lA78YtCsY9c+TLW0/IEoQ9ypk1aOImFH9j9PGPvuLZe/7eo0/KmmIoKIY7yjW3UyRNY/FUvSJS55DGIGs+1ohZi6C+0pNXkSLBvFxDfdUvtm6V2WNWFtxHe13WOedCGie/J5dALoFcArkELkwCOWFxYXLL78olkEsgl8BKCQAUsWhndW2AL4t9095nEwGYCknAJgEwCQKA380sGxAXcJu/WcijucSinusBXgGR2LgCCLO4Z0PE+TSIX/867mcjZpr3q7k5AOgGFOaaguse6zq8QPROaAOz20y/KQObOfI2koMNDfUzTSvT1KXuFlOCjbcB9+Rhlhf6mh4rd2JZYgDZ8Ew0TsmbjTzJdix8B1RgI8WmC/kZUGcuHZANG3/KasA04CWbLtNcRObIhXLyecYc/cxzSOauycpLGa0u5I/cKSPa++RlR3YTxfuV38z6g/stH7PE4T7qC7BEO9NugLsAoABVaMJPKSHDLCEEaQO5sZo1iBEb1q+ypJH1PeSClp3Jr+WqNw27hc/La84w9yE/5EBdkfNGDyPQzljunOmvlN+0sGkDyAb6HuViEwxAQxvgooYxcUAJrWOAGoBw+jdgHprHbL7ZZAOW0r7mKuoT+m6EHWVmA00+jDmuQb60GWUBREdDj3oyVhhnWDwB9lAOI1ywELCNcdofAm3xFTh7RMTDlFpSY8Y969+gTXzZ3aWWEAQmS422SCQ5dlftAB9/W+cJrj3rf/OVoxHYj5nRFrCPjKgj8oRGQb7vUVp5IPt/oPQB3ZMC1XIPRbvgYuqXlIiHgaUGB2SFHT/flynz2McEuK/pduViAGoqH23FHITG+juUTkip9dvPlJ/hpyCnXjJaCqLHC/FiM3LBoEgJv+QF3TARUBJ7RREQXrcX1hr1stxSiMQIFeUijEYEiCYFqbDWKqWufOIX5DN/QKCu5qLkn6h70Ofo7xYIGbDQSAnGA30eKwfGNzI39z30UUg8J0IDmTKPMiek43YdEsPmUvpy9l1DO9IOzJOAnYyBlQfjJ3VZ0j/o+4wz3g3v73/fKl8nC9Wjjzzpd5dui0t18nKt7ffceur+n/v4ju//t7mW6yqCPd+pNfp3SnBrfJg1DnMc/fgDSsyFzPXMU3et8zgAxe9Xov/w3tmvBABprgnP3t53C4W7pzn16/2KUdFS31YA3TTQtli4YLvcQMndixuUgz9PJIYn44qOzi2WioUj1ap/rNl2p6ABlGlyiUH+s/X4g0/vKzA+BYC2FVy7qy/lYlBodMKer/LGbREsigbgRLwMiW6OvAB3VnFHwK6GdDQlR5gLIiS/5MduoSznmHL3tmFrwk00/cpLGbe0r63neAfSRvzNPIKbvh/eRP6/p2sBpFkjMIdAkJplp60FN5HddXMp623eFYD1qTVETxYWsVY+hXIy25gIB4uVhadlNaA1izciN1DJwEirLIudRQWdXhQZUI0j75lDX9q+T4G29w5NLh5dnq1OyZrAEwlx1v+fiImktVBtRZVgUC6UNMqipcGJ5Wq53tXzikMiOKqsOnTPRLxUnlAcmXnle66rqo01ySk5gmqfPjB6i2JofH7X3YdOi1y5vX8r6yL6HGssc/vEWpoECcB6m74CSUYf5H3Fupm5hDmEe/ibuQp5zSgmxWtvev3zTzz3ud0HVP8ljUEsgl+nK5Yknx1PfeLmz9/xzq/MiLy5XxPbV1uLlWTuWGOw2yqx3kLpir0M70Y70vUsfKPyKnh+cCtTkgxYsoG3GSO8L1nP5aRFRnj511wCuQRyCVyrEsgJi2u1ZfN65RLIJXApJWAbUAPuAXnZ+KLhy+IfMBSQCgCJxT6a82wkWKwDTgDo4cKGRThALXMzYDILcoBT07hn82AupgAbuZ9NF3nbBokFvWnkm+Z9dmFvIJcB9tqyjUq7vlx2cozQf7Zt2skfsNdcGwHCUVaAdDbV1Nc2Qmxo1tpAGFjP8809CvVEe5eDzTbnzc3TI/oO0MaGkjqRqDvnTJb9W8+SBoB9yB4wjs2VATXUJ2slwWYeYJFNIZs0ACHKZaQC15sm60qChfPkCyBqJEaWtLAyWV48lzY2UslIBn4H/E1dqSiZ5QSgJhtIymSutsx6AvmYxQZ1NXKIZ9rzkJPJmPNGHkFCcA95AdQbqYastjpf9veQFVLLswro08iulTLIXHLma9+6AtmYiyzqw8aSZ3HOCAI+OQ9BQ99mfACc0o8oE+3Cb2xm+QTMQSsdmZMPbQ8ZwLWAM/yOHPnNXJF7/e0AACAASURBVENRJABb8qR9kSNjiLIgb9qDDTmufADjqSeWAZSNRJ9HjrTZcdecXQ5//58Wkv1u1KvLrU5drqDKIjmSdMw+pBYZUq8lmOVn5AYqlh7/UT3xI/r8is43sUqgQFfa0S/XskB+xhrjkL4A2M3cs/L4ZZ14q9I/V3pc4GtbACv9iZgWaN8jawiClce/1Im/7OcPkAbZ9pLksUZgbdqOfkP/AryF+HuVOq9YWNzbyNdNLK83fvTqRbf9ielo6thiXBvpeUHNL/rzwmVb0tVWoNBE7mK8srTHJ+UuptluhVLY9gYGKsVlaZsLF5Wzj6DQlNPuWGQH9f68En3rD5V+Vwkwhv6HfACA+m7X0rmN/ocmPBqu9EnGO32Yvsx7geu5jr/Pd9hcxXV8t9hB1Jv8cX/3I0opEXKeI0tW0Ca4/aKdGI/0a8qcWjJ1R/cuxMXqr+p7SljIZcevnnrzzwkk/be8e/Lj4krArPOYk8z9GmDifiX62M+s87jv0e+k/12JNmaew098T+O1l41fIJIhlhukpoi341GUdIpFbzEIghlxdBPiIUqJ5w2pqzdksVARhzetV8MpuaNXmRK5rPEWZNmwpN8vibu389V5bLjmREwUojCqNltBTZYSqnMyIfBZRlBJx3Wjssyi8G5Vl1VIWy+4luaCokgOEZWuKnKmh8s/WZSEvW4aYJj3yssFhGaJCtqSNQSfpgQBmPx/rtG+uP5ivrCDsv63fmKsMvbNgosxTR9aTWHl4vbYqzc33hcQyMy5qaY/ZIVcHLmZw0GzvRhNy+3Rq9V37lR/L7QXKwdELpSqjXYnGF9OBNI/IfdGI6M7Zr9DBJgna4tByAoB8+J5bZmX5relOVttaZWQiPzADVRQKIWDiu+gsSXTpVqvIOuDBVFrDXpe6prtzHokS/6vJWXaHeJBPqtkwyE3VfXxpR+QpcUn9PcBvSFYq2O9Sr82a2z6R2ohp8S7BgUc9iu8N219zJqLtRPlYc1F/+QeyvVpES8jkzed3rl0ut499vSWvao/8xR9+SCeQU/uG9/92Q+89jNTdx/6O1lWLJ54dmKL5HOHyBj2EW/uyzy7FqAsLb1Wnwk7y8OKmjOupFO2tE3Xcvzxco7RteSc/5ZLIJdALoFcApdBAjlhcRmEnj8yl0AugatTAtrYrlbwLJhrgK35/Qf0hJgAkGLlzZwLoMZGid+MNADYQkMOQgOQCYfJnDOyAJKDvAEg0ILlIE+ugbhgE8Hml4W8uXpiA7NagdmMmNUCu6q2tOtrLlxsSbGSMgISG3BL/hwPKOFaBFCT+6kfzzFw2kBxrjViIktQrCRJyJ8yc/CdjRHa2oD0lIH6spHnGnPhhCyoP5snNlFmuQDIYC6hLD+AQDZmbJ4A3qgv+QAIAiaaxQjX8SwjSrjfNLe4P7tbMpCQT8rAJs/a1K7jfqtrVvamRWZyop3MDQRAg5EHbFIhWqyOAI9YA7CRtPKQhxEx1A2ZrUZIsbnLRvmlXtSbjSp9kHvICxkvuqTbdr6K1N5Hv+Re5GuWHdy33mEWRlxr2qOmyUcbsRFmo4u2nvVnc4NBH8D6AjIMAgHZIBOICA7GBGWivbiGfpi6PVBCNmzIycvcofFcyAhzR0VejEPTGjQ3V+RFPhAYEIVmUWFgMfWP4mc/4yfPf3KLNxLc6k1EU2rhAfXa7RrBe/Sda6qKZzGob1+rkr9f5/7aKwoIKZwliPrVuGI/GBsAFvQ7yFXmIRvb2UKj4Y3rmYMiDU6J8EArnLZFXj+pBDBqRF/2PoDu9ykBeNAW1k4XSyD0N/o6cyLam8wTZwOKC5RM6QqOdjJ4sBUP7ujG0mQtbjkeuMa+MKpsF/Aq1/fxkpBN+fv2C12ATrm8EXMhJc9Yvj/iqvxd+MJhlqWN3oz8uOPjGCSJ5zwveHtfZtQLMAbi5zN9eZqLNsY1YwuSzuYS+h1/MybNbR2fyGitg/HC3AbhaiQ58wTff1oJMGgjB+QK87i5kKGMjE/mQ8YaYzLa8f3/Jv7iof+N/O2gn9wji5C/1edGLEHS+3Q9H4Y+vWieXM8l1kYqdI1dg2zpI7y3mNN+XelBpbuVfmGduv5r/f4Fpf1KEJIfVJrBnZtIC7NYTLMQ8dAqFgNZEkUtNYqsD9yYenrgRcluEXeK/eBEZHihi/22gP5OtxOe6PXiRRF6IjvOIbgvufghLBab3YFmMx6p10pDYilkBeJV5K5tIemEgfDbhty4eaVSUVRj3JA1hV9QsHGdn1Vdu8JDezK/qGh2GJCws5aVF6UuacyjFywhyZ91DcAu5C/zBkAwBOF3Kd2/xkN5T5FwEwa4Trv+D6W/UmLuTl0XKvGeT61eLkoFrt1MkBFrZI7sOim1tFg67UetBb01EleXhcCAH7imiIp9IhhuloXFqD5nFdhlW7ESvkIukEpzx4barYVKbeGklgHhC2QFmQPeC8yflyukgkgOglS3/ELlxmIpkhFB4oJC1OoslUVWpM/j4B3Ke2Gjh+0NdL3n2ovlryi/YbmX2lUZ7HxSxAV9jf7Bu4V3Nesq+gzfeVeaIhLvAd5hrKvIk/UR7wSuY43A+5VrmP/5flRusrxddx3CsqM0c3DkiyJwFlW/VOFEJM47lmdqdzz5sVt5p1AzlI14Z/H8P1Cy/Y5Z5NraeqsEI8d0ipQjE6jMvot3FW21rgLNRgWXX5dLIJdALoFcAle+BHLC4spvo7yEuQRyCVwhEpCW4Wol0Xo6DTTMYYSFza3sXEhorWKVACj/zUqAalwDgIVrHjYIAKws6rkGooBFPiAv4CwLew4W+3uU0KJj4wBoBVEBmMRmhIU/GwvAfX5bTUvXtO8zwKL2buHpyC198bir38rvbGIoNyAJ4Ni39stEfhAkbBooH5s+AOPsYbLgNwMAAMDMRZERAtSVawBTkAGbcAO6zVSdOrFhohw8B5mZJQLPJA9+JxlxYW4R2IQhUwNUp/TdiCM2/YCvWe0uQJzV3CjxHCMkKJ/VBWDegAE+7d6VsjAXU5w3oBIwmHbFkoJ6G3lAW0JC8Df5QywAaLCJBLTnfiM6yNfAT3sG95lbI7OoIB/O8TeyAwCjHbkHOUOOfdq1D+xx0VLRLT6yUvvd8svW63zfTR7InbajDyIX2idrKcPzucaAM74zFiAUbFxwL/nRn9k4s1k1bXLGD2MC+ZhGPeWkrQH3+J3z1JexQp3ZRNN+pp3H9VgHAPhQRsB2xiFjjPFHXwmT+YN+/MAvb/NKp+70xuM7/C0ab5Ebimfco3INtTctoUaOcqZ+T8qRw2dV2wOqRbvvekmnr+yjb2mBiyhIU4BO5IKLLrT0swey+c99ef2RrmeeCftxLZDzjyl9n9KUEnMR1xtg/7P6DoBKGzIXpn7VL4JkyI++wlhAixT3T8y3WDCkB2QFpIWgIQC9sdgVjwoYWpDXjtnYq48pbrackpflj1+sXTecwde9HHxNCsgsyENMOXD+snpIr9nqDUhXuyaNdPzO9Hzf64rQwBqFMWwEAuWhV9D3strnNi/ap82NZiXB/fR1xkSyErzvA5/0U65HpsiOv+nXb1T6biXcndm7Yi3RMsd8SOlPlRgHECaQdWYZyDkCaGfnAtqX+cqsbyBGPqn0IndD2QeLpMjW2+Y/I7O51N4Dnq7l+3n7xHVKaCAP+gVtwzuDOZtYPbwzeS+znjjfwXggAYbzDgUYf059CUuntto36rty6snSIlQQbQJwy3rI6xW94IuK99CUexrpinvTLHEU5KKl/06JyDsuC4ymgrd0Cdy9xvNf9p/mF9ue3DglzXZYKRT86kC15C80O8PqaLNBwTslYqUiwoWlW1vWF+VEMTdEQcqqAh9/3oICcDcVf8jXYCQWDePpogUQ749Z3rum1Q5Rwbz6TUpYWU0pQVqsd2D59BdKvAOZX2l7yMK/UWIsM681V4zX9fK8rn9/+MHfTV5z3/ebpSzjirXH2aOz7I0dfqJ6vDHpdlSHusdlDSHSIh71gmRO1hPj7aXyuNwuQUYk88cahZPPjeNm7FHFoXgz24QVuk3PyjJjbxJXmor3MKjrKstyVKb4Dq5YDkUwVORayl95D+sh1vVZ4oL1ja0zs66Uzpab54oc2SG3UM0o8hsj2+eHVG7cyrFupP8wZzMPs9ZkD0H+KL3QT1kz8X7hncLBd+7jncK6irUT37k/tVolzpMsRA4qnsWAYnrccPyZiWOSy6tF2tzUD6rN+jVrKU1f5R2XXROeu7FSRG7FsIg9mUDx5s68Eqgz62DWZtTlYqwf+lXNP3IJ5BLIJZBL4EqVQE5YXKktk5crl0AugatNAqYNyeKbRTnEAhrlAA1oxrHYBxj6fSU2CGiF71ZC446NAvexseU62zyRD+dTEEsJ6wo2LV9UAnBn84A2L0AS1xpIaxpjAN1NXB5ox26Le84BJDL/nyEIlh9vue0/WndD90zpb7SfABO5hg0dZQb8Z1NnliPUi2ezceDIujzKgve2EWGTxfO5jnJavAieD7BIuXkuCdkA9AECsllik2IbJ9PAMlCQZ1NGqwubGL5TPu5D7vv7+VMHNjtslJAdzwAIoizkZ2pxbBRpA37n+bZBtN/5Owvkca/VLwvEUbbs31mwjvwpJ8C6uYOgjdkoUmazLKF8WBzQR8iLa8yyxMpMXllrHcrJfeYTm3Jw2N/Il/JyDW1IPZVnUnG9hZorTnCdkRxGQGxUI57y0cb0FfoyJBP1o4/yPNqEccHv9GPOA+JAkJlWt1kdIQOrK3kA1FFX2g5ZQJzR/7jOyDHa0iyE9DXtrzzPrAeQExtowFnu4Txlpm+YViF/M34G5GC6F3/8Vxpe4dBrpC94kyRVSGZ1vX4RKHFQEo1Uy7Z61MNeSRvo2B3wGmfyvFrICoSUOWh7gAnki8ypC/LjACQzMPzn9J12BgiBfEjnGSVcItEugHAAqVkQiHOMddqR5zDWN+UeaoUrKJtb6GcG2vO8c8gKqxvuoFSpsu9Fn5+Jdj85G9wy03ODca8b1np+2a9W5Nle3rykbV76/9l7EzjLzrLO/9x9qb2r13RIVzaSsIQgBofNhEURwWVwFEeD4vIfBpX5j/8ZVNzB7S/z1z8uM6LIMCqIjKKIAoJGEsKSECAEQpZOp1O9d9det+5+tvl9T92ncvqmqru603u959Nv31vnnvOe933Ouz2/3/M8ryzHC8V8LipWcjEbp4ZhkCmXCy0BuL4A3Vy5lGuIuGjl87kZtQPCiQAm4sFD++ofH1aK0APcbRy2MYR+wdFMb6qd+m793MAaxgwjjOnLgJ9vsoec5PMj+p3xBbKZd0u75z3QFykPJMVaIBB973eU/rj3DOYvwC6IjFWPHllh4yZjKfLhkz5uSBRtgb85kjL00jqrdOlcdpI9XOLeHhf0NQhVvGM+qfSrSuwf8ysnkcQv6PdJJazyufdzPW+LhHDo7WnR1Z4US+oIHZF28kLwjsilaKCQywae4p8pbJT+xU0hq22Rdb76iRkfnLeX0NQQrYfXmx3/iMjDuXwuK8vuWNwLm2uz54bmHYWEUsGTtYv6rS8cNCcS4zLVcUwzv1/M5WeIpJOPI9rnU9qPI0UskhegLkYn1yhZ22dcxHNyvQdeNX+hxLhpnp0QT7QB5lHenwNu1yvN469j3GH8IqQf72jlEHfVnjuw/Rl7Pl8cGRjr5rdePT0mb4pSZaR1SF4RCgdVqM4dGo20J0M2aBdaIgmmFeroukK1q3BQGS/s5uUdsEJCDOq7NsTOEqps+YhyXlueGPK6SDwwVnHepl33e7Ye5wmydpUzQ3h7RPs2PbhlYi7cPDHLeodx3sI7MeegexjxzTxgHhT0E+Zyns/8ztqThFEJeoetAVgvsT4bzeajpjYj114wMujIRVsbcwOl+cMjeREXQ6rXhK5hfmYtiLzx2uNZlMU8pY+rCv02aDcLoZx+Y3lYpI5JfcfowZEVa79894uTgJOAk8AlJwFHWFxyr9RVyEnASeA8SMCsIFHgWdwDJAHCoxBgzYgCwHksjVAEsEw2kAhFgL8Zj1FQUEQBwJL4GToArIizCwgPGIbiiuUVgBMHIVxQWs2SD8sp/uaZq1n9GyBkILvUiFbeq32x65W2z3uVq3kuCgbKMOA+VliAmCjJWC9TR8oM2MjvAJtm7WXeB3wa2GwWtADLKCgo7gZi8RvnUJ6oH4oM+RqpwiflJX+u5T4+zeqfv80yGUCNclN+5MM93D+hhNcKVvqEXELhMmBRX5P8sfinLoBp/E3ZKUfa0szIB1M5rX4GlpNX2prYrqOMBvxzjYUzoo1wPRaSAO9GBgHqUh6UTABBZGLP4Jn23WRhXjzkzbvhvXJYaCYDBi0kAO+OfLgWwoC29w1e5ekDXv1B7WVSMUCRPAx8TRM0veyf9JEGVm1/CPOc4DlonhAK1mZQkgHDAbhRfnkGSjXlAgyFXEK5pQzIh3fBvRz8Rt7IkvbJs6kncqM9cCA/ZECaUKJf0W4og4VYeYG+f5MS7QVPC8oCoHtQZo+T8YEvPM1rPbglMxaOeX5hT7wULHrF+AUqaS72vUOZIfXtsrdL4Z8Oq2U+pjQjosIA6F4xLroP5Mj7wor7HUpY7f9HpbTlPgTTLyn9gVIgIgHvFEiaRQF2hEKi77y2r+b0Rdrz7yoBrn5MiWfR/tbTvvoFaVbLEBQvV3qpEn1oxbMifcNy5C7v8+1o+A/9uDraCMeGGmFpZ6FYLAsgybe7UYv9KWRm3ZYHRU7AZp19LGS1PdPpxn6pqF/UfgTU1mSJXVconFq5lBf4maWNUg/GeyMirT6RSIrTBRON4GQcQ/YQdcgPYI36mqdDv1xW+/v/7b0TgDn6Gn2PstInw/VYZlMPERB39WVOeDCILH5b2SC8R1RklhqdfKmYZ6wdkMyqkl1elvlDApDDoBslXkn5bLap3lsX0Gz766S93E5XduuRycV8DXLh/SF7xkwMFpjbflEJQqv/YExiXJ/oJdoTxBPeFnhVESYqAerlaZEQwIRW0ifhoCp6Z5pjMnJGiAwcjzSS8rt5aJxXWaqddcVQHGu1uo/rUwGgslvUXa9U+8qJxBjBfUKFL6tDFdQGmSOYMzcptE+nXMxNsj9HtxtQV+tzq9YnTSj2XWBzH/kCKjO3czAXYXAAKc9c1e+xdiK50R/+hnekhFcG6z3e9WeU+I2+m15XnNd3cJE+nPUABgx4q7AWWCbnxUIr2t9LQz+zefHYgMKGFa4qDXbC0R2LRW0Y3c0XglntybD98IPbGyIciiIcWGM8U3s6RJsuX9C9kadwTIcUmikX+vmcNtN+SNeMCLznOvM4hKiYlSmRGf30i9DW1Lxn+hrrGebKk5JdCfmhTeXlBbLw9dufvvuGlz76ldHttR2Fiv9toka2yNvwIdkv3d+rL2sp1sbM6damGFtIzDfm2Up50CkoA2WGgEhCdyqvm+QtcsPI9qWR6kh7pjFf/czSzEBZXiVXaF8Oxgz6B/kx99Ce0YWYv5gb+g8IUZE+8oZKKmJL6pXLkANrRFvzrZKFO+Uk4CTgJOAkcClJwBEWl9LbdHVxEnASON8SYIVtFv8GvgLeQjKwSAdM4xOFE+WIhT+ANZaSAK8AheSB0otlHh4VLPQBagFTDYxGkUDJQGkgtABKBNeRNweAIeP7ata+LPRRmnguZIHMwMK8V71G1y6rOr38eCbAllnvv07fUV5QFig/v5OXWcTzXAPUDcxH0eJZKPIGknMO5Yd8LQyTWZJxHUC0kSmA1P1ai1nn9qq6skEteQDgmFU916GMEXIKkA/Qxlzg03nyLO4xcIz7eIe8GwPPVuzienWh3NQ9AW2UACZMszKCwZQxAzMoL7LlWcid87xvysR5s0Amv3R5LB97N8jIQkDxnfuMlOAZlAnFkHPI3AgK8k0UzF69yANghfez32s+NKB9LLZ5nWPkyTs2IoeyPElr5EF9h5FURqjwHCPN+G2yVxbyph2heCI33hFgDn8DHnDf9UqEqqJtQ/hZaDDy4X4LN0U+1Jf3RJvE+o4+Rp0pt7Ur6m1eHtxPueiX/E77gKSgD5EH8lgKP/3uKDOcCb3c+EA8JRV/rHtldrNinXfVb9vaGPKIOsustyd3vcInbU7q4wuwP84cUOcu1gP5QPIBxiPTb1HC4yl9QIxyHhCcsWhKxEWr+1eJbAFDCFH0dqVXKfGOjGwij7cpAbr/phJEKOMj/eZkALUBirxb+g2gB4QF7QJAf9UwGcr2Y4ru9O52NDR4X+M7dmcKo9vbhfFRRbMf04g3IsCyJSCzlMvmO7LFbgqAEbkSN0rlfEWAp9fxA23qG0UCNw8EYXxE187n83nIC55Le2EjXPoS8vhArx7I598IvEd+9wrwRy7rPei3yIv6UD8s6BnbabsAVmmygrbHtf3recYA5g8AWt4lBBSkEWWmj0FUnEze/eUFGAd0fXfvB7w7/kFphaQzsqLR6ha0L8IQVuxiesYD9gkIovmOH28RaDYk8LumvULa8lbR7ZkjgHmQQPrDPC6ScfQpED7rlfXFfJ0RY7QtQFebTyAYIfDsYPxLHy/RHxC1P6WEMcQgG3In7/GOm/Gy6Yq4ME+9jrwT1O9W1gbkk8xFvXBS51V+O7YMRSIsMptHq+F8rX1EG21nRCSWRLhktA/NZrW/nPapoA7T6sKb1J8rAqTZhLtdKuRn6fu6Vh6o2cUoDow0W0+dbE6kATOfs15AzkYMMXbiVUbfxRhjvcfHdeGkEv2XdSEeAMyR9A3GSfpzer5fb77uuj4JKCxUpLBQyJd1CN4E5k3oReyfEHSvCtpeW5tKj2nviTkB8Y8Xy35bwm/OHxzdKkJgh7wpFClNIcVy2p1+S7277ZrpmsD7UCGR6tp0uqG9HeLWYnnP4rHhvSIRDqkXXSGigvU973Q9xg2M62bMxLy3rkPPKBEHUSGqtu/53JWPbr9uKhjdvvjQ0JY6m4iz91ZLe2fI42hlCqAstC3matZC6BCUEz2B9ZitsRhraOs2n9NO6TcF5ZfPDkbalcNriKgoaGPxh9nPQ2VhbQcxiiHKNyvRd+gn/etKxv6GbqiHgb+VIScJr/VEjelTPPcJY6t1ScNd5CTgJOAk4CRwMUvAERYX89tzZXcScBK40CRgC3CAS4AslEwsHgGdAABY3BuQCviEAgogi4UyoNeVvetZlKMscA4lwjwvWLujQJh1PfUHtIBYQIkw0A/gAsUDYKrfetkszVGYAMMpc+A1vh54uSHbK4F7uB/glzICSAKYAURSFwPozTuAepqlWJrEQAb8zTO5h3InYRcoePLcJ0gYK6fJcDUwjWtMWbHrUKAoN/kaYAPQh5KEAopMIXsgLbgHeVroLK4zDw6APCNYeLaRTChWJm/uR8Zm3WV1IQ8jbvo/+y3BLAQUsrF9KVDUAD1QEiFdUBCNtDAPDeZr8jIPEORn5ICFuwL4p7y0KerOe7PnWx14Pu0Q2aOkA6y2vIFnjmnj9by3eC91t2cja+TL+1vPQXlo1xZuy8JqWRgTFE7bm4M2w3uh3pSVcgPsID/kColA++Nd8V4hGHh3yIxy4SXBef4GLOZ+wvJwDwd14H2SF+XCi8K8LvhtUgm5AygbAYLsN3utWim767qi17x7S2aH9vXItnOK77Ddy8aP6smPyZ5yRk+7Pzvh1bS9JGW6WENA9UT1pA/aAO8Oa0jk+n8r/eMqF3+rzhEmgvb3z0p7ehv6BgJAAULZIwHCYjVLSoAL2uCvKPGOj+qeudVAdBEh1tfpM4yLkBW8ayyPGSMJs3Ki4/f9uPJQKxodbURji/PBc+ubitWBeisaaCsmlHwn4nKxsK1YFLYZxTMC2NVeMoPExg9zkXDOOGnTwk+m5HFxVGGhagodJcvbMBgeKAHuQLowLjIGUj7Gb/rejyvh3fDHAvIJ7UKbTULw2NG3LwP1pG1TT6yyaadYvn6P0sQaFaT9pw/KwnzCWPBhJUgLvidzwWmQFOm86Zt/ofRzShBYP6rE+4OcTx8ZyUyRhFR+gXkCkcvtrryUYm84jKNtquRVxBbKxoIEg0xHe4U8LHJjTla180Kojun3hv426/FTJVXWENMlfZr3wnwFMYXc6LdvUaJNfsMaNaeN/YbSpBJ9nE/G07b6Ybt02802H0NeZC4EcmK1ekBofezLh+KBapF9KWbU1tg4vCwXqSu01Yz22fC0P01mQKTEwbAl94uMV5XnFJuHy6EqqssDqCa6oqBGFmkcWC9pSptEfvRz+ihrPOYwwuNNKD1fCW/UtFfaiRogcxBrKTyYICkYA5inmR+ZX3i3Ccmo5PrDiSR56r8hUw7m/pUjg1tOJjOgVjIQaZZq1yqbko2xMbbIeJPyjCgIiF/xluBGEd1L1dHWpMiLtkJGFbZcObuQK4bHBNrH2lNiWmGjPlCfq1Zqx4Y2K0QUxC9r0vUezHl2fFFf8NbuDxnVn9erVcYXNBcqj+277/KHF7YP79d+E/PDW5auD4PcUe2f8Wh1pPVF7T1xd3Ws+ULdTJtjLUW+rBExIKENMtfS1mmnNtcyPrCGM8MP1ojzkkGpUPJb41fMH67PVpuSw6hkRd+AQMXQinUs/Yz1aP8hb5XYC7rtKb/dvKpvw22utXCdHfYgWa/g3HVOAk4CTgJOAhe3BBxhcXG/P1d6JwEngQtDAmbxhvLDopqFPMAp5wEDAGVRBlA+AbgAibkWABeQAEUIYMrAKrPcx8MApYi/sQRjzCb0A4oDyg7nAaPIn+uMvOCc5dEPmJuVPfcARi97QARLvlfZhcfGp5RuVaIegGvkA5BMnlgLAvoCggHOoZCbtbq+Js/neQaym1JixAjXIJM0iM4zzNrKPBfSJEvaCiut5Bg4Tn7IEtmiEFEuwv7widIFaIMS9rgSir8RF9TfykK5kL0REHwnT5RYgDkjBrjOymAKE592Dhlx2B4QvT9XrpyUxgAAIABJREFUPuw6rKINWKfcvH/Khix45zyXc+YlY+VJW5ZRPv7mMGLJSA/aFffyPimLvRcjbFB+UUABSSATxr1wMe9lS5G3cBfXkigLbQOgpN9Ct79e7Goasft871rzrkCJ5RxkAfnxHswDhffDc7C8s9jM/GbtEtDNyA/qSTs0UAEZcS/14x1zHXXiubRNQFzqz3euow1AgHA/xBtgMiAr5TEvGsgr6rvohX4ls/0Zee+RP/e98OGtcTE4EC/GJeX4uDbdXlTrjfPfpHoUl0NzXKT7VajoJzysX3ERQNr3Kv3/PdnZjbQnwOuf6cm/KXLhqOTBu+ZdENrul5XwtFjteJlOMp4BsgOMfElgqe2XkoxfPYDd+gHvFaAGAIQQHj92kjpApEDebStna1/qBNdOibTQTrvDhVxTmwbnso8LpMxWywXCQA35QVRWpdWv4rJOD7fbflFeANP5Qu6RZIOLTFwrZL2DrY4/JUvtxaWOH27dNEibhcj9LqVPK9GGIGsop40Nb9J3EmD/zwhkpT+sHKozbdCIbPLjb8ZaSAtkOXGSetrP/6IvWGgzxyBXiIskxA8XnGSPhHU+Ihnr6Hd2fJ++/J6SAX+ZVtsviLAoY+Uu8kchtzJbJbvr9fe2xGTWi7GeZbRogBpr+BzUNQflvaIxOm4qIIgcMuJQYHLERtzOy2JZ1Cd5f5HaEe+a94MnDH0VoBFPTcDR1Q7ARvoo4zt96UNKEPyHlJeN3ZG8LuK3iHo7Q+1nve1s3dd9+zfsDD/98LQ/PFjqqsENdzp+UcRiq9Hyg3rTb8g76nL5iKj/ZqbVIXOKGaUNvTJZtbeFoOkvqknKwyderJQLHe2JkV5vJGXo7UvBV1ufsU5hvoAMop/zN3Mw6Wd78lxv+f9VF0Ic8VzmPvNAZBzkfZJ3sr68UOW/3opeoNchW9YQEO/LRxKSKNQyoC07hYD1bZWVTRxmmYdYexyHnXC5PBVqIic6+UK4RaGXBovV7pJaWUv7XbDWnxm9bHFA3hgZeVvUHr7z2rz2eLidzbf1m4H4PJn1o5FVa+EzzA+E4lvPQb/WXi6ZqsiSwYVDo4dUpq3zB0ZZAxejKLO7VO0uXnHToRsKlW45Xwrb+p0ysEZijGcdzRxk6zrWwlYuxhnTJVg38xtrrP0KjVW9+t88PrP7rqs/szQ9xPqTccbWcOYx8qR+RoXUF0v5YjnKFQqTQac5sbykTA7Wx8ybrJ2PI/3XIwh3jZOAk4CTgJPAxSsBR1hcvO/OldxJwEngwpIAK2uUCcgKIwL4hGhAQQA0RQFFId2rBKAHKIBy8O1KkAIADQB3kBdYvwM0odCQBwoVfwPaEfbGLO9QBlAeWNCjBLCoN0s8zvcTFvY3CgQKxzJAXRe21T4IeYLSDYgM2GHglFm92/MBh22jXQC6dIiiNBmhn5KD5xgQZ4oKnyhsZknLs8yLwIA+I4LSyo09i99Qrkyj4TzKJMAfeSJbQHGuQfFCySMfe56RIkYiUD6en1jMK31EifeGwpm2pENuVhfqRj7cRz6QAGlZ2e9GNJA3ckvCDinxvnn/kEDkw3lAR96vhc4CxDDCJG1VZiQG5/iOEse7p/3RRpC5gR3WDigbZTRAGWUUYJNQUNNe8+FtnvY7pNC9+63cqyqXvevSH9xrpA3tnAPZ8J5JvAezCjQrdIgJ5Ml7o90BAvEeIVPM88SsWSkPdSQv8jGLQK4zRRarcsAkwg9AhPAdAHdCCYKCdsEzIS+4j08S/XPACzpTcXupEH3hncVM7a5ipryobVm9xUwpc8QrxONqQZTzsN4U77F7iZIVqtrKYf2Ftgq49kPpH3vf36FP2tHvK31SpMUk4bEE9EEY/LES+1W8X2m10CgA+cgS76J7lT6rBNHEWLQ3eGcyTjImAYjQnwmJRNs6EVnBO/4TJfoV+UK4zL9v7l3URf0izApUr23ZNLA78MNBhXbqyup6RJFvtpfyOV8darpW72RFZmg/Xm86l815mZzXFYD+qHiLOVlnN3R/VySHycbIQ8Ls3KHEWP3XSvSFv1Gy4/X6EgiE/7XhBz986PK//iHuIw/6OGM+8wUAM+39F5Vo3yc7eC8QQrRt2jF1TYg0JeSUHjNOltd6fidPvEbe1rsYS/73KgH6ebsnZzyICsmqXC7mt1bK+evyhfxE148GG01/JAiDTfKeqGhj5O5yiPJMKHD5Osl9WOBUpJsqxUJ2vtnyHxDpEQpENhmvp2wb/Zo0eU8IMEhZyEAssn9eibms/zAy+j36wQB45j7uoV/SpmhPjJVnui2dsfdVb8qFZ7jSFdFVVzs60u74o+1OUGq2tHOv5lK1qSify4S+2mExH7fz2njb9+NjuvahUrlwUC4W891Au1j0eaRqDDNglrnH4v3bZtfMGXh4MV4xLr3yFCrEWMocZ7Jl/OT51neNADyFLN2lpyEBxhfGXdo23i14DSaERdDtaBJrVvOFkjwlSvQTW7uwHmKMpk8kaz+B9HhUxCIqxkRe0E5Y67CWZ13+iIiA4UwuvkkeGA8861sfnjy2Z/P/euyeiU+ISHixfv/OXn54SLH301rYDGMszz2pAYmusfCt6A+sNcvaS+NHaGMiMAbLw+2njYw3Gtose1QeIVtq00OtylD7s5WR9pzKyrxNG6cstHFbI6NrpEMbmu7BWpXEePOPIh38fFG7jLeKe0SKTPTKyzrM1pZrrSdF/SD6YCj0uxNRoGXhE4QFskYP4j0hH9c/JAR3OAk4CTgJbAQJOMJiI7xlV0cnASeBsyoBWe6RPyajy+D/8mIaYNUs8VBesHrnb8KCoAwAUKGsYNGIhRILfuLpo7gCtpoyRD6ADrI+TSyVAHMtnA/PBYRAOSFPFCruO46kUPnSQAPX4RmBYgygi0Lf9VqPV732fv7mWsoAYWHEAQoSycgYLNQBFwE0eBb1BTBLICgKlTqsLMw3RhLws5ER3Gvgus1Jdo/llS5/mmBAebJN+JALwDQgHzKxsvOsdOgmIwb4pO4W/gj5A0pwLXmwfwJyQtZm4U1e9jf3Uz4D9a2M3GvPNiDT5AIwicW3EUW8e94HzzRlGNd8QkzwHAul0y9Xe5bJCznQvsgL8GRCCVKJPPtlifzIF6IEggDlesbLj0kxzZa8sG5kG9fwvimrkRDUf82j52WBTM1K0EKgEfKH9m6eFJAVPJ+y0HapB78BSPNMIzeQMYAzCjdtjnpzPWQe5cS6lbJBAGIRSB639q5BfhAhtHMs//iOPCyeMufoV1xHIvzBobhVm40++95s9OAdo9mt+aPeUn7ay9SvyozLNL+iezPJPQfYYFqfl9ShOiWHCIf0gcyRIcA4QDVtGuCj/4CM4B0QzizqkRZYfQPYIKsfVPodpVtWuZf2QKLfAt68R3Juq3V8Jm5ovOzqnRYUUmJ552xAkVtPIvif0O+TSng+UH7aChsEewpvQzvwtMkuXgBLija+R+TEFQOVYlVAe0kBoMqFYm4ql89MFRXvfkhW2wr/FMhkW/tWZGfqjaABkK4UPbpvNn7dS65iw2nGS9rQc5Xou/8gr4Alnf87fWe/CcDgl/TKjOy+r3HlLf9j5iVvec/I/X+5v1A7xNj1IiXIGUJH9Yd56q8u1wEk/39KzAvU00hL+kd6nD2JqE75Z+QJGWSEBYAYZBIAeSzgOFMp5bPaRJtNtscVPmuTom4VO92gBGinkD0jnh/GOj8keQ+2fUV5z2Q7QTm/SQTQVeU43OLF2X2S9eFkgO4EyLEjeZ7NOp2yEC6CG2iPkH70PfogY+rLe+3Mwjf2V+MneyfwfPozJeZ4RgPmLcD1U9mH5ZyKCC8LhYbqaj+LWXlONUVM0E/HRVRobsksjg6Xq/K+yC8stHIKS9bS/hXDpUJmTjHgjsqzqpbJ54LFpXZgoa96RIV5PjH3MAeZdx7zFTL8t0q9UTMhwddzvLP3Phjr8MSi3zB+zMqDwrXx9UjwDF7T28eCd8vam7XHzUpjCk/Hxs9e0G558cAI64q0dy/redY5nGM8bCsM0pyw9WkB9H5umbCg7ZAX6wqICNYeQyIzXlQa6HzD0559+A6RHI89cue1W0QksNZiHYqhyonaAOsoxv71HMyneNixDmReXlmLqozt8kAnGtpcv7bbLOS1H0e2MtLyB8ebczsGj96by8WEvaJdvjpVb9ZyrMVYN1FniBPyZd1pXuPU+UbV50vTe8frjYUKOgHlYA3JGHIizwh+C6RCNTrNpSv8Vl3eLcdxEoxhk0roT8kc7g4nAScBJwEngY0hAUdYbIz37GrpJOAkcG4kYMAySgeKBWCxeRfYYj1RXJSwGkYBZhEOKcG9gLpYGBPWA2UHQgCgEIWKRTp5oDCgEAEUAd4BUGO9hLIAoABgZWAtefYrQCgQgBcoP1yLoiTf92bNi/05aQkCCnOAbtxngLlZoXEt91NeyBOU729RAuDg+TyXOqcJkzTZYAQE5QRMof4oPhYmCLmkD/Ms4FyavDBiwaz3AaFRaLB2JD/b04Jno1ymD+4xLw0jK8jb6sr9KGYoRjzHgPX0ngjkZ0QF38nPrN7IC/IjHQaLa6wuxN0HRDLvEu4zYIm2QXn5HZkAZBrZYnJMy5c8zYsCcoW2wDtFuez3jrC2ySd5o0gvyzEKD3tBbcnrJBghyTxNaCP8zTtf72FtnzaCUk+bRnYA/dQVAJfnouTSrmnDWPPizQIwwLukjfOdd8HfaK68U/MeQhHmHOVE1rwjnsV7A0TgfvoNFnlcu0zKLYcS4jfy5XnIGbAXoIL204y/+tEo/Me3e5mRHY3YD9tR2Klmh6I9mU3qp3HyfIC7S9q6z4gL1dOOBDsWCQExBEgOULcaqG7jgI0RTUC43oa+tLf/qgSoD+C91sG7eRMtRATRSGbU+7I2On+OWmFGATQgOwwMsvvpp7xLOyCzABhv773XZCz6jaP3Zn79fSvXhIrmlDsyXfMEbs7IE6AoIJ1+1NJTFELDq1VLhZw+8wI9Kc+MQM7ppXpQlwEooWO6W6oD8Q+9/OnWJykDbY+D+PW0Sx+QXWD7nlxr4TVhefjNikLz671rBsLK2FumXvZLb2lcdeuPX/G+7/Zk+/3uE8gk/RMeDYTuYfylTdM/6PMc1n/XmdVpXwaBlYRK6eUA8X6fyKBosFrUbqs59XM2avYyIhzYYHuHwOKrFZRnXERESWByR94r8sIosN9ARtsJePl87jK9i3KzHTzWbAVRsZgfy2ajZrVSsBBhp13YDXwj7cE8If9c31lb0Dchev+LUrrf9Ivph3ttmXUM4/dB9WO8d9YkxM53yCI24Fb5GP+1yXZ0hH1RqpXisNraJnlejHbaQSmbz2abjW5NJhyztK1u6Gk/mqjd9cPgO7/+1iyhr3Qw5zKfMgcxV2F1z7x8qxJzyGpjH6TdWsdf6gc8zBgfIYHos+wJhCU7czXlTq+TTpCV++ksSICxH+IXwmDFqy0Ofc/vNOVl0crmS3SB4w7eYWL8kctHx8Z3zWdHt9e0dI4NV2GNxRjJGo52Y3tDkNGCiIv61qtmC/vue9pCc76i/Vcy/M61dhjBwN/kZetL8zS4QueeVKi+MjI+sz7iOtoxhwJaeoXa1NCC382PaGPsoL1UzupsQSGvnjO8ZWD/4OZ6V/XgHiMGmPeR0U1Kf6X0D0o/pMT6kDGE+YDEBtuXKb8jBx64rCPvEXQDvEwgNVhf0Yf6jW+syIkeIO+KmW5jcUibbvcuXakRdTHPYddX+l60+9NJwEnASeBSloAjLC7lt+vq5iTgJHA+JJAGhlESUGoApPkEoGXcNSAWEBdAAfAWMABFGXAVoHWZSFgmPrgvDRzzDLP+s2tQTMwCkt/TKS0HwK7/rGRWY+TNs6QI6ZaoPu1lR1DaKC+kCsAYB+WmrHyiWJH/J5QAIA0cT88pAFamiJslGuWjnJ9SAqgGPCGMCsoYMgGwN0s2u4dn2zmTLXUmf56HpSLlBPRGabKypQkFU3BMaUtAjd4zrZzcixwoI+XC+4HnmGU+nxbOyYggnm/AOefI18gP+9vKb8QRzyAB4CJbwHLe+6QScfnNMpbfjMjhOaawmgyMuEBu5EFZLQa2tY80aZG+D6X3ASXAF5myNUe87lTbm/mohW6iTRiRhFxoM+s6el4W1MG8I/gOaUF+tHMAL2RvxBqkAXVBdsjSQnpRBsrJJ8q5kTqQEyZ/Qu9YaAYUWq4HOCZ/ngVpQd4oyijMAETIkk/eJc/DMpb76GdR9kVvyGQ+978y8e47O4rmXMiMe0tx1ZvKjCTvhesTsqLPC8FbBeTnskvtoD0CPvxfSm9XAvhMH7RfyALa7qRkhIVnR7KBtLAQaOTxP5UARK0/PpFHz2dJRAVv7kfDB70fFVHxieyuVcOtTOoq2s/nlWj7vNMPKmEVzvvnvST9TmSFEZ7W37vaVFs4uSJQhPGsQMvFoYHSQRESTysXclU1sOySgE3h6l2FNZoT4B4K62wIVF+Uy0V3dqGZJoLpf4wZjF/X5peOVHokjfwQhhOSN6xu+tDis/7d16Ze9iu/FZWGIISTo3n5zX/aHb82Ks486mWiExqOMr79d6WPKtFPeSZtljon4+zZttBmg3ARMBSbZ2KN/95eNRhHsrJODz94195InhXL/Vmy0z4BA3JG2aG9t2PtZ9HV/gEKSRI1lpqK1yMXFu0FUiTgFpt0i7io+GE4rvvHyuX8YCGfHRbwzDiRc3tZWItZ+/MEhAHtY0FtEo86QEbeD548vENCvtBXGFf7D/o33kEcH1BiDDVyjvHwgjrY60TtJDoyveRtGx9c7PhBttuVAYbmUe1NcUwx3grDxYJijuVr8u7xc7mcwkTFS8/Y+8HuFZMfyV1W+xpeE6wfGL8I78TYwlxzW09Op1LfN+higF48p+gvtGO8VpAh3+nszCUOfD0VqZ6Fa3teFrQT1qR4vRDeSy9Go5ViArKxAnsp9DyprQSsSQTsR9Njly8c23rVTKE02AnkRYYhEYeRUXghAOqzPmEOZH1CG7tJXhk7rn3R3s9+7RM3fCjs5pgP8YbgoL2wJjHDG8gMO1grmpELa98nz6HLV7LOYVxmvoZMMyMicXeZfNDNDSxND1ZFWHjy9NhfnxmItb/G0Pbrju1SdZnLjDChzJSX+ZU2y/gBgcdEQDtmpqasi8r3UHuplJuZ3LRLG31PhX4Ob0mey/hyMnIFGTcVs20m6LRvTIWCsnoz3kASsbZzh5OAk4CTgJPABpKAIyw20Mt2VXUScBI4ZxIwcBiggMU6wBLAKp+2JwHKCMqAhakBGEb54HfzfgDEBUBHmUJR4RoLN2VxY/nbFvE8z4Dstaz2yMc8JsifZ1FG5aOtZbvHnu7lRwCHeSYW5WmLZoAyex6WgT+qhLLCufRz04JOu9JznjpgvQj4xhz0W0psWPvdSoAmZhWG0pQmf/hu5IDlyTUW1gnghb+RMcqNWZXxfTWlLk0AoHwBalMH3hMyB2RHQeId2XuzkEYGsFMf8k57gvCdcpq3yRf0Hatrs8pH/uYxANFCnkaEIEvAErMmQ0Ek/xN5rfA8C98EQAJIj6KIMmsgLeW0MiJHygY4swzAd4/u8jJ+5GWLPJ/feQ/IgGT5k8e6jh5pwbU8x8gJ5MpBu+G98wzKxzXUl/Mo10akodgb4YJ88IyA5LF2gWy4l7/tXVNW2he/mYL9uL7ThskbIpDfeJ8ka1O0J3uPUfFn7owF7iWxz+NZLyz+tgvV0Xt3yBcQD9B8UgnAGqvU9EHf/jElwAzAuQMiLvwUaUFItLcpYWn8ut47oN29ktYgrwoPsiKxN1XLwV5VpBHg4WrHhEJGvV9vtJkZ0h41gfeQSKbPRNPe4ViGsYW3PgEGvuWOm73/diuPTI4M4Lo8AthvYUmpJpAmr30p8uVSvtFo+8PaiDsUcI6nQKdalhmqYscUctk5f8897Vx9MX7dba+HhEn61575x2e6Y1daHPvry0e/Rn+3TVyxqt6Za84d2XTvn75k5IEPfXXpum/PzD/vR25o7fxG1a/sPfamu7NDj3zU23r7273SjKLDJJEFVw7GIMZjSEP6N/JlTKI900bNw2oNEZ2V0/Sbv++V6Xv0+WalfxJY/HHtYSECKMqJDKqK3BnRXhVZIWTZQj4jGcb6KQpFUrRVx1F9DilkD6G55pSh2CO9aW0WIov4I9r0XN4smYJuqLe7wZS8YC44gPysSPYsZipCw++FaCP8zaQSY+O3KwHQrkZYpEvz7/UHnlXszfKzSozPtH8jcS8I4L23QXsIcUH51KcbClPmF9XY5EWVaS3MZar5OOx2Gv6SN+Y/6563ZZ595O9HC2GL+YJwdoDLrAeQCYQNgPN6D+YUSCDGAuZk5jJIW7zymL8YO5PwdOvN0F13ziTAHMTaCcOh65QGGYcjv+sRnqhYGfQyeVsyrpQpL8Kik8uHR7L56EF5JTA2s9ZgDcd6gjWprX9oU6w96DN8dvRtaeyyhcLgWHN68dgQc6URFqxHzGAp7XXBgy3kKXOArVv719hcR3+kTVMe66O0ycQTWuQCHqM3Bp2CPEgKMjKIG4VyUGotla8dGGtNicS4S4mwqLR/8z6mfdNH0BfQW1i3sa5jLbmo/BTdL/brswMVkRUYMtn6k7GFPsC6z/KijOlDvHawuzF/LBcFq0aOwmMS78lFEUwXxFjTXwH3t5OAk4CTgJPA2ZGAIyzOjlxdrk4CTgJOAmYFzmdiva2EYsFq3MBgFBdAJxb9BpRzPddwPfcZMQEQa2FHOGfKgBET3GcJ6a+1qAeIBxw2TwTKBOjrewufXfI2v3pEIYI2ybfdvCHIh+cxX1AGs9RCuSK8D4q47dtgz7S6pgFzfsM6E6X97wRqfyYpZByj1H+jEhZrHMjB5iZTxAy4p9xmYU9+KG2Uk3i7KE/kYb7k+3p1tPAN6bLxHGRs7v8WNspkabHvyQsvGMI4oa0acdAr6spHupz2DjhHXQjtZc9Oh4lCueW8hZ3CMg/5ch/f+c3kYMSNyd4ebG0FBRKLPuoP0IKVO3kh23S7MBKF8yixXS8KtFvA/shr7hPs+wiypZ5WH8qGzGkzp3T0SAueTTmQtXlYWIgr6ki7Mg8f8ufZ/G79AoWcPFCIec8o9bRVKz+gOMBtOmxWmvCgTZhHB3lBfJAf9UO2Rt5Y3RJZYU2pQ9aS6eZ7StW/1C9mXAL0JMb1PUpmVZquN+Egfrf3bvIiLRjnIhEXXYGmWLK+X71pUq1/q97CiFrjKzN6ixnlZKRFNm1XuopEFWl7LtytPKvePt0Thnu9UlzzbhWEP6E89+o5B3Qbz6WtRyItgke2vCKe3PT87P6fviG37Y6bc/df9tqwXtwcD3ZnMvPjzw694e2LmVzOT/rF8DWZ/MBQZ2zuUbwGwkY37t58z9uyxbnHPOVNewYQinf92Wtyj/3EPY9ExcHEMjfbXbolzhUOK8wTZPAtSrTZWQFgb8w1Z73Rr/ylN/D4p70Dr3u/197O0KJOcN2rk3TF+/6tN7j3DuWaYJp4i3yan5UmlejjtlHvWoT0KpI6K6fou+lwe7+sv/8ZeYgAitR3AnlRyKnCy4roKcdxUNH5OJfJtLK5zDYhZpuzWc0F2nRb+4jEQRDMFofKI9lsPKjed4WymNPpQ+KJlKWigRWdunIm3mIvRBvtiXGZeQMSF9KCQY+56kQH8+XrlTBkIKwb+dh8y7y+QuLpOecVVOx5W3iEbxu45z3hUG1vvpMfzOXnJvMDC3tKpe5CFHda0VDnGHMLIc1e05MBbRoPqBOFeFpNRoTbYo8fW9vRV5EP/SQh18+2B9SZaB8bNY+elwVj651KrIN+iHUAm2/77aYXCkTPPkFYMCixplH/yezW/g8znUZxt4iLgwObmt+g86xjWDOxzqANsG6BHGQ9RR8zg6FGrhBtu+Kmg1965NPXPCKvh6tFJLDXj5bgWdoPpADrFuaR9EE+q4UlS1/D4oV1EWs+Bs9+4xXa/V5VkbpqzZRRBKxsd/7A2HB1uN2qjjUHRVhAvLGesvU8cx7tmTGDepK/EZeTKvNX4yizU4SFBvUcpH36gMT5nBIkYH99uG7abzW/4DeXbntin+2V29kL6pNKyPyEboh9z3R/Ogk4CTgJOAlcAhJwGsAl8BJdFZwEnAQuWAmY0m7u/2aZb8ApwF8S+1UHyo0pQoDEIFZ2zkIH8LcRISuV7ttU+2TCMBAY8AFFis9lUK92d+DVH2l41euPetlRnmPWhRbaCkWMsqCooLjsUnqFksUyXw2kMJAdcISQFFgwXiZlkDwBSggj80Il/kYWgIDmeWLyMvLGQg3xt23MTGgj7sOajXOUDRIFGeLej4KIUmZkgcnULJPN2pG6GQnCOSzcrlRCSaLclNMIjjQpkSaJzBshAWeVqDPhaagncqcc5NEfOguQhPjARkzo65OOBLnrnU0rn5QbUB4lkBAAyA4y6YmYxU+A9KZ4AjiBlD7kRa2qFzZyXuNrRiyYFwt/G6mVxIE51aPXLhWfOUFfaS+UibobcUd5kFW/F4l5ViB73htAgr17i8lu5o7kbf2LIhqpx71cY3Kz++19JX0KYJWbVEZ9PW5z+lOt7ka7HrnSjv6j0odXqTzt691KhI2j/QDA7BFxgbdAHKuVRo95X4h9gYOx9+zokPeb6nE3ZjcrRFzB26LPEx6h/DTieW+T0i9FGkVlmH+P8ioor9t7UCn72UCQQlzyjqE/Hrhm9s7M5Yv3ySC2W9Rep9XnHP5bYSvlfdkoHM8c+chAmM2HmUx2OFKkonZx7MCxXa88XBwc8nd+/f0D2fb8UFaoivKh/UIKMkZMi4R4RvnY18ebTyO6nepVGn6Zash4QTgY6+s/uFIhdYfC4gFPRIc39Ypf9eafh6Pa8rH/tr/zttzxm7ObP/t7uzNBC7ICTw0sSy08nHlBnVhAZ/9X+i2eNox6GgFBAAAgAElEQVT/HFQ+q43Iu1vHB9qbRwcWZdU+L++IukJu1bI5L9SgJTIjDgoiKeQ54deD0JfheyBQuaL9BCqJEbyErw0FPEXzCURSNLQ5t6/QPsq61E/Wnv0aXqJP6JEJYS9MG22LeQpyDHCSxvhTJ6n6W/Q7ibntrUqvop0qv8f0yfxD+Cn6CWHKzhlxYR5PtEOlgsKxmasS/RSA1zwdIVeYV+jDXMM654n+uXbl8XYyK3iuov1D0tFHIWGZ41jTUfekn57L+p/knbmfTy4BBhq82DCCIO2EsAjlZRFpTwW8LURm18WfHtQwxfphUBtMDy8eHc5p34ZvHhxv7JsYO0BYKOY71k/mTcsadVIJAx/zFmXtXdG12W3XTE/kS8HXjzy8jXXglm6rcKg+M/hF5X11GOQ2qQet5WF48hp53t/qou9VSnsZ0z9YZ7OunVMZXiPPiKomxVlF7tufK4aKhBXRzvE2wQjGPDRYW1Ev1v30G+pCSvQV5UH5affIkH6AsQ8emOgHRjQg1ycRFlEQ/Eu7vnC5GCIRG08aMhhTyIM83eEk4CTgJOAksMEk4AiLDfbCXXWdBJwEzp4E1rDINottU54tfJIVxEJdGFhtgLpZgnNd+l6773SBACycJpVQOlACUJzIq+WFrcDLy6hr8XMlbxyMPTlQRrgOK2HbSwEFwvZvsLBBBjqvVi7OARq8RAkyAZCLv7HMBmQHjOJv8iQfFB8Lg4V8uIdzWJyh+AD682kbgOLCvwxSLJ+DaLAwTgCkADFprw2uJS/kau+DMpqixT38BlCOtSUKKPU3IF1fV8gk80bgfrNAQ2kDwADQAbjkO2VKEy5YuHFQDo7V5EYZ0sSDkVjp6/kdwAUlMF1O5Ic80vM8ZaUMyBJwZdxrP1r0OofmvKkPAeJQFgtFwHfOTSr171XQK/L6PvC26F2p+PXJ5sbU1bxJ+omYflLGFF2Tj3m5mPLKeeqa/t2+G7ib9owxwu84eTuyYn3vsu8q3iVhun5bibBuhItIH/R3CENAUTwy6EMJWKgQTlfkbmL/FAGJsbcrfpauka+PPCWwdD7hAVkRQUOoZWhD7qQHq1VN6Bvt/fuV8F6yAxD1fUoQGI9mo2Ci6s9nYy+L98V4lMk3C2Gbfgq4VM+GASFcFCejeXOxszAw+PU/LWfjgPEHsBNSERKBtvd2Jcadg1m/OT72xfdcb4RFvj71/MwqZqLHVUrhRnLtBW/bJ97qFeb3fWnqFW9LvDM4pm/9+fHaM187Onbvu+/edO+7CaGVEHIXAviZ2seCfgvI/YaebCn69dfuGv/aoalaODpUaQ5Vi/VONzgicmKvwj3tVEioMW12PiICIijk891sBpIwmxCYihdVDoKwXipon/OQ8T0ekpeFQkLFofa6SJPCx4nR/XH6Eui1J8JEmZcavenjSoTGYX2AN0UaoO9/GPM47QBQE/B/UglQkzUDoRCnlTfvjnECD4PTXbMkz1Ve/YcZNJhBBXMXdWDuojyQFCTmOiy8ib1P/4ZkgEz8AyX69qoxaJ70NIU90zmsznnuTqW/UMK7k/UIYw9zWuJx8lTrusqz3amzLwHap4WevFvfv2fFy6LVEJauWSOf1w49mfvz5YGyPgfUopuNuYFd8gzT3jvxJnkYTGa0L5LuZY0MSc6ajbZHf2JteocSfYp2yXoMoP/q8SvmqmOXLdbFnkdKQ+1GcXTh8MgHDz5w2Qs79eIrZU9xurU3zyHup0wWUpM18ctFVhzR8+PBzY1k03CRJ1PlofY2nR/XMzv6pC9TdvoQfZt1K/M8fQ4vaXQD6rmDfCSPA7rPwt9SbzNmon+wFnhSXC0KJg+WIYWCUj1XrSbECvPuggsHdbrNwN3nJOAk4CRw8UrAERYX77tzJXcScBK4SCTQIzLSS/FVl+W9UDTp+MYoPqA6Z6Smsm7GqgorQWLT2qbDgG8oIShTI97etx30rv1dwHUUcRR/fkexMvdvSAZzVQfMN8UrXScrsJEwlB8FhzwAE6kXnhYoOjzb9smwmLyUDUUHoANFCUCB75QRcB7FyTbHBojkPpQqC3nEcyaUAEpxXScPIzuMYDCrMerHfShZlBEZ4QlBmCrqwW/foWRhtNIEgln9pusLeMHfZt0NkcCeEgC12I3zG3OvueobmJ9+yel803I1Mss8bbjOPBfID5lZ6CrzKEnfb6QEcuR41GsdeKY3/WGAFkgMziMn5ItcqCvK9ddoOwrng8L7lI4UeUE+1tZPCGT1+sWpdIJ+MuIpldndvKYEaLuQfFhx0mbe0XclfYl0qxLWpYB89C3GDc4tamShTb5YYZ2MwFvzYdithrJlxjsjISqM/lu+wwJIkX/6ILTLjykBYKrzqWnoX0ZNTwOrvmb9OJN9Y+aJfSMYM2hr9IdJkRWMVwCy6QPyhXGFg3HH074VXnH2UXlOHFwqzuymzv0HxA5eYOlDZEfrJ8fv/sNqoX40e/g173x7nK8koWg6W66/4eir3vGumW9+y2vHvvTew5ff9ltPCexdpTxn4hRjIp4zjMEc3/X0ic0PaM8AcQ9Rq9HqLuFloRBQDX1fEBExmMt4ZeF+cbmYW9JG5nEYhBWRGk2REnWBVfOtjq8/w5m4FdeqFRGd2qG71giikSFzbjsTxXZ5pCUgcJ1xuClCgDEfwPZfe78ThoW9pd50AonRplkvAGJCHOPVSJ9mLiIfgFGOw8qfedrC9zFvpee+tAdN/1qCeSjtnWc9n0/WA4wdzIlcYwYY9HfGgpcrAT4DnjIPsxcHBKsdJwk8t3Ldx/QNTxQaIiTi55Ugdowwb/f2CMk4siIl3YvoK2D48158G22XtS/t6Xus+J1GTaC67w1u3lGNo+hbNS7NytPiGoHzs34n/3Xt/eAVq90J/U37oz8REso2cKeNQZAza/27Xp7Ml1yTGAJpKooUgimnJGbEC8rD7RdXR1qfHdle+8L9H33mnwTdPHMY7du8ZE9FshjemDEK9bI1sNa8Ge1fFi8WK11fXh6jzcVKoLBWNc2AZTh1eS5a6EzGedbsRs7Rr1mDIy/67n6/nf/ywpGRHfI2Ye28mifFqmSF1nfdTDb7bHmylDTc99frr3QCL03zpD2VertrnQScBJwEnAQuAQk4wuISeImuCk4CTgKXhgTOgZU3Yz6bpaJko0ShQOxXApxDiWl6jQfq3vy/3umNvWxA+1igdKDoo1QBDqCAoVEANmDNaFbyvADyNCCdvw2AsHBWABXkg5KDsgN4CUnAPQAdFirJQA3O45nAPQAS5nnBs8kDUNA8BQAtzArXNhmkrISaAoDEQ4ByG5jPteYhQr2w4CKkCXlikU1+lInnoFQS+gZwgvyod5owMCDdNC3bCJe8IHcAO6k7skp7aKSVNyN2DKixTyMoeAb5G8lh15vnALIzUCdNdnC9WZ9yj8Uj5vtdCpS808uWjnpzn4So4FlGEtEmkJmFw/pIT176OPfHKoTfuS+Ee+JaEqA/0k/pZ8Rw/7k1LqRPva6X0pfQrwxAWfVWbax9d3TY+6r2rPD1vRt3vJ9e3pVi3S+lz0o8zaPGBW3urNEqK9wm6XbPTDk7MUatdhhZsfJbvnbQqxz8ohcXB4bIK5bjgAIf2e+AU2ZpyjkAT8YU4t7vVcDv4sj9H8g1rrzlVQs3fv+f6P5bkxszuZuDwe0fnL7lra+978Bbp3obCq+70ufgQt79u5QICcQBUDV4ZHqpNlgtdkQyTA1WS9pD2xvQJtrtSlXhtlQreU4w9hYFVGlvC29R/bshTwqFjtN8EOsNZzNt7V/h+0HY1m94ZYUXYN3PgXjP+SPoAOZtwLwBMUe//pAS3giredpBVtjBPGR9g0138WSgjQB2MsfergRwamEfIQCYr5gfjYKkDLauMK9NC+nEWoD5nTmW6yHM2CsHIPUflCgLxgXvV2Id8TNKeFLclirjqX79Yd0AKMsYAuhMeB/zKqWcaQMTz5EVpyreC+562itth7Ub7XNTFGoZJUYhpz0swtD3iuVBjFAsrNGYvCqyAvqnjuze+vXSYCcc3VHbqs24aS8WipT1q4WohOCjzViYI1tTJ2Oi0rR6RFNUer400H2lvBbuHBxv7l08OnRIZAhz6KniNsyt1In1JvljDEQf7K1b42ahJNZ4uL2ULwZlhaHa2WkW/cpQ28/mYzwk0RO4XvNisi62Nk8d8DqE3Dms1fc9QSc/qnBWElcW4hPDqH29Z9On6aOrHgq71dbeFY3Ip5hPOnjORC+/9c/4az3MnXcScBJwEnASuOgkcKoT30VXQVdgJwEnAScBJ4FlCchCfl6W8ihPANIo3yhlKDSEMQAIQJkZ9dqPKRZ8IEuxHGQFFpNY0DJfWKgmAAcUFwBw7jUrLFMo0gBkv2U8ILptnowiZJ4Pdi95AkRwH2VC0UIBAvTgN+4HwCBZHczqjHOmnFmoISykKa+B/nxa+czaE4vvO5UgJ4hLjTUb1wGQ8GxiVAN8oPClvSn058q+E0Ye8GnlJcwLQM1VSraRtpWDe63c6bIdh6amnofilvbusPpRF8qVJozIz8gKzlvYK8pFnXlnkkvwmPfYL/A3yjX5IW9+WyavlkFV2so4bYcCu2PjSkBtwNP40X/QvrDKZkNNwq0AzPxy6iL+pn2udeB5sfYRe5/MlL13ak+LetTV2LXVeyQ+INI18P6zbqJfY0HNgacH/ZcxoP8AcGQsSx2iKYSQZ3rdGW+LJ47VnHlO7OCQ69S96sF7RVTkvNL0IxLUcdgKYy6gL/2JfvSPSmQIaMW4ltAvI195f3fhOT+AVS8gKRuWc0CS/qnSjygxbp73IxUWijrckyoQYPHgq2+5bvGjdz7i77pstJ7PZWeiKN5TyOfKErU2lPUqQSvKtrr+9ko57yuDSqutnS0kr5LiQWk/i2wll1mQm8VB3480x8T6Vb4Z7jjXEkDmtFWbC/6LvkPg0V9/Wulk+iNzCbHzOQixyHzyq0p4JmA1jZcncxSEJR2OvsH8DoDL9fRtIyoAPzGeAOx9sRJeTRgC0B+YVyFS2EuH9QnHm5VOtilx79InfeBVQpuGxOf5lJd1Ec+ZVGI8M+8QM5JYKy93/iKTQM/LwsbZFZIZ0sLvtrxI++t4JVz0VuaI5fWXQiHNHRgb6DaLjRtf9eBeeUcwJ9JXzIAE4J92y1zIuM86ywgIIy+Qls1T9IsbFWYqXxlu3bd4bKimZ3D9qR6QiPQp1nlmMENfZN1NW14olP3Z8lCnItJiWOTF1SJbphUKakqJtTPkIO2ecvN86kGizPRZ1udDmkmf0WmU7j62Zwt7bhCWEdnRb3kOz3vyEccH5GzXlGdFpbkwk42iJ/ER6Bg8H2/leRcO6lRfvbveScBJwEng0pDAyRacl0YtXS2cBJwEnAScBEwCWI2h7N+vhNUTwAEu4ygeKBkl79hfL3mbv3O7t/02LIHZ8A/FwazvDYxHgUcZMoAdgAPlLQ3op639eT4gBIoPCgwKG2VBOcRaDcUGBYdrsGJE2WOOMgtMwAgs1lCyuA4wwTwGDMinLChmHOYFgQLIebQh86owsJ/rqANAJ5ah1AEwgnMoZNzLd8K0AFogI4AQIyd6j1rx7khidfeeRzmR8729c2lZGGGS9rgw0sJ+SxMX6frwnd+4l3eB/FAkjaQw8sjKyDVWH8LSWJinlrf/HQVv6cvIEYXWNgzlvRiYRBshH96TO5wE1pIA/QarVNrQB5S+qPQrShB2JyIrVssv2exU6a+VHlPr26vWfq9acCTiohAdVD/uJG0e6oQxATADsgJCAOLt15SMxLD8ab99hIX9tExEpLdbh7w46R4UT5QckuYmTxtpV/d91mtd9ly5EHQiAVrUA7AFQgJi9X/2yomMkjj3StbnEuBz3w/DlSZ97Y+UGJt/ovcY4pB/4r4DtW/TJ2N1ckAcXAAH5aWOBqYRGuiQSIsY0uKKHSM1eUvsr5YLUS6X1QavXi30ogG916w21K53taG2zo1VysVj2mR7pljKhdp8+xF5VuyVJ8aRZsv3tZH3idmiC0AIl2gRLGwihB+EPnMFcwkhWthRYkKJeY6NdftDsaVFwvxqB+2avTHsgBRhjDAvQTtv3oT2t3lhriVqIyv4/XTICryd/p9eWRi3eD7rH+rO3M96gLmUtYNrj2u9hUvjvHmWMo/hNbYcj05vvduqax+LnFJxJlcodTVO0daY+75FnhadTqP4Z3670I6H288T4G8eev0hAlmDseYyDGa1EIJVeVT8vTwWBOZXSnr2pK6/UsnW2Kux6mtJP+3dx/rY1sjycstcplBOc0pZzaalbCHMiLSY0fjMmp/5lPmN/ssaGOKdMYF+wFqSUJCQiOKbM3ONuaqcBXPPL1b8ouRwR2/fDQvN1l+2hjYrWtJm5q3G3LHrgg5ZHnfw/HcqYfBD3emP7nAScBJwEnAS2IAScITFBnzprspOAk4CG1oCKACABCjhWFABwrOZrMyCE4AdAHDRW/j0qAgLFDXiUL9WCVDBrAvRLriPvwExDEBHsAbMp4Vs57jONqZG8UEpQRnCopL8SJAZlCPtOQDAR1gVfud5gCPmKZEO85QmS6xMdh1/m9eBlcc8HMiffFHk3qiEdRwygkghJAaKG9dQXhRU82agjkZ+WF7cC+GCQoqVJuFSUBhN0ewHO/r/ThMb9luavDAiBtnzfpLY/DoAP42s4G+Ld8w1yJT7eN98Iu/f9x77ZTYhRSaTSgBJeFNcpwTJQn3fo4SXCYDrJX/Ie8D2MUksaPEocMfxEjiBTCLJD1ARIGOfEv2VceMHlSA313MQJ/6DSgCF5hnUVav2M3lvKXO1/L7uXen3f65rACkt5Bx9k/72X5UYUwg/BcBD2/2MEv2acW6Nw7raamTFcV2UelE/yki/whobguT6XHNmVhtwT+faNd0Q05foR4SYoy/R5wC27DDr7NXAT+T4s717f6d3A4Tq7/XqkewlIwLjvJEWKS8L6vYWJcLwcABk36XE+BTvP7LY3rF5cFYhn6JSMbuYy3pzuVxOY2OsOmaiaqU4Wy5H8rYoFAI/PNzthFPZcmZfq+1PtbtBWx4awS/edrMDiFMN52x9VTijtQ7mNtvjgvmJdv/7SrZ/FR6Yv3Ga5bLQOv239+unZ2oTE/P4Yt4jjBRjA3M/8x8AM2GwbL8ByIoVJNWFezrNN3zx3UbbYOyGfGd9ebNSVqGLFBYq7+WLFREWBdZ3dthK4V6RFa/Zf9/OR66/dc9+eS6wdwrjdv/8xxosHW7Q1o5pSeGpMKETw7liOCfwn/BqeAKzhjuj2I3fLj5r7uDY4cpwJy5W/XYUZkLtOzSiFSRECh5+kP3MScxpX1Ciz9L3CfvGWpw5+JtGdy6+vN0oFbrNQmN2/6Zme6mEZzF1NU+tFYZd+4BMd5tLD9SnD90S+j6MR38rgUCk/z2u5DyZ+qXj/nYScBJwEthAEjijk94GkpurqpOAk4CTwMUqAfNQQMkAWCdOLaAa8wGAGiDfkjd35+e9KBiTZoZiAkAHaI+igoKC4gFwAYgAUAio3U9UGMhu4D6fKP8AXNxvhAUgI+A6yhCWmig3AHLkmQAlvd+x7jJCg7Ka9wXn0sC+Pc/Kk7ZIMy8G3bICfFIOy4/nUUc+J5XY7wP3d1zfCTthxAO/m6Wl5W9EAgSCWVCj+HIPcrLf7dl8pr9byCfKz/0Wa9jCUBmAa3G9LVQWJIt5oaTlYPkZ8cMnZBR1fdh74Ac+rU/27cCaFMWUd89vtAVkD+jIe0D+FtfcynzJfQpsRz60bd4XynlL5xYF0D9Jk77kKn+GKiRZJW20R1w8rO9/rPQ+JcaOb1bCcwcLfLynAHNoo/QR9kHASt/6LAAPYwVkIW2Q9xF3/2oFuOCd0D9IRkjy/minEK+0YSxD6bO2Fw3jFM/HE4D+iGcAYw4EI8+GdBCZGwNYQmxA3DEWQfAeTD0LMot43vQRAz8Jh3V7vjG9t7Cw/3BUKKs/ZQFbyJt6GOByQuvsFAmgW5K6/WGvrAYG/3v9jcz+Qy/f80paUMjeAZhmB+FAflXpkZ6XhXdkpt6Z2Dk6qxfVFfCmfSziRWF/M34UjIuQQJ5HRVYUFVZkruMHs9q0e06bbze7fth502ue6fpfSrjn+au1Y9o2YRIhDOl/9A+A1O9SSntTPJXimqfVU8kjfS/9mPGEeQ1rceY1QGm8tZj/IC5YlzC/0m8ZN5w3xZmS/sWVD22atRBrPzwItClRrC2/Ag9PALwsCpWBKJcvmjes1W6HRvqn+53CDu3j8E/5OHO/vCy+ph+ZW2hzRs4x/5CYGyDL+vMhv6p61q36PFIdbY3Ujg0/GnRz9D9rk7aWNSMd5lv6JZ7KrGOMEGHe49yahwiKI/KOuG9mctMo+wjJ26KhfTj2agNw5mHutfBwkBX0dfoLG9hTJ8q+V/cVtHH3+JaJ2YdmJse/qP0whjOZovLLML7jEW3r/qQcUehXG/PHnhP4nW3Itu9gTQA5j4wmlS759eeJ3o/7zUnAScBJYKNLwBEWG70FuPo7CTgJbDQJAAB2BC52BCwCYAMgohBgvYUVMKTBrNfafZ136F13eE/7KcBGLMxQrFCWUIogMQxIt3BMJkeuSYdoQqExgB/FBwXI/uY3lBnAd5RDQHMAeIBCnosyBnAHCWD5cg9zF8oeilmaODBvB8piVmtGFBiBYn9buAv+pk4oVAAwKEnka5ZjgJwoaChRRqJQLiMEeFbaA4LfUBYtf+pje0wYOcI96cMUV8uL+vFMkxN5kpCTAXg807xbrL58oiAaiWHl4h7qR/l5xx/3jn2AUAcAs7x7QPq9SoBN7FlCeWkbEDXk1WXvgkvV40B1M8IH+VJfkzGyXD3+8vHvz/2VkgDEhWRKH6ZfIU/aHAQBfZ1wMlhkY32JdwLEAm0PkNDCwNAfLGwcfSY5+izA0+Rc8r462PYvH7xPgBrb1Je/J5XuVLLxh/sZW3gWFqTmVUXIJbwoIFToD5SJvsO4AIhJffAiMQKWsY58+bsTFQeC2rO/N7PjH/6TeX48lY146ZtmyY4XA8dtShAkkEFJvc+np0WvTInHR+rg/RKDPe55R8S//r57u9fuGl9QmKeWH0SlrNAskRXajDuTkTVvU2GjvGIxlwnCsDlfa7bna21f97owIH2CvUD+pN3ZxtdmQf2bOgfBj8EDa4gXKEHsmUcl/Xktb4rVqpW2QD9RtTF46A8BxXjCeuJflfDEop9DklJWSEpAZMZ6xgf6u5XRQrTZHhUXiLhdMc6xBBjLmb8gsQDmV8KddZpLnkJBKYxdNpsbKHT0xcIrUcTLCYNUOza0pJBIMwqtJHuf6FGRFjfqN9Zb/YeRDatWT2GWalGQfUB7Y+REgPxYrxzMa6wPWftZKEbb44U2D5HImt72rWDesrXwWmLcoee8cP7wSDWXj7zLbji6XRwCaz/KRz+nP12hhEcFfduMBOg7ec18W6IgN6eTxULFH88VgoV8KdgxMN68028Vdsrj4mWSC+t5PCkW4jCc79Rrtcj3n7MKWcFl/1uJfsr6gffgPOzWenPuvJOAk4CTwAaQgCMsNsBLdlV0EnAScBIwCfTARAMBiUELaP1qJYA7LAxReFAUtnq735wRYYEFIgq8WUOjFJkShCIBqIRCxDVmLcZ5wADAQe7nHoA95hw+AeLMqwJggmcDDgIMohzxLAAOnmObcJrSCLgOSAGgb88HfDBPB6tb2mqt37OC56Foch8H38kfZZDv3IsrPwoZ9bP41QD+HObFYd95JmU3coa/AUH420IzmZJnpIopq+TFtdzPtZaHhXey68z63JQ3O09+XGtKqSnQlIH6AcQiQ+rGOUAcNv19Q68eWKPzjvBg4dmQUwTT/9veJsthz3J+ueaX9sH7RvlHTshiNcvHS1sCZ6h2KW8L+hqJNob3A2PEx5WwyOa8eSKYRTOyPy2r+hShYZbgjEl2tERo8Czrh+maAmhy2H0WQm2fztEnGQO4jz7a3w/tvgwhYzo/fldm0y/eddoAS5+XBXlTtncoQVSY9fr/0HfC2WDteiEcyOc9SoBqHOaJFhqZ0iMuuC744F17O9pUO+MHYS2bzURD5VI0t9jMLDW6mWIhF0FWXAiVOtNlEGlzoizT88Gq10mGZ7pIp5TfKiGjjFDnvR5Q/4LoI+7/PykBcNIP6PfMpbuUsMh+sRJW6xyMB8zj69lM+FO67qW9+/CCIk+e/5+U8IYijy8pQZhg+DCpxNwHIUo5+Js1CWMAh1mrM970y/60+28vb/dxEUtAmztHz3vxbcwdtE88clZCCWrPBa9dn5eHRbIUTJMVKzUO/NyISIZydaQ9ms2HrIHx9EsfrLnoC2uGORNZcaBVK08+8M/Xb28tll8gwD+9ZxvrX/NqZn7CQ5AxF4OblymxlrWysYaBeCG0E+MqiT5HHsy5Sbgq5T8WdPLe3MFRb2jL0tDQ1qVtUZhtagNu29sOspFn0rcwQMCgheNKecZt0nVbtd9GKLJmTJtvXz843mAD76qIm6tm948Vu01tw6FeFQdBp11fONhpLDEOrHZAJlJGnkdottNaC6yRtzvtJOAk4CTgJHARSuCE7P5FWB9XZCcBJwEnASeBU5CALKH/uy7HwhjFB8ssPnH9RpF5zLvyF+/zrvq179Z3FB+ABggGIwfMVdu8HszqEiWHfFA80kod54xkMCto8jDSA7AYZQ4LXUB8lD2UMMuH37CUxOrK4mdzrwHL5omABIwY4F7zcOA8zwe8Byy1zaY5Tx7pDYKTGOxKgJbUgXL0W3KmgQ2ejTJnIYXSVvuUxazH7R7qitwNDKUM9nzz3kiTEny3PLjW6mJkjMmW+lI3ymFhswBpUL5RAB/ybs9gEU6Mf5RmLOmer8QzCSvA57QA55+0h2yUz15YKHtvKMxNyYG25o4zIAG8dHTY2JG2EqW9mqfUmmDhpdLv554AACAASURBVOrhs5poAfpTB20Sgud+pfQYhOcZoXOS43xswt0rJ+Vjv5K/6RUFIgWQLiGCrFyrAPZpMtaqYaTRk8RyvgH7M9AFTpiF5MMYbuP5k4C6i6H+Ii1sLgZgtTmceQaQlPmbdQUhcpiLmFeZf75ZCU9GgFfIBwBXwqFxDRbdzMG0iwklgGRCWUJQsM4gT/oEc6N5Szyu75AVtrYwUuJMeD2d8B26Hy8NCYiwoB0zvrIn0pv7a1Ud2+JVhse9fHmgIyexfuKiO7Jt6a+f/W0PhqVq95i8LFh/fYcSITg5IMTTG2Gns6+JPPjfU49t3jO1d/OLBPa/ip18dI71G/us9Bua0u7xVMQjELIO4yDmCtbp5ulMf8HDIfFySB3pckA2YrTiKQSVt+O6YwsiHR4cv2J+UKGh0Avoy4zneOBSlozKNCTPjE1BN19uzlcGl2YG4jjO0meHFb5qIPSzBZEefm1q8PDC4bLIwsIr4yioaJvtSJ4qg536ghf6x0V7oo+zF9LtShjVsPZa8bAUkdRXfPenk4CTgJOAk8BGkIDzsNgIb9nV0UnAScBJYG0JYE3/E0ooM3hXoEhBFOBVsMN7/NdnRVigQGDha9bGgAZm4WUbyk7onHkUQFwAIpiyYeA/IAaHAemAM1yHAgR5QF4AEYANlIPrzfIahQmyAgXNSI/0Jtic6ycnyJ/7KAf5oDgaEMQ5lCvAUpQ8nsV38wKxzbyxFLWwQGZdzb3mAUF9DHjDQ4U8LOyMXWNACeXjOwnlEGCP65ElzwckNxmmyQkjYiwklJWDZ5u3R5oIQnaAN9QZuQLgAGwCDmFZ9wolrLV5x5QVJZQ6Il+IFNrERjxo39b+kT/vxh1nVgLW//i0cSF5wkYiJE4m0j5PC/o2YwUW5uwXYRu+/qC+/67S+Q6dRPnMcp2qXa4QT2O5bMY8V5LqrgK4Gzm1ISza1+FhYV5yppuZt9FFIx95YVj/boi8SHtQAeoy/00qEVIN63JICv5mjmauAjT9iBLzIDLg7z9SwlgAIgPvS2trrBlg9Sxkm3mBMjfaHGskaNL+TrCpePK7O5wETAI9LwvWUO9WYryFkF0hJhTSyFMsO68QBIdLA0NH9Z02SlhVjmJjofKt8pD4fGmgC3lAW14hlvWddcZqpAX947A8HaYPPbh9fGlqqKTvecJM6YA0WO0g7xcpEX4N8o6+BOFH3+AZrCtJ/N1PWLDWYQ3MWjAhKzhUbu/oo1tHhxeXdoi8aIm4MEMa1o+EKHyWyjQcdnODIiYWa9ND091G8brigD+g8E9j+WJ4eaHSjZvz1YcyGX9fdWQqM39oey0Ovf1Bt/XcdmNRe4G0kz1B+g70jDuUCHnIOnWFrFi96u6sk4CTgJOAk8BGkIAjLDbCW3Z1dBJwEnASWFsCKAhYfhEWCgKAA+ULRQaPipd5nyp80Hupj3aB0gMwMNG7jjmEhCUaQIIpYQAVXEdC6bOQS9yW9uwDLEd5w3IM60oSfwNkoiQCavA3wJft1wCgT354A0AQ8HwL1YRiZZ4VBvijBHIOQI18uZb8qB8gCeAIyhrlMkKFcqIs8SxIAu7hORbKijLZc7g2fVBmIxgoA9eaBwryIWQGCiWWpg/1fqM81PclqYzShIidRsarWSVzzsgHyk05IX74juUdyh/Pe9j7yrdTV8IG8K4BjlCokQ1/U07CatyRrtAG+k5bQQ6kDReKoM+q31572muJc2tawJ/Mwr+PkLhoQNjz1f775Bnp/bBx8C1KbB7M8dtKkJEfVjrfYZTYsyI5kgYSx5d/9M7dB9l4+3zJ7yJ9rhHQzDvmechYZOTFRVOtFHkRibwwQwPKD/nGvEiIJuZcwkZ9Xol5i7mIOZS5yMIYsu6ASDdPLAMy7dPG6jSRf9HIyRX0gpUA7XFS6bd6bY+xF28heQZ0vHZtnjBHVxbKlSNZduLJPLG0jcPslsZ8dUybV+NZBCHAGpkxmjxZu9LP0/taEC/usEJBNRVGaVhExSMKsbSeUGkmPAx/MDixdSxrb56DFy/rTvoK+aU9O+h3rPfob3g9JSFSVQavtVjxBsaaVW3GXRJpsU8hn8iH/oeeoOvi0dDPNdr18mw2G18+vH1pXJ4gxeZCpVIe7AQiORbyRT/yW/Gw9rPYVB4s755+XDsU+b4Xdjt6Rqh03BKL9SvrcfOOcmSFvVn36STgJOAksMEl4AiLDd4AXPWdBJwENrYEBCI2FaoFzYHYsShVAPgABWwUCEhQ8qJgwAvbX/ZyZay4EoVNB4oRyhdKDuA/1lsQBoAQKGkADwD9nLONd43Y6AfdUZhQ6nguShT5AqzjaYH3A3OVeTzwbPLD8wHCIz2PGdjDNRaagnMobyhEKGs8m3IZSUH5yANAxaxAAVMsPAfXG3mQzpNnpAkE/uawuhmpYcQGdeN6sx7F9f2DSr/QKxfXm+eG5W3PM0tRy7s/NBS/myLKbwBCXIsyChGCDO/3wmbBm/04cuAaPnnHKKHIAvd72kBEm7DKbKTPHqB+vq3Vz5vI0wC5wHHaj4Vvsn1V0nu0JOXUPQ6QPndvjH4OCPVGJTbd5mCD0lcq4Xlxzt9FyhOEcfsOpVt7DBckNOTs+SZSzt3bOcmTThLSiY3JbXxnHrB9osiV8wX9bqEFV0IbpR95IYeMWt7f5TgBUQfWCmlC1OZTCPz03Mr3BnmcRMQn+/2CaQuuIBe+BORlESo0FGshyNgPKLF+tfVvEs7Ib9e9KBq/RmyFGc1QsbqIjMHa1NA3bbt6Zq82op7VxtsYhhgJiUEQ68E9Shjd0K/b8lqo+e1CrA225xVmCVL6205BSuTBetjWjBjFYHAE2Uc/o3ysyW0POJ7LOp01IOP0p5QgZBIvkijMePOHRu5ROKh4ZEdtv0Jb3ZTJxqxdb1EvPKJNth+WJ8aVraXyDnlZKPRTJlR4qHh4cz2bKwX7wiCeD9qdbHspLgedYFNrcfo1nXr8tChQF4XYYUOLJw68Twhb9SEl1qzHeeadggzcpU4CTgJOAk4Cl6AEHGFxCb5UVyUnAScBJ4FTlABhGF6vRNxbLB5RfiAQbOPoG70Dv/tJb+LnAXMnlGxzakAHlDAstwDADdw3IoPfUIpQQPo9Hyhi2tuCEA8oS4QnIl/c27Hm4j6su9LmWID7tk8G+djzzMIyHWqE68gPQgVwnrJYPF+UN8qdDiFB3mZFbvmhBHLOPCb4buGxbB5NAyzmnUGZLY4wdUP5vUrp75XwPGHjUEgZnsO+HemQT5xLe3EYsMM5nmkkhpWXvMmT8yirlOG5SvuUlkNhHf1ziAy8OKg3yjdEBRso8s6RC6QFbcEdG1gCIiuMqDDijrZLu6Kd0AeMfMPqn/ORIy7OWYNB3oBnv9TrwzwYAuPTSlionq+DdjFpD9dm2gObRqq5j975iCegPQHYextvn6/ynffnpvb7sLIch9rRh3pho5CXbRjPWG1ee5A/nLf5dE1vp/Ne2VUKsEZIpv46pGXiCIgL8UVuoDL1SAvmQ9ZprBVTR+wF7abXXpwtZMe27ssVihAEKx6/2iy72FysjA0VwnkB/6zPWAszh7L2og9D8uJV7MurYfexR7d8SZteX7N4bLirPSEwZrHQf+uRuBEVdi3rRYx62PeIUE6EVMPTlvGEccS8t1grQqBAWkCS/LRlIPLkO6cfH39YZMVXtl07de/wlvqtWqn6IlaKfju/TR4gY/ostZfKnW6zuDAw2tzZqpeWpr+2/eHBTTMDUbh4ebcRXdWqZXZ06oGXy2dk+/QksuIret5fKBHujb04kIvzrljPG3fXOAk4CTgJbBAJOMJig7xoV00nAScBJ4G1JCDL8vvkZfEG/Y6lEwoVwDUWWIAjgJaT3qE/2urt+rmSAvdyDYoQB0oRXhjMJXy3zbABziAFABxQjvide/ieuJ33fuMTAA5ly65/gb6jPOG1AVBqlmv9CpkpXgbe80yUMJRCAFWszfg0rwoURizEOCgryiDX40pviqh5hVgYJyMMjIxIW5xzLk1WpOtiJIURHUbkUB8IhOf1ygKBcGWvDIBS/QCNkRaWD8+gzLbPhYE9nLP4xXxHETavFOpwTCZzde/hNyH7SSXeBUoh8sH6jnx4rznawrKI3LHRJIBXxexCM9dodXO5XFZbEGS02WdczmWz4wKg6bs59ZyqztO+GBvocxbmwoGL567BAOq8SolY38T5J8Tbi/T+sJJdIXZPFqLrDBeXsWolTrvCoyyODpVyc4tNxjUHQi0L27yW0qI34hlih/M2ptO/GOeNhGJcx4CAuYWx3UJEOXDvDDdkl52TQJ8EbH31Hp3H4GNlLwjCGrWX5scyuVw4MLZtIZPNbsaBQARFvTLcDhQ2qVSfq+7XJtz0WzxdORgTWQuy7vywCIAJgf77935x15C8FnbFYeb1OncqZIWNG2kDIKsCxjx44EFMsPbEQ481pxnyUDeMk1gvG4mxstZW+a9fmhn8pctuOIpBEWvllpwjDi4cHfnU0d1bX6S9K66Vd0WczcVLfivf9rJhIexGz4oCf0zeFdcuTWe9+qxYjrbICnlt9A7GNNYQdyoxzkFW4FnBXJY2TLLrPbfh9ooo3BcnAScBJ4ENJwFHWGy4V+4q7CTgJOAksKoE/lZnv18Jiydi66JMAZCgXF3vdWf2ewu33+ONfcvNvbsBVix0BYoOigceDCT2S8DanzkGxcyIC9sU25SS/nAQWLGhyOBtQDxe28PCQJw0AWCVQMnhOZANKIVpa1S7HmAebwLKC4FhYA/3cU86FBS/9QNLacLCnsunEQr23TSydB6cMw8OyoMiisUb4bUgUZAVFncQRZA//N6fb9pjxMghKxN1m1QyTxEjM5AH74R3M+VNfQDrNZTtCSWUU5RG7sF7BYKIfGkD7thAEhBIaiSct3vfTK5cyFfanaA6WC0aITis6NzVoigMrCvzuexIlPWiHmlBO00AaYHltLXYeVqcvcaTCr9E38cT7flKxFf/bqU/UPpeJQCpBMTGov8ckhbmfWYC6KiQ5g2WhMdLAfJPEtKFHM7oqbzRXmg1srAQgxaCENmYF0UyH2q/j3SINeTFe2Y+tTB1Rl6k91CyOccRhk/lRbl7nQROLAHWrngr3KH0felLo6DrdesLm/PF8r7S4Gglk/WaQ1vqnxNh8ZxiRWGjOnmMQCb6src15gPypvj8I3ddPdiulf+D9r645fhoSet+LauRFdzMOhoPCg7GGYx2+ITIsD3b8PqFTCEsE2FBWX8nB+RLvqhYT3Fmm1JXoa3YquOqfCF4dHR7bbO8QhaXZqvNbDbY1G0Pi6/pllpLwc6pPbmd+ULWa4mqDruQFYSZWqkLawa8KpAnRjvs5ZaEKhUx4caxdb9yd6GTgJOAk8DGkEC/xerGqLWrpZOAk4CTgJPAcRKQZT3WTgDXzAuoFhb+BQv8rV7U3ulNvuNGL2yhXACcALwAfGOpBbjJJ+A5igeACp4OKEqQASTu4RMAhri6gDAA9igoKE98B7gn9jneHc9SwqKLIx02wsB8lC6eZyEyIC54pm38nSYNzNuCMlo4pzQpYJ4cfFqIJRTUJJSJks2VaaXQ7rdr7LOf3LC/LdwTcmDzXGTAOQBGnmUbi5Ov3UPdjdSxc/xtABayhOD5E6Uv9/JEBlgAQkQsW+m2Dx/0vv565Pm03m+8U/LgHVv4qi/22gDPdMfGkQBtu1Iu5kdn5pqbF5Y6m+Rhsane8rd1/PCGbMa7SUDDMxqt4IpG07+q0fJzIjTKQRCRjICknydEWgqg3TgSPD81Zfwjtvq7eo+/QZ8fVeJzLfDqrJQUUkSJceRfUg+4ZufWYeYIzjOe8/2cluusVPbUM6XO1J1xGW9BSwCHfKfv2F5Mx/WfXggtI/sZry0xrqfnJwfynfp7cXc4CaxLAj0Qnb6HEQhGHXgbrBzyQpQHQctrzBzZ1a7PfyHstj4pz4v9Iiy+WhlpzY1dtoiRz4r3mb4zdrN/xX6RAEPyVGguHBm5WXtX3HSaZMWJ6mFkBdc8QwnvivQakjWgrd9ZM5p3cJIn5em2ip48P2aU2CeprL0sLt90+cIPbLp8biCbb84FneZAY36pXDsWa98Lf7A+s7izOd/xalPavHtBy896ptVtZbTJ9koxCXf1r0roHMiBUFW+IyvW1RzdRU4CTgJOAhtOAs7DYsO9cldhJwEnASeBNSVwl34B2Ab8xnrXwiwBruS8uX+5wWt8Zc4bfgHKGwA7AL8BMmQKIA5xAJGAFRXWUyhDy/cvn4ecSKyxlVCmLLQM4A33kidzk20infbC4BkG3AOEUQ68FXB3t9BP5qlAfrYfB4om5Af1ARwy0oL8OIwA4DzPJrQVZAJgrpUjTRgYQGRWsmlPEMszHarDCA9kgFLIZorIASALDwsjDfoJEe5bDsWznHgeZaWMkA6PKn1MCYs4C+NFuZEJefI+HvTmPob1HO+Td2b7dpAXefKuuZZ3744NIoGeZwXtj/62SWaTURTFW7p+UC2XsmO+H14RR/GoUIaSH+j/ODpQzGfrzXYcVcuFrdmK+kYmUws6UbtYyI30QkZZX7b+tEGkee6qmfKy4KH04buV2IeGsB67lLCQpd8z9p5rL4t9eiTjEuPxLw8OlN6vT8Zcxn/Guw21AXdvLxjGasgK5p+EMNcxov7GPMC8xBjP+wO0S+ZH3RfqPSfwXoq0OHeNzD3JScBJ4DgJAKZrA27Gstt7Y9x36PPNdlEsNN7vtrylo/tK3YHS7M5nhgubJxaHFBpqhzwSMCAhxClex0buj4kMeKC9VKrMHx4JojDL+s3CK35e3/GGnVRinGD8OFMHYxDexhAF7Llh4U9ZL+NpwThta1NN/BltLp6dDTr5fKdZ3CoChrXiohbAxVwhKJcHF5t+Kx4Mu8HWbqs+jrcJ+3pEQahFtpazyytl8+Tg+2eVMCqytTn1XjUM1JmqsMvHScBJwEnASeDiloAjLC7u9+dK7yTgJOAkcMYkIAv73drLgrBMeDqgREwqXa0EkIJCs+Tt+fmS95xPzihIL4oX6gjgpHkbAIZzX5pEwLoWUIbzKDvkw3UoReSb9ugA+AfwAnzjGvNu4NMAduprxAIKJF4GgHOQHebRwdwGGGskg3l2QFZw2DONSEB5wuOBkEzUhY0QURRNDua+b/mZS72FvEIB4xk80/a9ME8Jewb3oixSb56D0shm5RbGit8BrbjGwj7xG9cjFyNAkDeKL1Z+k0oonQCFEBKcR97IhefPeZ2Dd3u7f/ql+o7ni+3vQVkfU8Iam/Id5t3r0x0bQAKpMFC01Ujg6Y4wivIiJjbr8+p8PjsgoGJwttUZLhbyXrWS98VODIrQWNTv2wpBthuEeU8BumvdblgfG6ls19427G1B+8XjxxEWp9GOeiGTuDPtZbViPW9hk/pIC0Bv9v1hLLDjv+nLG5SSkEPnMDQUYwlkBceANkFhnDGvO8C4ZB7YCJtv98gKG9shK9g3qKQ+hGyYJ64UcdFS39NYHQ/okzmTeYT5t6H7fRde7TQ6kbvFSeAsSaC3ATcAO4QCa8kVwiJ5pBiIKAxf2Gm2rpveG7z3smfEe0e1ks3kFFJ1eS3Kfexfxrqv2VqsfHLP56/s1I4NXa35lvUm8zFjwy29KkAgnI2D9SVlSh88l8TakbVwsoeGQkDJe6QwHkWZimrQ0p4WH89mIy/oxjdmc/5j5aHuHnmU3BJF2XGIijDwvUgLiTWOn9V5vLiZlx5XYq2fNuw5G3V1eToJOAk4CTgJXOQScCGhLvIX6IrvJOAk4CRwhiXwAeWHJf5+JYBwADEs+SEadnvzd7S85kM5aWYoHSgbtlk0BAPKHGAbbucAVRAIbKjHtYBXFj/XgBwUFoB0SAfuA6xHUcL6i8OICr4byWAAHloRIDsAPRbF3Jfen8JAP7PqNRKDvPq9NriGekJcYAnHM7B6pTxp4sPupfxcSz7IijpAQlAfzpkSRplNe7OwVyilO3vXGIGCfLgXEoNnkoeFpuI7QBb3c1A28od84Fo23EXeKIKcMyu+QZm51byj73uBF9apA7LiHfIuqSvvlndM+Xnn7tgAEkiRFbSdijbXLssCdBsW38WCiIrYG683u5cvtdqXKyTU5Y1m97Klpe4uhYR6mh8GzwnC+BtrjfaW6bl6cane3d5sByOtTlCTCwbtlH7kwkKdQjvS+8hY0m2MUYwZtndQ4uXVIyqS6yzrXhgm26OCfvzG1GPZiwivq/O5xmecYtxiHuCTsqzsl3IKIrpYL7XNsQdFTGyJ4ngijOJr9f0F+n6z3JmuEXnxjUEU3ag+d5USBMaEKgu5wdzCu3eHk4CTwAUkAUgLFYf1KmvUP1utaHEYj0/tyb7xwX8pTHfqmaNyvqhr1UZ/NqD+CwoFdf/s/k1fbcxXQ3lXvEq/PVdpZTPvVfKFRIDMPJsHdWMOtz3hplVOhXQqLS0eHXwoX+oGCnW1zcvEO7VmGPA73uiez0Wv99udrd3mkjwrWiIrkuW27c1jZSX006eUWHviEWhegayNXTi7s/lGXd5OAk4CTgKXgASch8Ul8BJdFZwEnAScBM6UBGRpv09eFgDpgGYvVIIIgGwAlCcG7oB37ANN78pfQ7kB1MdaLAE/lQCkAKhQRMiDvRqw4udvAHd+5zxaDQkCA/DcYp3znd/J0zZxNQLANi39P+y9CYAe11mme2r5t97VWi3Jlmx5iUmcmGwkgcQhQJIJXCBAthn2bZjhAgMzw1zmZm4mTAYuS0IuyzBAEsKahTUJgTgksbOvJk7i3ZYt2dbearV6/bequu9TXV+71OpNUkvqdp+yj/6/6686deo9S9V53/N9n4kN5PdMJcgwAkoTXBArC9wfsdIb8p5nHOXmHHPthGBAOcxagskV12dlOGXnOH6HOKIMZjHB7ya4kJ+ZzXMc37kWx3A+q9Q4z0z5KSN4gROY4QbKzgNb9nPfVi59nZs4IihYXrmvXyXuiXIjFlFGCEtW8JIP+REXI3bto0fcI/8veDARJn/O49pWp5Srlzrngn7bMAjQTmh/PRIa6nLnJOsIt1VihNpQtlWxKQaSOBxWXIt6kmRpJ0u7maiKuF1pddJuLXDhrnp/3JTIcbynGkvHSI83293Rei2uRGFIHxklCLdfIb50e5IAYf7CGU9MrCi7w8styHTcHLGDFcZ8CwVwFt5/rmO/U+nbi6v+uj4Jxs2YcamsLMqEGvf09M1DPR87OTZtLu0Yu570BFXJuoJnwU4ZVeyVOHGN+tjVgfqaRvOOXMh01d8UzDbbHMSRXLJlEpqDB8Iwm1K/og2MKZ9TqltvrbRhhmV/o2sdAbmFooi8y0G+/1XxLmVjbl584j50mkH/o3fGr5NY0XfDi7rjjcFsJqpkJ6PY3aOg3NtlkaDFPd1+XEJJFOB9F1es8zeuY8GxWWzCu935buRjFrvmosnegcmTd0zGZywf8rhDEidO6c25mrQ6xx75QjA2dbKx/9rnt492mi6dHA026f6eP3aktanbVtZnBt+wcrJ4hucQi4B4NwYzW+h0vvfhz/MIeAQ8Ah6BDYaAFyw2WIX72/UIeAQ8AitA4D/qmLcqQXYRBBsynAkPk6YZN/5ZLbt6ZMQ1rtnhwghCnf0QKxDj71bC4oFV/0xY+I6lhcVg4PKQWRD3nGergI1EhUTHxROTKQh/SHlbWVxeMWyWD3xCypP4zjGU2SZg5GuuoyDtKYcFAOcaTK64N7NcMGsQiH2sFphM8p2tvELYAg5TNoQOLD1wh8J+vjPpI2E5weo4rmtltfgYJr7MrZwu7rVsAUJelIlzzB0UxCBYY6mBCIHbLnAzy5gbZFVxu7v7dSdcchrBiA2RwsqM1QsrBCGtqWu/bSwEzHUP/W9SJCrtSTErFAMhCNSGs4FWq9uQmBGrIcYuC9OuYmdOt7od6Repy5JI5/QrpsXDnShJKnEUyyoj2b6lT5xs5iSA0A6tT20sZFd4t4WlSy7CVuKw0emmgXAbCFwwpIFI3rVcS4mVuWE3Sen/5ue7rXPPcqPxwY/fP/3tt9zwgzoO0ZYNtyKsAH610vwVryss5Tkflvs3V7JAr1sU38TG1bLl2TlnvM5OyEUZ1VsYR1gtZVuVqqkLBrJuWstcNqFeNCnFQtqEGwqSIH/Gqf71fAj06ar6gbYxWcSzeNKLPOusfn1xPQKMqcRjgEfBvebPliGBv0+77kWPfy12Iwci1781/VsJFXdNjgTtbfvSTAG249ZUO006neNBFNsCm4VQtcU8jAcXIljY+3LZHWpZsGB/PU26PLs1CEVbkk5zpNtuaTwP2s2J5g0PfiYdOPjlOoscnkoAbY1hLsmf8mcNT1jzMn8AG1yXfkGJI5uyUPHxKnzf8Qh4BDwCHoFzQsALFucElz/YI+AR8Ag8+RHQivu2rCyYjEF2QT5hKUE8h9nJU/NQzXVPttyM1o42rg0lWtgKWkzlIdiZ9OCTG4EAcYAVXeZGCQCZtJj1g/3GhIlj+WSfrSqG7KcMFsPCJlkQYBA9/G4WHEyKuDb+gPmNlV2Q+kagca5ZVJjLKM7hO+KIiS7cAyIEwskNSpCA5GMuqixGhLk9KQf8NgsOEwfI18zsrczlSVv5fsAG0o99lAWxg3MpP1YUYAjG5v4KsYKyIFYgaFDuQDPlj7jHfusFbuxTBORmH/docTe4J6xRmPy+l7rmon7bMAhYuzdRrC4NQnR5NCiKNFLnE8EaQJhCWyjkpmsrEPdAGIdtubLR31nYSVyj3k3bcS3c2Wonx0W0jtWq0ZBW0h/cNtyrNipqxm+LIlC4dsotKUToK36B21atRpkw3yYyaFg4xyKE9OGaigMxVavEx/XHZKeb0PcZlxjjuvMtLb5dK/K1/0eU/ri4OBYXL1b6sNKlIL1tbLV7P3bkxATjDuUuC89P9tZB3wqTJEV5GlLqdVGA1ifLFe//jQAAIABJREFUinxc75MVk+rbxQpMGykujLS/sKEKqiVZNpIm7mglDnhu8PxkfPZ+3p/sLcbf33pEgHfPTygdUOL98HvLNwGPrxjUbmo0UIq+R789R/tOTYyExzQaD0XVYPfgFVmjErmXLnDzjPE8R80y2A6xd1Czxj1UjK28m9t77mJYMi6VRQ/GIltY87hE1Z5uu9lIFT280ui9R2LFlvbURNBpTlXTNLlGgbSvaXLHc+uHFtIq3D06gBhwlItPFi3xDuvFivXYwn2ZPQIeAY/AGkDACxZroBJ8ETwCHgGPwBpE4G9VJvzqEgCbwM6Q5Uw8Ehc1Kq51eIuLBxuOxb9ZreuiyCY/L9QxxHNg1RgkFau4IdWZTJmbJyZdWC1AqO9R4m+z4OB6/AYJzwbhzu9ld0lGvpm7DKw5zHoCSwtIMq5PTAjKwrUpC4SaBfM2oQCiH2FgrxKWJEzqsD5gZdjTlZgIkreJDOZeylxfUQaepUwwLai1uWxCODHLCCw17JlrrmCKW8w/rDx2r2ZxAtnH5M/u6YC+v0gJvMAOYQjMuLctii0SuYk7bnb7/x/KQ3wLW9nMtakL6pL8sHChjv22sRAwd2b0i0hE+Hgc8pE1RaiyaDKLY4Jsu5b29apxy5giyGREIX9PAX2yLjOKtFqN20qbRGT0KQL3TH9vtT490yGksBEql4IgX3c1V4gV9H/Eiq2KIbJJxPXVkicmJBBtF7F9rVwFVcJYY2bg2hIxJlVhg2HmToRhPC4SfDIMQ0SkZAH3UGCOhdtrlF5egPMhfTKeXmz/51yOMZpxyFyOzMjqw8n6g7ErF2I3QsDtYswFiz51rB3qP7sk9NE5emR1MSCBoqF9PbKmOan6lTjoQrmK71V826qOv0bHKrSFS1TP5qaQZ4DfPAIegbWFAOMaFmX3KhFQmnfMM9xDUdySAQLWxldincCWJukX1Pf1riiZOtPCmyyblnkVwoe+ZmMa93km3Kg/xvTJuMr7rL0r8xyf1nF3agwZ0jFX6IcZfWfsRZRQWTJZOgRck3fJhfieis7rKG95fUwfTLrtsdbE2AskUOxxYyMPJJ3W9TIBUenMK+qyj/T36TqPKPHufKcS79W8+9sinLVVe740HgGPgEfAI7AuEPCCxbqoJl9Ij4BHwCNwaRHQyvsZWVn8ta76SiWIbqwMnqrUdZNf67iZ/Y+7dGaPi4f7XBRrQhJZwGtIza/NTphyEYBZDhMmW+UP+c+zh/0Q77cpWZwJYlJArOWEnhKiAJMvi18BCOVZk8V2MAsLhAnIHfKjzAgPB5RuKfYzmbMVq+RLXhZLAzdJnM8xiAvcByvEcL1kFh52vAVQNDN7Jq2cw3W5N8qLuyUTGSy+BOVnMxdQ5Xux7ybMUE5WpzFR5frUxQuUnl/s49rgQxmJG8B93ylXXYG765WUHSsKXBVQfsoDHncrMenFyuLvqGMrkP/cUAg8IT6qnYsg75EYQduFvJiNbi+xQu5ssixxnSTIOpk8P2VhNNRsJxIwXP/UTLbDBekp+Y7YWgmDnVEUjW4eqgzIV39TrY3+GMqdTerjWJzVrnLLlka9UhNZNCji+mpZqOyNK+GMgjLLn3m2R1YVkQQL3EFN6e9h1c9mud06oBMflTjUUL1M9vVUk9HT013cQ80TASCICMD9QSXzi44f8Z9TyuNZXMSNe0NAZexju0mJAKvmnm9Zxusilu1SZg0OschDCXrypyY8iFUhOXALweljuX6qVuJhuYYaVd1q9XIWtdvdqgQKyVBpX6MWi7QMJnXOiPI4pX6UPzt9X7qUVeiv5RFYEQI2tmHNyzhrccxetdzZabfz02OHH3E9Q1u6lXpvFlXrwxoptQag02Tcl1BwPNY6gCxN4qTbmYgq1VYYRnUdICFbVhouixQJZ3enNX2MY9Nu+/Fa3yZ5c4oqvGGmSfIY44dEkKvkYa5fn7wDnrFxMT2H0ubE6AtmxkcHlZ/OQ6TIrjnzVfusoZs4aU9RIi4F1ths71fiPZrFEMwXNkTMouXq2f/uEfAIeAQ8AheGgBcsLgw/f7ZHwCPgEXjSIiBC+3MSLYgHAQEJkQ/BPUt+n/qk1vX/QOK6o/KyLpdQ3b7HXVyHDIdcf54SLoyYzGFEzqoxVvyb8MDKK0h2JjZYR/AbZDp/8xsuj7jeXiVmSiRWadn5NnsyIYRnGcQ+XCtkPcfx92eVsPiA3OcYBADKaC6cKJ+JENyn+YrnOFYl4waL49nIm3KST+6Ptzj3M/pkFRvlhahDCKGs5haHfZTTXFrxad+LrPMPymFCC5NeBB8LTk55wIa/yReMDyphwcG9MBE97WYeO+0OvEklO2KCC0HSZ+OOzCYISywr7qVuyxf33zcUAvQH2iTtaLNWdJ8WWXpMthQTIss78lVD/Iqebjer1CrRiFrzaZEaA2qgcagvOlYObZyW+Ythr8e1aiXcImLkRByHPbgxUp70o41CTp9zwxnorVY1ZFZlLdEnvAbATS6BrhShLfdB7opUhLZW346Ic5JlS6hV92lFnX6flCIZv4STWonfqdWi6a3DvdMnRqdsDCuXA0ES11BfLHb+oD6vEPH9KpHeiKsXa2Nc/EulXy4u8C36fJuSWVikWIUstEl0uVhluhz5Zm2Fopf2Bx7jEiSmpERskjVNs1INT6veh1odCYByrzYz0+kSu0SdRW7Vwil1L8b9msQrBbd3m+I44Hlifepy3Iu/pkfAI1AgoBgMC2GRWz0oIDeDG+/KvNvy7vmW5YBL2k3XHD8lQaI7XKlpuGDQmJ7sYVVA0mk/szGwmeA2BJVoJ+2WS7UyQC6bGmGl2lUgjFPTYyNXt6fHr5VgcVQH7ZLocCiMK+/T8/tQ2m09SyLI9sbAcBBXG6243tOj53T+XiqNIjf9kEVFjwQP15w4JZFCr63aJ7HE4tItVnzGI+71diXej7lnrCt4p+Q3b1WxXMX73z0CHgGPgEdgxQh4wWLFUPkDPQIeAY/AhkTgy7priHsIb1bsP0Op7mrbZ1zcW3XJRMd10qa8ccsVU53JEOQUwacRKjANx62UTWIgSskHEgZynuMgTpngQbx/RYnJD3lohVd+HPlAuvPdbNOtIrge50PyIFSYSxKIWMh9xAI+IVARMRBCTDxgFayJHDwLEUo4HpIJsYK8zN8vAoRNwrg2pD/nsLoMt0y4ZCJvttx/uRJl5ZOysXF9I3E5pnwv9t3cWiFO4LqJ8nE+foF/SAkcLFD53uJ3xA1Wtd2hYOjf6478CRNJE2jsfO4LbLlH8KVO/bYxEaCt0Qbof/StvYgMWumdhlk600qyjuIpTIjYgLkYFMk63dGqy06SDofdQJ6hwm69FqsvKOJFmvWqIUenJmZGTk40Tw/310/19lTHqpUGfc75FeELN7CaVCBZVoRSIypyD1SpVMKKvG4odkWySUJGT5RlDaijUBYuEodcTxzIhVA0JPLaKSzCUXFZB/t6awREr0rQMLd44O0kSnBR6hiXHD+j9DtFKb5Nn9+t3//0ItYL4xsrb21j3AnlFirRNTdSHIZM7r66EikQhw7K38v9+j6uJ8POMAh3iEzsTDc7KbFLMKmQa7W4XokaqmvZY8ioKc2q3TQZlIkG7hD7JFJRqTwzvAi4Mcdsf9frAAGJGTMSLb6kovL+yTvc65W+Scnc8511FxIHXLs55RAN0BJkRaEQZDJ01LiPg0aJE07iBEIC78paGxRjgqG4U8nTFG/iZNrpSDDQoxp3pMpL517nWjP/yS6kINp5frLMcPXBzU7ChQ5LJIrgiYqjpH7PyJgvSWZzmfVfdZYlRpEfzxqsKJgH8G6LFR/vmDzveUflu3f/tA7aqi+iR8Aj4BFYTwh4wWI91ZYvq0fAI+ARuMQIaCX+3bKygJD/cSXIeVb73+FOf2azG/qm0FW2SbTo9rtKUHXt05GL+09odoSrIiZsHA/5D4FuogOTG8zFzaKA4yDTsQZApEAw4Jg7lMwVE+dD2CA2mPWCuU4yIofrQNRB8nA8kyquyXfcTCE+MOlDMEEYYD/7uB55IZrk7lqUsJbgOoW34bw8CAdm7YHFCJMz3DERt2I22PUTliAmWmhXnr+JJPzNb7nLHP4oNvtuFh77inJyfVa74QaKPCgzGzEoKNOsFYu4Znfgja9wD/8yZCH3weQRN1RsiBl8B1/u+23Uaena/usGQkAr2VnlTvujLUGEagF4tl2EhYjyUEJcsEehtrviTrpq7JUkSRqdbiprADmAqrhmNVCo0MzVJWCcFNlSm261o6SbpdV6HPfUK+mmgQZtGXHO+s4GQndltyrBIRQJ3T/T6u4OA/kez4KhJE16hXei6MunhatW0SZDqgPFO8hmJBKNiUcKiG2hIWa6Wqv0iufeIrzHhgYa3bffel/7x172lPmCAHX8h0qMWb9blIwVv5BMiJwXY+NaWH3ZZoJwLqQgqGyETfeZ6n67ilExpXoaT5NsUiLFjGqiOtXs9CZSI9TnoljLqCuVqCPViert6XS6HVlbKH5Fbs0kHzFBXU+LcpDcjQCfv0ePwHpGgPc9xlfeMxn/7lIiVtizlIivhttTezebvc9ZqwaXsUagxTChjaevtrbEBtfUSJL/NfuKOasz5P+a9e+ieBF/IrfMkAAyM3ZCggieCHllnLWwkPiBJcesxcXiG1bEvHP+htIjRfk5gQVJZi2cv7tKtPGi6lJI+t88Ah4Bj4BH4JwR8ILFOUPmT/AIeAQ8AhsLARHcH5FoQfwKSE4I8avd1D0Trn286XpvqLIS27WOnHTx0DaXxD0Kwt2ruBYQl6wwtRVYiAdM5sgDawpEAawW+CQ2Az6ALQ4GEzHYLYh7c0dlQkU5/oN95xMCn/zZME23eBKILQgoTBbt+ha/gsmVEUKWlwkT5GMCBmU2aw6EAyajlAdrEwQci2XB8ZC1XIfnq51DXmZhYcJLecWsTfLM0oLYG7h1YT8+4XGxZUGzKS8iCS4Helz3VNtNPVB1j/0WYgyCBW5Y/okL5r/P3jdlxirks9Rl8Zv/2LgImFsy2jHtdydBP0WFYDHRaUukUK/r1QpwReNO+0WUR+I7mmJUWqI6mq1OimsJgnJPK/hzq7dRafX3VEaTzCWtduJq1civsly8bWWyWoklAvXLzEIrZXNRtSIBI2m3g/5uN63LwgXLitw9UFgJNZ66WkcxRHRcb0UuofTZlbCRaJV+RbEs2lds7U9EkGcQ5SUrC0rAOPRnSoyv/1qJMeINOva/6biLFc8CEdU2xnGL97PRepvMJTLZToR9lUrQE0XBZvWxnmrs2h0F2taDodXpJGNyDSW/9NjRSLYKQgkWYSA5g4Dr0zrHnguM/Twr/eYR8AisfQTot7xzsjBEga/zd8y/V/oGpfcUn9+hT9yQsn1VaWsROPvsu0PMyPeenxaQCxQyzUOc6LYwjpy9BCKJWVnMu6j8vebvq7zrY6FHUHHeORmDOJu/59z86TvPmWwRd1ln34/f4xHwCHgEPAIegXNAwAsW5wCWP9Qj4BHwCGxUBER0/38SLRAgEBEI5HyFG/to3fU8ZcDVtgWK1Fdx6aRsz6tyFQO5rslQVLG4CUa2myWBuTXCjRKkOqIEZJoR/IgcTPKYHCEgQNJxnFk4mLhg/ttNKDAhAhdWWGewcQznMqnCwoCNfMxCw6rU8rYVY+XfbfWyEbG2gpz7wu2JiQ/mBgqSriyslK0pLBZH+V44lnuERET8YGJI+YmNcbMSeHEtcDqlhJix0yXyJXD6s5E78OuHXWeCCbK5vHq6vjPBZKUfK+KwYtmvOnyn3az/3LgIFFYWCHyIehAqtLcB8RpXZ4GbiFIFqg+Ju50Fsp6YiqRO4EdCvvePNtvdhgJEu1olnhDfcUCk+0in406LPJ+QsNGdabbbV10xhAug82NXnuTVct2ezYGIavnWUjwQsdTtdiJjlaxHK14ZoxRQNe1ziX4QoS3Nd0Yr8xExavLo0YlROuKwodqotXRSt9OptDpho69RZZxdyDUUaFLHb1BCsGD7P5VaEi1erzq6GCQ4Vme2sap4o84zFIok4Dk2qvo+LKuJa+TSq6qIuDOyuqgpDUmbiOvVeDSOgqYWPKt6g1P63pnuZG31vW6lIqFQT9acOvQuoZ7kI4O/vScZAjz/eNcj2UKZL+g774b/qIQQQNBqWzTz2uL+WXBi7kVXF5Jc+DCRIn+X59nA+6tZ4mGVbO+ilIv35Q8pYRHNxjsDzxmSd1G3urXjc/MIeAQ8Ah6BRRDYqBMJ3yA8Ah4Bj4BH4NwRYPLyq0q4RBpxI7c+4CrbO27b9/W6yrCEhf6Om94vp+tXyda8MeGizbhpYrJztRITNYtPASlvQgJkPmQ7EyfiUJjLJlsFDumDFQYTJAg2EyX428QF7sSsE2xCZeQ+ZD/kvwWxhv4pWzswMTNLCvLgGubDlwkax1oQQpuk8ezEAoTJKGXjWtyfkbQmULDfxI1yeW0ya6IIf1tgVTBg1TtuoPgdPLgen/xmgbcfdzMPttzRP5dw9HEsPZhsInCYWymIQybKYA/ev6fkN4+AIUCbo33Q5hG25D0/Oy5tYlyuiCYVZUE8eTotUjWpRNGUiI498ssvCUOSRpq1ut2kLaL8cCdLR7VU/LQLFNciC2YeODjS/a7nqv/7bUEErt+7JTt0bLwld1By+pHJ40faSuSwo5vkAqNWtAb1VjcP2JxUKnEnkeGFhIspEd5NKRuBYl40my13qq+nomjn1XSov96QeMQYYwLp/OtSF4wNrOj9h+LH/6hPgmP/y0WoprJrKsadjRS7ogxnInFJ8V/Slup5VLVzUBrTJlksSchQpwuCbRIoKoHEKgkaPYpFEujvPn6KIndULtgUVUZupBTIQpn6/nQRGqrP0iOw2ggsYmWQv1cqvgXPW3sPNLepvD9iBfynxbMYMcPehYk7xG+fUGJBzy1KuGZ6SfHJ/pcWefLex0IdNlys3qRk76Hv1nfeKZ9bnGfvyuwjrhmWuXzn/dLeyw/qOwtdcos+pfkWFH5MKsD2Hx4Bj4BHwCNwcRFYbIJzca/qc/cIeAQ8Ah6BdYmArCyY9EB4YWUx7fqffqPb9e963fBL5PV+sqZogXJlEtZcbWvogqoEjc2IBRBqJlJA7DNJY4KEyxB+s2B9TLCYHEHQM3HCJN3IOCNubMIHfvOfYUyizNUJLpP2KjH5M3dUll8Ze7N4YB/XRBAwN1Fm9k65mLyxH+GA61gcCrMC4Tqza2GfEED4bpYU5Zgbdg8WnJvjyNfcB0BegheflAHRh/xxt4IQ8YBrHrjW3f9zoprfb663CNKNqT7iBfjiVopV25T7zbKuYHWf3zwCZyCgeBa0H1ZSknZLsBgSceqiKLpRAsbTtEq8FmRZR6T5ddVKPCN3NeNaHa4oDG68Vq08pGMe73TSeypx8IgI2cmf+a6b8oDbflscgX/40uO9U9PtK9Wxb+6m2TfIV8dws51slnstmaq5XrkFquCvo6q42sJb/7vH9W8WV6K64nUf09fHexvV+wYHGvf31uPTCtp8UIQ3K2YXtWyRRQXjyX9X+qWiZIwru2Rlgcu5VdmKgN8QaweUGLvYWC2cr9DdKDEsDEzhwfNgs/rF1RIltqpKny6harsEjIbqa1hPhkh9Sa6ggk0SBqelWaQSBUNZMt2nxdD3y/3XgTiODug33PlNb7DA5avSJn0mHoG1hIBEi3JxzDLY3nd5N+Ydk3dmxk3ceWIFgXhAbKAblD6vxCIUxhbe73gvZGxnjCAfy5NzseBg/xeVWBCDoEH8DGK6YaXLM4PFCiR+513VxAw+c6FCKd+8yydDwn96BDwCHgGPwKVEwFtYXEq0/bU8Ah4Bj8A6RwDiW6LFO3UbL1MacJP3bned0Zobv7Pieq6JFc1PPtcVKbD56JRr7NnluvDw0X4XV3fqS+6HnR1KWAPwiWDAhIuJGZMkToDsIjFhggC1CR2TOYsOaAJG2aqB71g+4AaJiZpNABEqLKaExcKwmjDRgE9L5tqJYzie1XBYaEC8MWFEtOFYmywycSyvhDWrDbOwMIHCXFFZ/nYvTBaZlJo1CfdOQGTyN1cvrIK7W26gtrvpe/rc5FdTiRUcA64myjBBJU/2Mynl81YvVlhV+89FEKDP0c9aWs+9Xa6hertZcjwK3UOiU69NFWRbDqHGRaxOiz8/QnTQMAtOS6gYaXeTE91ud7LdDtutTnfOLZFHenEEKpWwW6vFE8L6lNxotdutRJ6BsvEgi53wHZBgNNDpZNVmq1snQLcGmiH5C2rWK7H+CLNKxU3L+uJ4NQqbGlCaCEgiwLngoqvxRXa3RaCzitcEC074Qe17K7+tYn0xluGT/RuLPPfq01yKrOJl1kVWjMU8146oXnGhFhD7Nk0lArpgopOmWxTnIqiEwYSsKQJiwKSxa0qkOCQLpjGn/qb6pW/mdau6Oqt+N5oItC5q3RfSI7AIAvNIf1v4Ys9NxuEpiRosumFxii3IYaxmgQ/vgFhBEO+Nd2Hen3nHZZwxSwh7h2XRCguC2M+YzLF3FMezj+d9nr/KtFGt4Hw79Qh4BDwCHoF1gIAXLNZBJfkiegQ8Ah6BtYSACPB/kmiByPDNLusccmOfGXVDL6q7mcf2uOrWiqvI+KI7Ilrt4bZrXC8XMq1BF2wfViBuC4TNxOx+JQh2JlMQ/ggZmKcfUGI1GfuJxcCEbG5ype8mBpRdOVmQa7OQgOS5RokJmwklHG/WE+WVZGVomTiaJYitFGdSxwSSa1A2Jo4ch6iAiMHGJNIChptFCJNA8/VbdmtlIoVd16xCsAJBWKHsXIuJp7mH4pj7XHei6pr7e9zoRzP30C+aoAGOuN4itgUBtXElxWSV32+jrso36L97BMoIEM9Cf6eytMhXVMr1UFsrvYcIyJkkQaLYCfozSMW09ug3Bdp2R7Uv1ULwMRGsp9MkOSoh47jEihnl5d1ErKB5JYr1IYGh02p3pyRYHBVpvU0r8OMwDo8GWcT40xdG2bh+7ygAdz2O4kTUUqfdJc5F0umrV6ZkARN0s7SjEaYpj1CcY7FvlirBg/rxR5T+uDhIJlrub0WE71/FmCOM1wT5to3xF6Jso270J8WpiAhSv0V96TFikMixWigLiliCX1WxcNuB1CpZXkjXSI9GUdwKI1kqumwCT1ECrhwDaaPi6O/bI7AhEJCAMP8dkfsui8q8Wy4Zf0iiB7/zTjgncirfTPtNpPDP6g3RmvxNegQ8Ah6B9Y+AFyzWfx36O/AIeAQ8ApccARHh75NoAXn/anfyg091W15+lavtGnRps+PGbktd45q6C+OqxIppWVsMuKhHkydx8lEFl0ZYBEBkYQUB2Y4FA2IGpum4NIKggYAzk3QIf/62IN6IG5jN8zu/2Uo0vvPbXiXibCA6QKCZFQfHcS32mTBRditlLp3Akwki5zPxMzcnrEzDpN6sQbgXrkMeXINrWwwN8wVMXogZbGX3UPzN/VjMDq7Hd8rFxrVMzLhL7raOu9YjN7qj76q4g7/O6rvvVkKYwMyf8iDOvFKJMt+t9F7V0WeKvPyHR2BJBIpA3ByjeM4pK+KJX3FaAoXaWtbptJNeIgCrpSNqRFoRTlyFaSVZCaQIa35bIQITU61M7rVyMbIaBw9ruLvCEb8gCOROL5NomfZJhOjIp16tUg0zWVUQNyRIXdaqRHFFsRF0rBzuVaKOTDMSnWdjVVa4ZTqjJLYKH5dC+v3v9eNblBBHGYN/TQk/JbaSf4V3sehhjJdvVvpPxREIx2ZJd6F5r8fzc8GhVo0m5erpflkrnVbd7ZZw0aPBvaKHRCcL0+k4jhty9YUOdVS9bFyC1ikdY0Fu+cxWUVRajzj6MnsEPAIrRABxojj0DGGitH+FOfnDPAIeAY+AR8AjcHkR8DEsLi/+/uoeAY+AR2BdIyDR4l/pBvYofa+7/revklDR44JKzUW1zHVGElfbGbug0RXRmbp4x7ir74CQx5wdF0j7lPChjnsoI+gh2yH/b4akUYJYw1qA71hecDyWGJyLEIAwgAiBWMAzjWPZD8kDkcd+NoQE9kPMmUsmBA72iTTMLTIsiDakm4kbnEvZ8PlLnlhVIBSY1QTlQYDB5zBxPVgIYL6EzdS/LITY6jkLpI3ow3cEB+7R8qPslAs/w8fcyQ/F7thfbnZH/gwyGRwoA+UFSyxATOT5G30/6C0rqDa/nS8CsrjIg9OLFK/JAqAm4aIiwrUi7lw8atDW6vC2LAU6nW5Cf+oWlhrne7kNd977vvBoZXyiuUnyw9VaVX+TRJ99URgqwHk4KMFosyxa+pvNTlXqEPEO6NtNxa+YqtYqB+We6+7+3voD/X21Q9o3FkUh4xPjBePBWStny26DJFiQF2Nr2erh+3QM48YFbYVYwrj5bCWLmfNn+v4TSq2N5r6ocOFEP2J8z60AJfAhMF+vPoTg3q8+1VQg7oPqVL3yDtWngPeHVd8ciwjNc4hnG8+ArhcsLqh5+pM9Ah4Bj4BHwCPgEfAIeATWGQLezHidVZgvrkfAI+ARWGMIENwakupT7oGfvcN1jh926cyMSybGJFZIpmjWXZCGrnkoct0TDdcet4DbuFSCmPmkksWVQGwgPgSEFwGov1YibRAKIEchb4yk53yujShBHnxHgDALCj4tDgbnsKqZPCD9uS5k0J1KCA0cayuBuRbCiokdlJlAh1iDsN1VysvEDX4z1yxmhk+eJNvMvzDXMesJYm7wnbJRVlxDIVqQ8FV8xB1+54S750cnJVZwb5QFgQiR4lDxyXHg8iklrk2d+M0jcN4ISICgP3XanWSm200nRKziXuKECNcRviu+woTECvqPFyvOA+Xveu5VncmZzujkVOsRddgv1RXAXNmMzLQ6h5qtzqNSgkZkUTEurI/01OLH+xrV6VolPiWLjHvrtapEimBcVhhtiRX0d8YdE0mXLI1IbwSoiBmhAAAgAElEQVRTxrz/UTrwr0WuI7qu1obVmW025q1W3usmn0JgyPtRMS4rBkkwpnSvrCxwDfWorGUelbuooxKoJqlTVSfH83yw5xbCuHffsm5q3RfUI+AR8Ah4BDwCHgGPgEdgtRDwgsVqIenz8Qh4BDwCGxABreSHOH+XEkTYtLvnJz7jWocm3PSjItCzCRdtasmjTN1VtyUu7chb9yGJFsf2ubQLkQ/Z/2IlXCthNUFQwduUPlgQNtv1SQBXhANWEXMNXDIhbLAPIoh9uJIyF4fkC8HDJ+Q/QgXJ3EMdL75jvfDe4lyehSYy8L1MECEQICZwPcrzdUoElGWFLH9fpwTZZ0EQ9XXORVUeF4AdxT4TVdjHb1hVgAF5c03uC6EiD9QqjOru8B/e7B74D9e79hGOw8qDa4ITIgX5QWiRKCN5vquok+KyF/4h3+u5NSafSmGR+G6JfeW/7bjy8XYM+ZyRLryEPoeLhABtkjaGMGjtjHbI3/mKfm9Zcf7IDw820i2bek4ryPJRGVF8ZVN//UBvo3KqUqkcrdcrXx3qqz++eahndNNQz4P1WnyvYlw8VI3jw7298aN9PbUxSRXUBX3e4uWsiNguRIv/qfMY/2y7GYsArCQsneudFRYUlAFXf7YhppRF23PNdl0fX4gWYGLPGOqMZ+YjSljXjUjASCVUtPWpQOwBzwbEQY5BhKbfLeTTfl3j4gvvEfAIeAQ8Ah4Bj4BHwCPgEVgOAe8SajmE/O8eAY+AR+BJiACks92WSJILJkTkGgpi/78qVVw8dKPb9WNdN/TC7S7su07Boruu7+v63NT9j7mgG7n6taG8enddvLPiqn1mlXAsP/eJ4LEQ91gfQIzibglRAAsDCByOo/wIFVhHmLsnnmnsR5wwd0lzt6kvFkMCQgjhAmEAP+6IHYgGCBzljePJG+KIfDmO61MezkVgoIzstwDchmv5+Qq+c8EPSxdApKGcWH2wWp2N+BQnXPv4Pjd664i7+we/or9xVwUOiDVG/hGfApHkWiWC6XLPvyKxYrV80ecCRXHfFqODeyuTjybAmMhT9ptcvl8Lcs792X47dv57iNWRHevUPldExJZw9V89AusCgbffel/U11OtSIAYjEK3S/EtdjW7aW+9Es3IuuIqrbzfot9Pqg80W83ORKUS3Tc4UB+rE7E5Dhl/GDcYXzrEqFjpTRfuil6n4/+iOAcB9zlKjEn5dj4unAq3UIyJjJm2PUVf7j+f/FZ6P2v5uAJrxjmSuYhi7OY5gtDM2G3CDt95tphLQ+rWx69YyxXsy+YR8Ah4BDwCHgGPgEfAI3BREPCCxUWB1WfqEfAIeATWJgIloQKS3cj1fMX/KgkXL1NeL1YadDt/5Klu07de46rbe1w8HLrWY/vlImqzi3sjV9lSd5VNEjeG2y4cOuqiGMIfkgYCDuIN4ox9PKcoK8ICBA+/YW1hLqIQLHDxhOWBud6AVDdivByvwoQMRAdWuvI3AbUtFgYkEpsR8CY0UCaLGcF12Y+AAG7mNsquw/kQ7OXna5lwtxXREFQQU8TyYB8usCKXTH5VsSqe5U68f4cb+SD3Zatz+f1ZShZ8HMEFjCAGb5dQcWtR9gv+KNqIrQgGE/AEKxL3y99mtcL17J5MbOC+2AxX8La2ZuIF92EkHvvI21xl8Z2N38tiWk7ezb9BtdsLvmefgUfgciHwnk8+HMqCIpKbrd5WO9F4lvXUqnFLgsUOYlnIFdRIrRYFcRi0ZHlxtLdRzbQin0aPOElfYxw6Z1JbRDrxgeYECn2/RQlXeXN97FxFhpJgcY/yMddQz9T3L59rXperPi7mdYsYIjYWMoZSjzxLTBA36zuzbjrner2Y5fd5ewQ8Ah4Bj4BHwCPgEfAIeAQuFQLmQuNSXc9fxyPgEfAIeAQuAwIlEhpiBPKdxAYZn6+g1zEQwhckXECcy9oCV0dPc4f/+EFX2Tbs6ntSV7/qpGvs3e7SVp+beWTEVXeErj2m61UmXdRUINItMy6qG+kPCYe1A8Q1RD3fKSNWGDy3cMeEcMBKXkg7yDGuiZBhAbFNSOB+IYGMHCJvYj9grQCRTv43ln439tt8iZOnWV5YXvzG9Y18N3IfPI20n29RMesyq8C6+I4gYa6dTrjp+3rdyX/6drf/je93yenn6zfIRGJ9IMZwX/+iBPkHLpQLtyF3rZZYUWoj3AfXZUNE4F5JWKZYXA7EI8pEGUyQMIGBemG/ucoCc3MpBA4QpWCaB2wu8uF+LI4I3813ezlguQlSZYsNyugtMIrK8h/rD4HXvPCafNxVIO6pyenW4cwF1STpxAp2Pt6oxQp4nraDIJIlRi2V26AZiRW5RYWlCwjGTB8lZpAFyP59fX+REuPShWyU7yNKP1Rk8jR9Yil2wZZ8F1KotXAu7rgKUYcxi/HPnhN8mlCbP0MuoF7Xwq36MngEPAIeAY+AR8Aj4BHwCHgELggBL1hcEHz+ZI+AR8AjsK4QgHQ2It+sCSBNII8hk3KrAxHX3Qu0tni38vlOpRvdwV+L3c4ffZqLBrEeOOZaisUQVPtcdbjqutO6nriZqD9y4UzmKlfUXNwjvi5k9b358n6evvOsYh8EOH6/EVkg8xEpIL/3FbXAPXE/kNzcC0JCOYipuX6CQEO0IFA2q1vJzwJuQxZxLc41AcSINj7Jw1b6m3uq+YR52S2UiTBcw6wKOJ7yfVpp2mXpaTfyvu3u4G9E7vRnOe5KJeoJ6xHKBbFo1hyUCQz2K92r9P7i3lfrw7AGV4QGro9ggiXKFUrEz0B44V4oJ/uw9qC8JEQNfkd84Dzwx3UXOHO81S1uriDocEXDtciH48AGywzqkb/BD4GKcpm7K/Ky+CXidXP3ZiYUeQsMgeG39YcAgbjf9OdfTK66YrAlC4uom6RBrVZxg321LFG089OTzeyKrf30pzm3aRdCanOuyHPE3i8rfb0S8XneovSjRb89XxAZF3FtZxtxfjb8VggV4FAWbspu9PhtbvwqHZ9j5y1UNnwTuqgAtH48z75sCXnGs7T2tot6eZ+5R8Aj4BHwCHgEPAIegbMQ8IKFbxQeAY+AR+BJigDBjbXZCnXzmQ35C/Fr7n0gwNlYFQ8Zxv74QkQLrfhPZWXx4SK/ne7wO77ijvxJj9v7S5vd8Lf1uKx7woX1ba79aNdV5Rqqc6TjkmkR9fedlDVGw9WuqSjGxZiLKhDXkPVmPWHl26t9kD4mUJRdQXEvFtgUKwCzmDAXUpzDpBz/7+TxeaVnF+dwHfDid1wt8d1Ico6HtCdvygW45DU/5gJ/Q9hxrrlSIg++kyfXBHMFJ3/8Tjdxxw539w+FrnuafDkHQt/KQRwP4lNYbA+EJfYhCNyl9FGw1udqbdw316AtID7YfUJkYnHB7yagcAx/W8BvAqfjqx4xiP0fU8KNF/nwrsF536C0VQnMqRdZ1uT1y73z3SxorL7NMgNhibIQzNeEJY41d2F8ll2pgMdq4kJ+fvMIXFQECoI6t7ZQstX2ds0FXcyVSe3zJLQZm35aiZg4bD+o9OtKd/MH+Z9HvozTuLorb4xr9PMNuy2Ao7cM27Ct4ewb1zuT9XHahX0vx3wyF4pnPdv0HnDem4SK8gIL3pPovzxPTRw977z9iR4Bj4BHwCPgEfAIeAQuBAEvWFwIev5cj4BHwCOwhhAoBAor0fwgn5DeTEYh2S1INc8ACGpWrEMs8zvuQCChsbRonq+lhSbQ04VoATn/XJclDffIm7bIHVTHDd7yFJeebrmgHrjOqcdd6+ju3EXUzP2BhIoJxbnoldVFQ6LGjGtcjSUFRNcjSjcpUWZzHwRxT5lNWOC+zOUV94VAgJUCE28m+WY5AUbPKHDYo0+ugbslBA7IcshCiHTyYPU/BAKfuEAqu/EgH37j+mZ1wfXBGHKdlcsvUKL8lMVcHX3c3fmKB+T+CcwpE+XD3zv3Q164qcIagbKTF9Yg5r6K6+PC5TPCmH2rshVWCogC3DMYUxbuycSDh/QdqwhwIFGmvUomKiA4cC7CBvtpR7Q5XM6QzI0X+HxJ6f7inhCBuB7Bw7k+7rnAgxXanI+VBZsFFOYafKfNcrwFHrb3GSN8y/EvPDFYgOg/1i4CywgDF6UNFy6KvihU/qfS/12g8/f6fLpSLtaeh2hBH8QSy7bH9cVI0bVbAcuUTM+z+ZuRymXCd74rQCOf7flAHgvW5YWQzusW1A1U8FL7KYuPPO/tWYUFKc9Pc0NJuzLx0uJZWewo3inOe0yQSGHvh+THM5hrcQ1rv/Y85Z3Kbx4Bj4BHwCPgEfAIeAQuCwJesLgssPuLegQ8Ah6Bi4oAk06Lq8CE2FwkQcKzQTKbeyPIZyaquBmCsL9KieMsmCvE8HltBaF+mybqWAP8vFLDHf2Lo+6UFt9f8aPDbvB517uwoSDcfTUX1UJXuzJz7ZHNbuqBqut/Zibx4qgb/9Je1/fUcVe/5loXVqtyF/Ue5fP9SuaCyIJ1W3wFyspviA6Q7ZBuCA3zVy2aqyaOZ9IOYX5ACVdLuDBhVb+tNIREIB+uhcCAUGABwW2CT364c4Jkh2zHTRJ5QnN1XZpMuWym4aYf2umO/dnNEisQMLA4QASAlEfggDggX8QLPnH5xL2YCMO1f0+4UlervZlbJcgScONa3A/CBIlyQGJeXVwYCweO5TiEJO7FgpNzH09VQpSgbbFam/rA7YyJQtQhBI1ZdXD/5P0SJbBmhTbWGuAAnggT7KdsCDnUE0QobWtvkT/tlvwQW6gj2m7bYrPou5MAd94kD+dfzK1wybHQJXKCSy458rKzErctp2vR01yglN8Wu0npYy4Mr5z9ntw1a10VDMqm6dMutfMv5j34vBdHYAHCu1x3duJ8wnsuw4tFaEu06EqU+EtdyAQLxq3vU/oLpfO1VGLMsI1nCmMw/fKibQUJa887rsNYzMZYYAQt8x4jjM0qi3GefZxL3+GezTLRxOikI5tB9aVIo1AUbFUacmGwxVWDitzZKSKTzsH6za7PNRkbSWaNxliIOG7PlYuGhc94TSLAs8neyywGF5+0Q55vPENZ4MD7gL1v8Fyk73xVie+I9DxneZ6es5hQWFNYObB2xBUjz3baPYsBeNbau9H59v01Cb4vlEfAI+AR8Ah4BDwC6w+B8iqP9Vd6X2KPgEfAI+ARmEOgZGFhrnsgTyDbmeSyj0/IE0gUCCWLAwHZD8GCtQGTWMhiCPXc3c/5WlmUq0ZkHfEMXqjEanvEgMz1P/Vqt/X76q66c7OY5LaLh7bK4uKY67m+JhdRsrDoiUUjZe70J6fdwPNarr5PAbrrU662kwk7ogLPMLMAYOJvqw75zmQbcpxjbUJuogXnMeHn/vgNcQbyHcIJnMgHEQOXRhBcYMg5Zt3BORa/gnw4B8KKa/4vJfAjaPazlL7mWof3uOn7j7vRj0ocal/lDv/JQdc+znnUDwQBohHCBfEcuJbVCwQF16VcWFV8UqQlQsGqb2o73Bvtg3tDMGHjumAGjlDjEI8WB+Qf9Z17frESeH2jElYYtC3uAVIOYYG6QLzht71FfuxH0OBaiA5YXxB8nOthqUGdEZcEAQLxA4sM2ii42HngAV4IF+A862ZrVgShbiB9yIc6oX7NQoOg8mtWtFA557aCXJq1jKq5NLzCpYF6hb7nK2+zU24wvEb4dEU0dSUMha6RNV1voFaVtdS+O6qH1DXDXW4sHXWj2THXTA+rP9fl8m3WOY+1Wbum4bIgUeV9mJdrZ+XfC1cvNiablZcR47RLc5lmoqEFoy+vyncXS7DgTiRY0M5+V+knizujrzEm8RzIt3NxDaX86NufVULMvEPpFTqfceC8twUEPRPmLU+IXcYqxjFaOOMKmGKdx3gO9oy7e5V41lEuxg2O41zGJfoE40WfRl7wrwS9bkrCxAmNIKly2xL0uLr61Nfn9G7ijqpP7tEvD2qk/BdJJLfoEyJ5m87HRR44MFaZGHJbUTbGdq49JzZezPo9b9D9iReEQNH3qWOzbrXn5/Xah1hgriVpi7covVKJZx0iP+0USyX6IG2SwPU880ys4DmXj9m0nSUE7/wQJa5NO2ej9WLFyd8WS4pjEE7YGJfOsOLw43+BjP/wCHgEPAIeAY+AR+CSIeAtLC4Z1P5CHgGPgEfgkiHA2G7kF0QJk2UIKSahfEIKQ9KwUp/fLPj03GpS7YN0Mb/jF7zSDqK9cBGF1cBrlK5yE3efdu2xT7jem14uESJwPftOuSBWMO7RzSL0NRFPZhTPoqrf63IPFbtUIkbzkcR1xwdddVdV+zLFuSB2AgQVk3om3Nyj+WFmQm8TdAOfCb4F4jbhATKLe2RlMXmAEUS6uXuCLGAfE3gEHz45Dozsmkz6P6iEq6nNLuk8zaVjWo37yF4d1i/RInKd0a47+q5DLhmjvNQRQgXiACIE5ac8XIdAuAg7XB/xA6uSx4ShkQl2L6v5aauKKZu5rmIf5YO45P4oI0QL+IIVQgKrpi04NrFA+E5itSjtB2whLRHCEDLYsKSgzUHasX9vka+5wgAPBC42juGa1COkDlYeiBlgz3nfpQSOHyqO51hIR8hRrk9bRxQib4jgsBD2LrlwsQJCiVvIY6hoJTd32JN1RCoFbpdIUrlJE8mU5nTokFIkovQFkmR26i4H0sfd+0WsTgjtZ6mFRkJgv469TufPKJTN8XCTO5ZMuHYwLBwTd0Kixox+fyRri8xN8nYFVuAIdpDVYGWkugkZ60LoKdrBZf0oEZWMw/QXW1GNAGfjCYQhf9OvaO+0e/o/LuFspTP9zsasCx6HFwNFYkJHIsP/0O8vV0KYpFx8f29x/XPFk3KzKpy+T1+fVP7m4mZB8WOR/mELq/gs3z/jJ2MLIoO522OsAlPGYFzLQfreqoR4DK5mJcZ4BinMGMXxbLgE5HtN/e0LSk9TL7o2CN1osNk9oPRYUFUdRRIEoXoj992yrNiezUhorasMofIPisUAZy8Fw5rMNsZzyvRxJYQMRNU8qc2cIVCVzsm/ekFjPiJr9++i/9sznnZHn7KFEy/Sd8Za3kO+SYlnGmMuff7m4q6+U5+I+Gy0Y55fnMMiCsaJc7FWMpGEfkgf5L2IvOijvANyTfKjZdM+aY8Wu6sogv/wCHgEPAIeAY+AR8AjcOkR8ILFpcfcX9Ej4BHwCKwqAgUBa6tNmZBC5EA8Qz6ayT/7zSUUk1QLCg2RVnYHxMQZcseeDwTghty9YLKsINzv1mT+Lcr/ZUrf4VqHtrl05l/cdN8+d/rTD7pUFgi1nYnb/ppe1x2TW6heLC9iJ2bVHf+bSTfwzC1u6qsTburOKRfvOO4GniZiqi6yqH7QRbGRUtwfGDDx5v4tkLbdE/ebBxdXgqiFEOTT3HnwN6QWxCIkA/tx5wGxC3EOFkauM8EnnxHpK6KH9+9yUc9TXefEcZemQ671aMdlnapcW9XlCuuIxArKyPnUF8Q++XE+lgIQCgg6EGfU1T8p3SrcrN7058XZqF/VM5hwz7QdCEv+NvHAViuDEwThASULEA4ZA+FB+REjECEMM+4TcpB8wRRilrzZOM82BCKEIIQQEyv4jfojsRH827Zv0RewpC7ZqA9zUUXd36lkgguk5gElAphbgPaAfrMGrC2s384KFQ2RRqG7IaipTQy7nqApLFKt8t7phsNt7uuzafdMHbdZ5OkwXUKkaSoRItR/N2bjusfA7QyHRIQNuVcIHVkq6X4D18wm3b3hDhGrktJkZfHxDHuMPndL2O/ek53QEYnbqvxautbDStQrbc5coUFeJSKUzSopdzlVqov8q1+BO+uuq2iTYEe/ZgzGCgyLMFb/m6s12vSPKVHviG1mZcHv4M0Yxgp98qG/HVbe9BELhHvWeLwKhDYWTm9Q+uOibt+mT8ag8xFKuS9cwrExHgxKFDkXktWEYxuzzUKKfG3cYaxgrELIBFvEke9QQrhgrHipEuImhDDWfaxOBzfGGTB+TlE+Pr4n/85VA/cS9cOrqBEskQK1+gxZXKNIqKvI7ZqTtVNeM8GmubGslNWSX7HswIqFRL1/Wglhh3ugnvO+ttLM/HFrBwH1T55FZsXAM8jEM6wCGS+x9OH5yGIE2mN545loz0Xbz3ML0YJWichAW2cMpo3MWVcsgsBsS55NLLJAlGAM4n2PZznjCv2Rls1+fsfqlmco74DL5b/IZf1uj4BHwCPgEfAIeAQ8AquHgBcsVg9Ln5NHwCPgEbhcCNjEFAKXZIQOE2gjzphAQ75DoEG+MzlmUsqqPiaukGpMZs0lBgQz53dXQ6woAwMBr8k9gV3Jf7MsD0iUBUKuV1YUpyVeMDFnNWFHAobY0B07XbxlUr5umnIXNej6b+661p1bXDqxXxYYT1Fsi20uqfW6cPCEixWsexYHJvhMwsEHTCC1zPrEXHRAJEBgIRxwXNltlJGIZrUBAcHvrO7nE4wkShz5pGseeL4sP3pcOqV8ssdc9QoFFp+cdMmkyjgz6kb+SWLGAxD05uece0ewoJzkB7mHwMI+6of096sZWFv5LbdR97QXEu0DsgRCAxwQCCACwcpcCbEfMhMcLL4H9cY5kHAQgrQ5go9zPm2MVZwLbWAAAckGYUI+ZeFi/jm05/KGyyraC/kgkNCWyMPcWtyg71hdQAqCOe0tkWiRrXb7XuT+2F1eLe7UYsNsSmRuqCQaVau1d6lVDcs3/kskQtRkMREJ1adkY+5KWUSkWtm9WQSpCTSzjbWpv1UL4U4du9PtkzAx29LtSqz8xq3NkHuuUr4pxsW+hNamHqBr/EhGzWVuv65zh1xHnRBqFf39cSXqkfqiD1k8AIQ1sGMzbM0SY4lbf/L/pDGNMcVWQYMXYh8WPrgse50S/QHycP4GoTl/w70Z4w7CBZjTx95VYE/bp41T2xaHYTWsX8iLcfmNSoxV1P2/UjonKwuCdGuj77EyHJEAofKbtP9v9Jku4VrK3GaZkEyLJR9aKHmYGEofRojAAoR9/L7Y9tOlH8jDNsbXMzeurlqTGHhVAFUMorqSrCvy7xG2W6rhCPlluc2eIksfR/lJn1f6AyWwwtKD5xfCygUvEliumP7380NgXjwaRlsT0njHQCBjbHxeUZeMBT+sxMhslqsruTDPTRZEYHHFhuBh8S2Waxu0ZsYi+hACBa2Y5yPiBHlQRhtHGN+5Bvkz5vM+uFz+Kym/P8Yj4BHwCHgEPAIeAY/ABSHgBYsLgs+f7BHwCHgE1gQCZcGCySmEMvsgvMz/MQVlMs0klkkzq80hk9mMkLdgyxBhPB8uGmlSEPEQcKxKZnUfK08h9A4oMZk2EvyE3Cl18sSEevTDlAvyGVdBfIfcHnUDz+11O1632zX2TbvanmnX2Pu4rDO2uzCCdIOoZnJeXv0MwWACBYQCmIEDIgf3zXc+WWluFifs45y2S7qa1GcV13zwhEtbt7hkSlEGpkVI1CJXHeqXdYj8nff0usm72m701gMSK2DxINcsP8QPSAWuB7mPSECA7oPCBuuAy7HRLiAraDNmbQHGlI32widEJm2IdsYndcU9IPhAyJjoATHC/bIfgpu2Z6RO+d6IhcHv5dXOEL1gvZBggaiDyyyIGGvP5Ee5SJQTSpHV65C+iCC0ZzbaO7E0+BvSJrfKmNUsLk5ciyIQsK0Wn7UIqblMLp6GFWdin/56toSI52SS30RxtWT0EctC4hkSM24UDVsNQBy7lUU2xaM4cwNhao6aWGxTjUZlilwtMT2usiRuX6iSSkRxsuT4yTlZbjYfVoB/QulzStCxkF9gCckKyTWle80tL2Rp8aQkuxYJmg02BdWdt1fa8TcrQTbiMu2nlF6lNH/19BIVlP9E8N35G2PkPysRvB7BgvqgL9DnOiqfWV8smPcKLTAYp35B6a+LTH5Anx9QOhfrCE6lDTDu8kxho79m88WKon/YynQjWJELTBRDUH+1Em50sJoAg9XYGL+e2Oih6he4e5J1kwtVkxINZ/uS+lTGU4a+tdJtZYKF5YZrKhIxCrBuoe3Qt8AvUb2thhi10pL74xZBYIH+X7Sa/LmIzQ2jKu8y9j5Ttgi0XHkPoU2XrQvtN955zG0izyYEBPodogWigr2jLNYeTKbmGrRens08C8kXd42/WFzIXDjerr951vK+wbjC8x8h76zx21vP+W7hEfAIeAQ8Ah4Bj8DlQMALFpcDdX9Nj4BHwCOwCgiUXEGRGxQlxDFEDCs0Z1f/z67whW4xdztMZplc20p+zoXIhQhiNS/HmT/7fKWnrrPqVhbl2y8I+jtFCFisDXyQf1zJVtpSLlYm4yKF+yIQpVmIMLmuuPEvPCR3TA03/G1NN/jcAdfcE7v6nparXTXh4uFTEi6YuJtYAB78zQSfa3IdyGRbtU+ekALmKguqCizG5OZpQMLEiJt5eNRVhrTKtzsgN09tl3Urrrqt6TrjkZu6d8SdvHXCZWnsTvydiKcMyhmCdzaPWUsFLAC4x/9DiRW2HeHwvjIul/p74RYKQcCsWxAcIBzBifbCimlIDfaDGYQMggQkiwXv5HzwQjig3rB84L7NAgMLE6PgweJrRT60U75Tz/ift432WKblzQKItg7BOX+jHNQlBCf1yUpsyk+56BsfVWIVM/to9xBCC7o4WiDvFe8qiFiON8FHMVd0b6G7Wn7xr5XLmX6h9HxRQ7tUkmfo7xnt/4qOviq8zu2WEDFnSbHii3JT8yO2rPBkCSS5yxu5lXKKh+FS6DFRxnlwbmp81kqAZBttgYRLG4Qh2gdkN66jwDoRyfVkJlpN/AQPGz/pN5CRjF+3KGGhhIUCaK7GhghHYkM4om/9afE3RCMEJ33qQnBn7GMcQmj5vaL8XId4CyvaECUKKwvIUBMGaM8mEBMguCyy87wxtzW0NvotfR4XT4w//25FF55tg4iYK9lm5z9PWCI5xMFQoxAWFYFKE+ASSiNXhpXFmfJGjns50McAACAASURBVHAqyZzjcqHDRihGJ90N/Si3YOJOlhIPzywp7eatyvtPVa5/0HeEi0f1XOTZcCF1uhI8/DErR8DaLrXLswxLCt6paCW4eiIuxVIbz0WON6s1O/Z/6wsCMIssyBshmOcozyjGlkXFq6I/0aZpkbwbURbOQxj5WSVGeNvoIzxrsabC1s7esxhDZkd7v3kEPAIeAY+AR8Aj4BFYAwh4wWINVIIvgkfAI+AROE8EzBUBE19IY1bYQo5BDpFYpccxTKoh6VmNC5XCCkCoTSbFdhxEsrlLgvgxxzLsuySTWJEy7xE5w/VYWQpJdpcSVJBZNkAGQpabFYmtBIS8vtl1Tt7rjr17QOm067spdbt/dqvLPl13fc8YcPHW0EWNR5VCV90BwcgKZSbx4MAkHywg+0z4MVKi49qjD8ha43oxV7FrHh0RG9Vw8ea9buLLky6qN1zYgNo65SbvUfyBeuqSia4b+/SYax8BN8rK/SBKQB5wXeoAKpj7epPSx3TvlwRjXWu5DUzNzQx1AflBO4LkgDSjPgwbhAlWf7KSE6sMs8zAYgQx4ZXFPULCgC++uyFxWUlMDBMEte8u8qZcEJTzN9onpApWNWzkC9lTFjXK5yB8IJAYSQz5Q5k5jzYOicOnCRb0C0S58EJdQ5VECvKmHVH3tC3EiSGt3r5e6RX65WrFnjiulrdbpSFYbyqLh54sEY5NN3CW1cQCoCy1C7dQeWDg89ggYCPJUGrNLpCsBlmbghZ02ZnrbllNTGL1O+PKf1OCBINgRrA4LjzoT+0nmXBhQgVjTkFX5+34e5Xo0wihRlgyhrEhUK72BklK+n6l31GC3GR8JKAzbZrtfElu+v+nlMymgFgLWIRRryvdGDvKNgkIiO9QStUu6NP2/LEy0sIQomk/WHi8ZqUXKh23UrFi9hSVQu6f8pFArtYeVFyKK/RZVY+sMgIqpkumkSOgP+aWTmzEswCd3KZF32nhEvZS4snQ22kB2mQ9NXv3CB4FauRB/wqXtxF5tZ4Me3T1DyqH2/T9Pj0Xp7xocR4tYvVPoe3aOwJ9gnaOZRXvTLSS5cQKSkSLwGKN/oul6AElFjAgUtGyaGG0JAQ/vnN81+p/geD0ZuHFex79h+cwzzusvXi/WGgjT8rPmMHxvKOcFWjbW1Ysgp7f7RHwCHgEPAIeAY/AJUHACxaXBGZ/EY+AR8AjcOEIFBYVllHZ3zcEPAQQE08mulCLEMSQQUxEWd3Pd1ZE25pSo10g06BamBwzySUfPskDYr19oUTuudx5Qdx/WAQN7lT2KnFvlAdykDgItiqR5xdEOO5RmGizEhHrCybtmZv8WuTu+wnRrvFmN/ySh9zml16peBI7XW234gLsbrvphx5w217ZcWH/dsWgOKYYGdcr5kRbwgReykUehDXXPqwIAbUh1z21T/EpFJC4Pa2/Yzd9X83Vrw21BBdaOHRpIso5nXHtkyfc+KcrbuQfoKsoGz7TwZ0yUweQiWCKaAFhcED3a+TiucB00Y4trCxoGxCgUG60M8pqsVEICs4+iBWEhL1KUNoQNtQThAmCGGQt4gHHgRMiBdYO7EPksA1hYSF3Oawgh9CBHDKxws6hvX5RCYsboxJLWeZtmHZdJoqxAvikEuQyq9/pJ5SD+6SMy5K7CxBFdk361Ky7p9kNMhsyiNW2O9XjBkV6PlWE5RERoDu0+lqB2V0zusZdI5Izth6pTAbyM5faUpfJ6mE2doTCuef/tt3J5DHXVP6p0lckgkxnx903BltEdnUk7gSz1KliWOxeqd1GDNXFSnHVvNxX5aJFHh+DlnE2UljaEJ8AcgwCDDdc4IrgeES4QcaZX/RFrVkuNzm2hMsnasSEChOiqCnaF/eOSIFgc64b4xZtFdqbflXkqZpbcFu0if6MDv9IkRd9g0DZFuNixQGcS5YRXJ3zbaNf41IGi7Bz2cqteWdl/HCstkB56LOMjc9Xou+z4vyZSq9QYnxYbptvdVU+nns3aznGYJ4LPNvoA09XLcZq1x+XJVKPxIkeuX56ofYc1feuRMRXqX9sVv8a1b5YFhandfzsaneC14euIYuLcbX/GfWznYr/Igdu+k99Uv0jUBwZpwD2uYUSokYuZnC3hXihQPf5ligiCceq/y9sfRFolIjyMeoWXfUjEk7erLw+q/bJs2PRRrBCl1/LYet/XxwBxnfaA89ynmUseOCd6juVvnkFwNESaJtvU+L5hnUl72xYL/GewwhrorpJxDZeZgs8f2zhAGMSfYpykT95/poS70YLbYzNtyuZC0dEk+knmbC8gurwh3gEPAIeAY+AR8AjsNYR8ILFWq8hXz6PgEfAI3A2AkaeMTlFWLDApEyImYRaoEVzD8IEFiIfgpZJNkQv1COBFnkOQJBxHvlBLCJ2IHSY+HHJ66Ag8ufIfJE1kAX4WobEpvwQBtynBQznXnGJAgFo/tY12e8eV9yLa5VGXRDtkHWFnO3Ep1w09Ax36O0TLuoRQZAqlHHvI27ztwy7yftPuNqmabf1tde71uMDspJouwktHK9uqbr6lTXXOVVxjd0zbuqurs5tuNq22I19bNodfsf7XHuEckFDcX3KRr0QMJeVwxAU9+i+1rx//0K0gMSHSIToox2wipRPVtPTzvjNYkGYCxfaFO3IAm1DVCM0QXhC4CNq7FXCusI2fofwnb9Rz4ttEDOkc/GrDyHK8bSjjynhboXNrHf4vqxoUSqQuQujz3B/WP7QzyB6n62rXKH0HXIJs03E5ox62Y3qVV8vonQ02uc2STx49px0WL5LWkzJUYjI0/vUYu5WS9qn4xEoDkvweK9q5TmyfuhRL56UNcRXhbrcleleFAlDwkJdBOetQeLu1wry7Tp3T3pMBGyv2yvLi70SSabkn/9lymMhP+qzpSnc2OgcF+qoVGQrQbuxuMhb9cJIUa/gYq6j/krfIeIhxCDUDZ+1Yk1URn6p7/QBaoVEv4ZkZ2zCggh3RfMjiSyVFwGs6TtYMNB/LD4OVkPDWRBpnAieFWQJ4uzVWRDy+0yQpRKBTGteEPxvLS76jfqE7CaGzAElxnGE3HMddyD5/6vSrxT5/qTcPCH6UftuicDZuIOioNQx9f6XSv9aMttVfQ/eihhBWbC0+nYlXCAhjZ2r+zPwRpjgmQYpSx/+c6V3KlFX1A/jzUNKPPMQFo5INPxHteshuX1qqf0/U4LEUxAe9NtTBW0rF/YCBajvmxNQGZvO2GQh8YSYZKWWdI0AwRZoJAvGJVY31e6nJZDU3Hb1x0CSbyVTDeBmKhA6mVBI9LQKcT+1lF1IxX2renaklvK27n73wfRRN+6J5fm1snp/LyFa0q4Y53nG885Ev/x5JawCLUbSQgXBopC2+BYl+jwCJ8ITz0IEdJ6zCGt0ar6bO8rlnkUmklMOxnHGIhYJmAUifWux7bP6gYUCuEbk2ozL5zo+LJG9/8kj4BHwCHgEPAIeAY/A6iBgs5/Vyc3n4hHwCHgEPAIXDYGShYW5goK4YZLLxso/Jq+scIesYkIMacR3860O4Y8rHchbVs1DQLGxKtcIWDuPT/Yll9LCYjnwijgXONUg4ZIGAoByMuGGROTeIBQgy1gBzSpfVjLbPXIc+EGyQzRYwHFIREgCBJ2m2/TNAwrgPeB6b9IK+CRzzce6WkertbQdnRPXXfvohDv1sftdZwS6CZyZ/EOUWVkg9ll9CWFGIO3CWchyd7h2fld7MzIV+hq8aW9gDAGDMAR+EDiQuBCRtEXwxzUQ+L9ECesISBSIfIgSSEAIFnBjJb6tqIaAxN//am/Ur7mmgZz5hNKHlSDSaR9YfiBkzPkJtwKo3Z9RlmKFq61qpf2wqpW+Rd9jlS1t6F61gBu1YntGlgm/LEL0OrXME2pxu0Vqsh77iH6DnJ7dsJiYdMfxeS/icrPiWEzKNdR+EZu5hZP2/27ysDsa3ag4F7VZd0v6/Q6t5D4h8aAlxGcC2QjpWm387as1h1rJnUkyikJZWOQ++BXBRcdGuvaQ3N7slmBRl3BypfZUdGS/yvvzlG854IlrkUrihGzNY1ucTXExZiBSYWFT3iDEflqJ1e4mcpn0MZfLGrSwoC8zlpCoYwjy65Vow9+hBEm4kg1iE0GLfkDbQ1zFbZqNP4wf9TRoNNrVqxX9PRgK05lKnI6pfpLniQ7fEqZTX9V3rvc6dKvZoWpJTpO8X6/EmM84dHKlLoWK+BPcl7mMsXuEBKXc+baUaMHvX9l/eHNa6f0dMfSvyzN77795Xf+9H2AMAUMwORehxy7L9Q0/AGAsoX//LyVESIRVxhr2nZIwMSXRLVB7D+R2bbda/I25fBHmQa4RAV+uz4WstOx65/wpq6R7lP/tql369VXpCTeYHXW9spRAnJnQb/S9iHgzuKTSfhfJqZ6JHmddMJP93iH3ofSwe2N2yN0jd1MIxl0vXJxz1Sx5whJiBWM+YwBjJO2FdwqEShZNLLW9Xz/yXoCoxtjI37wP0D55VjC+8PzIRcDl+mfp+WMCKuXZq8R4+31KCIGLbbSZP1BiHOLZR/wKnn247FtvAvIysPufPQIeAY+AR8Aj4BF4siDgLSyeLDXp78Mj4BHYCAgYWcq92spuC2iMyw4IHFbvQQRBMkOMQuBAXpHYx4TZLDA4jr8hayH0IZ3JL2fCRNjmE+m1tBXEP66ISLiOgmxidTFEArEUcHcANha3gL+ZpHNv3KO5OeJvNghtjoeAN2Iicadum1LS/YfKX0LF7HGQrFyPa7Omlrwg5sGJa+MO5x+VPqJyWv7FZdbfB/Uv0cJiWrBSlPZjgclpI+bLG/ELAgbBBjIRPHGHBD5YmECsYM2DSxmI3xcrWUwMSOy/KzCkrSJ4rOZW9qNvliEQsZDOiDC8B5kVAHVsK1wXKgPHcv8QVrQDCCII+nG1nLbSVUrXi4S8Ntyax6gYZtW2SMspWSkkWn0d6/sTYbFT9bWO3ILVlWeY45aKvLxLAsMfZZmEja3qu3V3SCu+H5OocY8ECySGADuK8ErXSk4r9sUzi766gqC8hUsZ6tGEqIry6lP6uK7/aqXv12/FWvGzbz9E3mm5Q+moxM4TbkJlelbeK57YqNOF1ovT72wFPCv36ZP/nOM2S95dNkuuRRoaRCJjAZZCiES0a1y+YD2Fj/qFYq3Mz4q4D7+rhLUDfYP7xgKMMYIxlmQOtuhL01+9/lhQ6R6u9c588VSUjkWN5p2VauexU2HW3BslY61uvPWXo+TkH9XaD785zGa+XlYYIkMz7F4o1/yNfgZRSn0y/t2m+n9c49KKXUTpHMY2hIB/X2SOYIH4sWwexKk48rW/Ssee8brRLFZcHw2kQXsaghfLClxBrWRDgODeEHnoZ7QVcCUf+hEr1Gk7tEysKehDEMO51VSk9eZK9Fn6KuMAz4l/o0R7ZKxBQCpsiVZSnCWPmXUBmLkPqZ8q5pF7NB1z71J/3qXxYFuaSKRIczd2D+vzYdU8ff2lWeD+rUq4LT2gX9QiwoUo8MCFsgp5hYSQ03L19nbi30i0OCSMT4tsXrYuLvjONm4GjAG8R1gQbMaB/65UDmC9EDoI9m9XYiykPf5vJd6zqGXaqy1qWFRxXML9E88eLBLJhzgv9HHGqaXECkS+31Ji3P9bJawrcFDG89BbVmzc9u3v3CPgEfAIeAQ8AmseAW9hsearyBfQI+AR2OgIFJYVZlUBYWpunBAeINH57cVKrOpnIopbEAgdjkOowCURk2T8I/M7+yGGmcBaYEfIHhLkOyvlWyKsl3NLsGaqRmQcE3mIRMg18OBv7h3CAXLKBAzub3Yt+uz9c69gaO4/IFEhtCCyOBaiCyw51shVMIMwgMhA7AEniL2viRA8FzdFawa/pQqi9gee4EEybPkOjli5gDVtDIsJyFHaGeQO+EB6QvrS5vDVzepqyF9+R+SByEEAgnSEwH1x8RtF4m8IlQshFalb6pP6RkyCAIUwZ+Ur5fsTpQNKuWCglJUtiooAwfQd2g/3QLnJg7Kxyp4YFJPqXV0JD1uFxF4RirslMoyp1dwgoWKLWkon2LzIavJE1ihdBdVNhFkqcqvpvph13F2ywgiUD62Pdka7K6+CXbBfnosPe/UXe//jk/uDKsUahvGFIM70mYU2vPnfqvK+L/msa6QjImKT/NzvXuT4hXYTy2WWvJ0lmhGzIPaWEovcxbbAKDChjsGDsRVi3ayH3qjvEIXLkZW0K6yQuB+EOLbPKyFaMNYk81dSFy6UOI7rMg7V2x3FxcnFwqAnDmaqtfRY2HY9US0bz7af+q1n9E1/el8lOX63gucMBFnnF9VsZel0VrMw6yIISwjUv1DK2/lSq7lLFhaUCSKU8rP9kdIvKM25wFnIykJ9BgwHkp7N1xz8gff/anPHTbm7ql1/95Nu8GvyiJVroMtuYIeYSdtnbKHc4Mp4AtFKf0QoNQtD7jUzq4OiLmnb1BnjEn0WN3O000VFOf1msQNMmF22oMUBf1iUi5XrWJ011Jo/oDQqi6Tp5CHXSffnZSZfymxCy/eoJ75RY0dvHpBbo2m4WAsTbN3P6Hldc3+QHXN3y8rpdo0KYJLqvlcE6kpvZiMeN8/Cgr5IXWHBSfulTnmOEXdise3Xi7qlrdIOGDtMrGyv0IJiobwpi72DMNbyjKWzE6diOSsPBOo3K9FvsEb6gBLP3Dxuk7fS2Ygt3d+zR8Aj4BHwCHgE1g8C3sJi/dSVL6lHwCOwcRFgwmrEOatFbXW7EajmTRuyHBIZIpbj8V/OMeYaCUKSFe9MYtn4DTKXFeZGxptrqPWGNvfNpJzJOVQvhCs+nZncQ9hBOLCi1oKQQyyyD2zYf0dxw7jtgPxhUg9RhrADwQ2NZOQZK/RZLU1QYcQLSC5ICsrwpNsQrrRBcECaQwJCtkHmQBLicoaVpNy/EYtgRx0Qy4C2Bta0RwhGCBZ+/5IS4hDY7lWiHbJ6GrHNtqXeUVglSt0tt3ENiHGOp53zN+W5XYm2Qf1Rr2ewvSJdTSCkDKxg5X4pP32IxDkjOqqjO/2SfNFfKfczqaSVFwqlfvWsL4XD2idXNDr7Cdc3Cgev3z8vNLYIvfdqpfStWoE9JRdQ3TzYb13WGFvmiPs5An85sstAeNOff9HGguC6PZuzBw+ezF7//c+Zuzcjx4MrBzK+i3DmGqnIOsjhA0qUFVIaywDu8b/MAxgrj1fIW9Y9ElU+HLDqezJ3LfdOpZcp7VVazrUXx5Goe7O8MHEVjC+XixLqnLYMhohkiGus7GcVM8IcG4IvxOX8jTEGQY6VzLhngRRHjOEeT2DZYELAl230PTMH+ket202HkzQdmG52sk4nmQrDsBFX4igOdw9qoX3vdLjlWGfoF/ZvqT7l4ah18GS3emW67fQfXVlJjr1RFhfK4oxmbNZFCINvVYJAfYfScdV3Z7E2NS/4NqvF6ZdYsP2EEkQs7tvOUkfUZ8xVDdi9MOi2dgTdmTkLp26voJXp0BIbwiVu4xiPwZPxBGEL0ZF+m7fV4tqIJpZZ/jlP0LI65N4RXW5XsnqZXwRzB0f9M0aw4TLqz5TIB+GK+2CsQGzj/hBCEAuwbGRsZLEAdc35PGMqOnMUyyn1k6TyS3lZO8KIcptYCJn9Yf1yQuNAohH02cmd7j9ksovEOuSsGDcqSXS9YmI03Xcl43Iv1dIzLlTfS90p5cs16TuLAnyxBb/5oK7Tv6mbXHBTQpzm+c+7BO8FNgYsdGuMge9WYqygjmmvtrDhLJFyhdjYex/PRoQTxiPaMuMybXkhy6r5WVvMHJ559CXK1PJCxQprwB/mEfAIeAQ8Ah4Bj8BlRcBbWFxW+P3FPQIeAY/A4ggUlhVMWo18Qaxg8gppY25p+Nv8guOGCMKH32CvmDzzG+dBqkDKQ6KZ731WATMphxCC7DAyJXeQvp4sLOajKEIOwhziE/KrLF5AEoENRORLlHCbBZFnK2pZvQv5jvjxMSXcGUFWQVCVRQpIg1ik35pzmzUfi9X6u7C04L1hfrLVn2Z9ASaQPhYYm/1gSn3ghgksaZdm5QP21AFkH+Qgx5AHghL1iECCaFDe3qM/XqVkBH35N65FfuWNvN+lhJsZhCXKdECJfpFbFBWfTbX7pLCsoFyIfxDUlIN+QwwYVqpCUCXKZbtWRlflf/5FSj2662tE4CscgdyCDed++rUIXqJNJgsKIlgE6r+ZVt4HucswSE7aFCTSabUlWy0+r+izf0qMWHC/doI1Ka1V41zkGeyruXotrkxMtdPdOwaag311JxI8qFaidPNQT076ipg+g9wsVhibiEnsG4SlFyv95SIX/rxq6SfS47q/1E13PycBKcnrHLLvh5VercSYAiG8lGUC5fjtAlNIasQTW+l+0WNcFKvxrQ2ympqV+Fh9ILx8m1LZrdhCUGC9AEbEuIDQZkylT1C308u5YUI4mml2auLyazOtzpZOkl45MdkaDOVOLFRQk1a3e7KnVtkVR2FPFEfjlTisVSI3IqOe8Wo0M7779FuvGJ56/75qcuSmIOvKt/6SogD9hrJ+TmlUZVtQHJpnZQFR+04lSFjGzx9X28mtLAphj6/0Q+6b8ZL6fm0WRgMjL/ovN5245f8CQ7flk7/ptt32poUsLP5UP9O/qfdPK1EmI/7nAhGvlHAv6pP+z/MPKyhEC8Zr6nb+uEDR2BBeb1P6RFH+b9EnQB5Q4hnCMxJLE56Z9H/GKNoMZWW8QWABG5tX5XEmhO9c+13AzQ/XBTfGF55Ru9WLXxZudz8a7nUDcvu26JaqZSWKQJB1tWI+cL+n3oJgQZtlrKTcZ1lcrBS/xa/65P6lGP+sHWOVQ5tBqPspJZ5FC22/r520GcZLxi7eK1gUgph1TkLFvPbB84a2Sj0ilnyP0gGlVyghXPAMXWp7VD8ioJgLKNpmbrHoxYplkPM/ewQ8Ah4Bj4BHwCOwZhDwFhZrpip8QTwCHgGPwFkImLsWJtGIEJA6TKQheyFQID1ZZQ7hAanG7zcrQaww2eZviCXIQia/rACFSIGEZcU5xIatXIXEN+uKdSVWiEin3Lmf9AJBvkN48veoCGjIg3zlrEgJcLpORBLkwsf0N0QRZHEeFLsI6j2ovyGR+Rui4sFFSMcNI1aARSFgYW1RdifEd3ODBbaIAXyyH3wgSYx0hPCn3ULG0Abxhw8BCNbQcxDkrOimTdN+IRtpo7RVEwxoyxCg1Bu+7SGU5m+IePM3CBxb246FBMQSBOve4pr0jZzkK0hY3o8ghSgzhCWJMpBPR3dH4Nx8k2CxUz7m9yjANoGtOeqA/Ng/RcdQ9lPai4UH8SwgNSf1yf1AzIIFRGOrTGwuUPZ8lywlFvxJQobFEpkWyV1TRfWlWVaVWyER3kF8eqI52mwlba3c70xMtdoHD49lR05MLMZqU1/0Fwhc7pcyy+WQw93J/O0bdMQ/KrbFz6uWv6xV4ePJvarDdj7GULcfV8JNG2MPsQsWC25MW/k5JSxeqAdW9COsgrWtGl+ShV8Ms+X2F+MBbZH2hPUPMSpeq8S4uZgFj5XlN3UMK5cZOxiLETkZT0lsZ5k8LFaebpr1pGm6aXK6s0OeoK5M02zrZKtzRdJN03Y3aU1XO7t6GpWkEkWtMAomJDwdlZjxsKwuDgf11z6QdpvHdky/62jkuhqvgm9eQrTA7z39A0HlC0Vci7PGsXlWFvRLxG6woY6wQpksWSEhUJEnYuNLlXg+vSZQ4IbGY+gis1tnADjPWCf1Ee2gx9xeYIb1ClYWfJo7uMUgW2o/eSJSYK2FldeLlskEJZC6oxyQzYxnB5ToVxYTgzqnLXID9A/q3Z47ZE9dg+Os2L+CmDJFmRhzyI/28xj9SHFuPpM+5n4qPeZeImsrJ/HirC2kFoRQekQWXbG7Nz2q+pmVOxHJ6H8+PsHZsC26p+QOjjGKtoO4xXMJoWAxsQJrJRJWNh9VQjBCvDonoWJeocpWFQj69D0WVnyn0mJu+spZmFBBm2YMYzzFRWMe68SLFefQKPyhHgGPgEfAI+AR8AhcdgS8YHHZq8AXwCPgEfAIzCJQWFQYHOaSBtLQVv9C/DFuQwpDdEKoMEEmQZ9CEiJSQF2wChSR44ASBAwTcMQMCGFzewBJYgzSnHuN9WRZUYgVYAYWNtk3Ai4noMHV4hIUwgNiRb6ZMFH6G/IxFy+K3+eOtX0b/bPUPvI2I3zzILdKJk6w38QLvpsvfRM3EA5ox7RrSBXOg6Cm3SIk0HYRMCBfaKMQ3zhJgRQlX8Qn2vYnlRAdsHowMhzCDgKaT6xnyIc2T9+AGKQvID5ARO4tzuP6tjJ5rh9oH+2JvoV4AkXIKlVY134R9Q9pBfQ2+Z4PJFTcLfr3OTr6OqGwKehFNMjJfgQJrgOB/UElCFqIRO6J34zgRBijLa54K1w/mfVVTrhHYZhEUUj+AzPNbm8ch4MivhvpVPbI+GTrVDdJxyan29bf5669wEXBADyojwNKrMoHcy2Pd8+Ydzwr6n9ftfmG6Ab3KRGp+zt/n59L/dyuxDhF/VNXr1OC9F5sg5Rjw/0J10R4RdwBq1V1t1YQlIwZtB/GReqX61ALtLOFRC8rN/EVWL0MyU2boIy0ZdoWq+oz8l8JaY11xYFDp6r9MqFodrr9cgO13QXZsOpqYGamvSOV5YpEp4rqUyv6s269Vu2EifpLlm7qadR747Cnp1m94fiBoddPTtaffe/eid/8lUr3yDvCdEauY9KfWQRoRD76Xd42VVYE26XccIE9fQBLi38Okk69iFPBswZLA0QBRAsEC8QB+l2+he0nQvp0B3djtqfby38CO/KEFKZtkcza6bwCSes+rD8wRlAu2hHjxkIbfZB7Roh5nxLjj4lPtF8rA8+QvM+sRFRc5Fr57iUsHLgWVl352KCYFx/UmHKX0reqF02kh93Py3oLEv2MLdSafqWh9EH3ixI3GK0mJZe8XOmAeZZC7gAAIABJREFU/qJtg7F3/7NUpTzxG88j2i0iAW0YUZz3LcY3NsQILBts470AqzBErE8pIUo3l2sji1jZkCdtl2cG/cieQVgISXx0/3kFt0B7fosSfYh6R3hDqOCZl/dtb2GzAhT9IR4Bj4BHwCPgEfAIrCkEvGCxpqrDF8Yj4BHwCOQIQJCYYMFqVQgYVsQyeeYTwpeJKaQEpC6T0hcoQc5igcFklVWwkDYQcRzH6jzygZQhb9yX8AzgN/KClErWoVhh7rLAhQ28IH4gZCGC8nWnItVT3dtSpFxxuv84VwSEawHxrH5RtK+chCu+cwDfzRWTETKQPbQ/CHcT0WwFM2QqxIsF7oYsol3j0gkf+hCRxBCBLPoRJVbFU9eQyVwLphTCCSsJIyLNVRV9gvaCkGHiB+0m94vPKlQRS7QVc5EGGcTx7DskamlYvuQPhXvcoCwprlIvgrw6rjvYrAQBjqhB+VktjhUIZBcrXUnkxZavxC6+n+9H7gZKqaMqGFAbr8pl0P5KFEQiujfp70onTSpJmm1KkvRUS0v1iwvlWEv06JTjWyxQCPK2oPImWPzVAscx1vy2cHmzBJwPVF/rPtd+d44d931AydxB/YO+X6OE26ilNghDErhyDtYon1edgCl1sCBuKyXkCmKb+tyrRF3h+glyD7IQK4v5W0GsBwhp92ZBKAuAqNuNtt5T6R4CIwjufPW9iRQrESvsIrJ6Sccnm6qyoN5pd3erDndpwNqifrWlUglGVXczspgJWh1XzVwnqkShS5O0nqatvp5afKXEjWqj3vPYyb5XTXR6n3XXztNv/fLgxAc+F6XjYPe9Sj+5wD3hAx9x5g1KtwoTBL4z4lqUAmoTf4N6/2FZTfSFnenXz+x61q82Dt1B3yIPSFWzUDnjUvHUCYkWUy6t9rrmtq9zaX3oSDQ9ggUNK8Cx4kEkol+bO7QV9Yl5AZK5Jm0aAQXSmbrAuoIxYaGN+mTcgCDmE/duB5QQFheyillRmRa51tzuJVy65eX/jScWD8z859ufc190hTsZVNwLJQffnc3IKrCRj0FnbblwwRvAjOvLptxHdewX1EvoO+D7V+o3J31Q7oVrpxAuzYIVgYB3JgvmbmIFJ5fFCt65aL+MFwiWiOwE1T7LDVf5qguIFSYem3Us9UvsFERhroErKsqz3EZ/4plIOaw/MVYuGdNkuUz97x4Bj4BHwCPgEfAIeAQuNwJesLjcNeCv7xHwCHgEzkSASaxZCkDmQqRC5kC28p0E4QcxykSXleWs7mWyDQFjvo8hR/kd4pBzLQYAxzKZhcyF3OE7hBuE/qoQM5eiQgvLChNcuCdwMUIWkpX7ZT/YgcOUzuE+u2ZtcSnKuZGuUQgX3HK5HeFCin206/mEDvWS+3ov6ohP2j7Eoa0Upa1zLgQcx7KaHWGO+qWt07bxO5O3YSXijiBymDUShDTEE0QO53Ecv9O3WBVrQZ4XIpsQF2hXlAlCuyL3R4la1Sl99smSoq1fWImPeIIVCAIF7qZYiW7CCnlQZpKVUV8veKNM9g6newk6QRj0VuOwIddC/z975wEgWVWl//cqdZwcmAEGGhhykAxKEBVUUBAVE7qKYXFXd3XddQ2rKxvcvzmtrgHMIIKKmBUDICAiOefQQ5icO1d47//93rwz1tRU5+qZ7plz9VA1VS/c+93wur7vnnM6SuVob8WD6paHxSoR3plSuQK2eD1YmK4knI1I1MowogWdh9CEeERb3i/7RJ3a05eEjmK9uUeiBa+ERukVUQf5xjoDMUz/IFogSLxjGBQIxYJxPG0lPBX1qE64PCog0xBQrJ1cF88KSD7G19kyRNx65VcaAtfJT+vkIMxUorD1qjAoPzxQ2HtjT8ux8azjrrR1Z0zrp/oqVLLt3EC5kg0jCWDF6NA4iNtiCU3ymJk9UI6KSnvfrhBQ5YFiJS5nK7G8aXbp6S/19RZyvdPbmsrtrflQHjXd5dz+xa7S8wZmdv3UQpoxxtl/Xy+cDHPkIzJyR7BmctxWeVQI/bT8lgsf3XjQyy+uNE1/VaV5xrP7Fh33QMvSO5cEcYWY+jx76pZs39pg1i0XBb0dJwaVltnry23zLpdgAbmKZ4N5+BVHGqqmjlBh92UtwHMKbyvGeT2Rxo5lLfm5DO8fPK+SMG+jEZkGa+9Qn1eHdNO8M7LawkrRX8yhRFT/1Cm3RM/pvGj1cc3f/0NzoWudVo4urURv1EhlPdqq5ERzR4zk/qBJrydF6xQqqqT5EiX9/hv1Ie1krfMcBlvDx/MAgevtMsY/AiueFrWFecJYQbxdIuNvLKQinktjmfuMWcYB90cMZf6xLv5zvT6u8xl1+YKMNZEwatSLZwyCnG/OGCGIfpgj4Ag4Ao6AI+AITF4EXLCYvH3jNXMEHIGdDwHzrKDl/ACGzDBhgveW1NNCyhCCgx/XELEQGfyA5Ucw3/OeH9+3yiCmLJROZ/pjluvzQzshFmVD7g6cpF1BmyCeqT/PMwhHiGnahhiDmEP7aKdhC/m6FSk3Sdu3Q1SrxgOjuk2QKvQLJLoReHxv3gcW390SGPM5/QshyY5wiB7GPUSN5SxB7EA4wNOIccExHM+9CO8EwYT4wHF8x1yB4GFMbCadUgJ1QERfUjflZ4jDOUE5M1/zLZuMK8YeSSXYecvYYzc7hDy0IfXhXrxCQkEGjyeuuU5Pkm5XY2QCEO1HvMHm9RfLrBcHiQCfOaD0BxIsDtAOfNrI99TFRCIEhGRfduppMdT8N9ECMuwiGTlzINXq/Q15nj6HyAOLZOc8u7uFI2Qpxn0RHgiP9TPZx2UIB/UKuNF3xJFnRzMkIaQ0xCH4jmrNEtnN2ohXgMIlJbkWSJTLLmn+TUkSSdcpItejpXHY/HUJFmD5WCbq6W3vvX7cffrLPz4UTG9vEo5haxxFzcpPIX0pJtBYMZMJ+jNhnJeM3CThIttUkASliqg/lUQm3EWdEpeiqFAqye+iFBWz2WhuOQi71zS/aG3T7Hd1zl/zua5M3GdCtcXhP6+mfdaX1+nzXwqj+8nnk+anYIwx93Lz//Cf84uz9oq79zkVYjUemLP4XIV3OkB147k0aAmjsoSKWcuKc/adGZZ6V/ftduTtTaseQDAAxyR030jFikFuYus6r4wtrvnyQY5FRGT95/54VuCp2DdcUvSh2jfO75iLzF/qzDjnveX4CW7s+NvepwtHdZ8z8323tsQbClrBipq9LxHieIhtVZRHZ1NhddJMiVcGh8W9CiUVa5d+HHxVnzIfncxOYUo9rUALkZlxzVxAqBjst/EX07GD0MXzg+fIWMQK25TC32WsP6xLJ8nwiCEU1UgKIfYImdcXhdnuSpi/d/n0g1cuWn8bgtSo1sWR3MyPcQQcAUfAEXAEHAFHYHsg4ILF9kDd7+kIOAKOwOAIQGJYiADIJnZw265zfiQTsoQfpKzfELIIE3wO2UHoFHaYQgZBXELms/ubXeacw2cQduzGg7jgs4SonQpeBzU5PsAIDwoM4pm22Y9/i9ts8fMhqy2Ja07XcS+LwcffhH1T5YFRfQ8TCcwTo/Y7SGvzTGAeWMgoiEf6nTnA98wHCCB2FPOeMQARCHnO93wHOUWYIq6DxwNjwq6fhK+qnQdG/qRkNyIYZCHEFnMLkovzeI9AQlsQUtjNbLteo5Hu3B4iZIyRslyfcc+/bfwzf9szmbCUy4QbtQP/CH25RyUK5jBf9H8INch98gxA1NJeEzz1dtM6onsrUfAxQ+0SJi8D33MuMf+Za+xIrhZRWIc6ZJ+WfUb2NZ2zjvwIaZgt7mehwqj3n2XvkSH8EFoIEYF+Yy5TIHGtfCx98xW9XiWDYLcQPpsPGmQHPnWkj/DWof8QeXnPPasL46m6sH5ADLJWPhhnmlfFYaGcK6+E5G4YKaiE6GE2GxbkHTNf/ZWVHtGnHBVzM7ms6h2W9F1LJisPgDjoLlXi3nK5MkMjtbm5KZcpS7HoL5Wa+4q5ojonF4fluLWpLbN8zgdox4oFq/8fY/17MkQZCPrzatrIP8EBW6Qe/nr588G9lXsTEhVxqEPWlhnoOnX2zRdO7194+IbcxqWF0ow9DpIQERDyaYjyO3ljXNS/8FlvU0ioE4NcU37jQWcvmXnn95iTldEKFUN4V9C/jGPq+zlZdfie6uohIHJvvKF4bvaOdG4O1cjRfpcKj+YdyJpkggX1t3nNPGl6snhk5ZK1X+0/e+aHbpiXffwxjbpb1Efn6qgXDXbfjFZArKLWRqxy3cGbFFZqnc79NP5hEqOYx8n4HW0fjLatk/H4NAwU45v1hXWbNfEnsrek46hetRG7EFxvThD9q6g+Gs8KW8cRATGeJ4imSE3m6XTokJiFWYTx5iibv6Y/N+3HfYU5Xeva9iw+M/vovpvnnZ2Ihx89pX64wWoPn8nYL14nR8ARcAQcAUfAEXAEahFwwcLHhCPgCDgC2xmBqpA5/OC08EYQbJAK7NiGYIOIhXTkRy4ELKIDpB0hP/jhzS5lSClEDog3rtUpsx/J/MjmM+LN82Md4sYyoo7mR/d2Riu5vYXM4hmGUX92jyPaQCrAoiHMVO+gh+C2ZNyToQ1ehxoE6ggaSagdzQ8jxZkPvGfcQsSbNw2HkY+CsU2ByGa3tYlZkOOMDUQLSFs+hxhkPFQnn647D9KduIgUiIXcn/HFNa6VIVAw9+xzvDsYa10N3rm9WdjRtRn/zHmI/WROK3zQ/HIczI7iaLHEC4VQCmlrl7Cj7RChRv5bgmjqyJwxshdsR7IOIPKQEwQcIfkQHIw8RcSgcO8Pysgxcl2a1NnCJqWHbBY/8JxA4FHYpWRnPOIFcdtrk3vbeaxxrIfUHU8L5nuyy3kIsQJyEKy47tEyPNOIFV9bWCNNtLhC7/k3niAIJOuzlfUWZqXuvUaTNN1uTDiuT1x+hyI+BYr4FComVGatIvOtjYK4JUvS9Eq8SyarUE+lSm5jsX/XXD7Xk8lk+pXDQppGHGU1isuVeEZPb3mXnr7yKnlklJvmTiv19BVjiRYVCRbgzlqP8ML8sLBlW7c+DvaPB5J8FHtqdM+WlN2uXuL5Ql/Mb3vi2oNbl9zYUpq+sHlg/oHxwC6HVnKPX137O+J+Hcuzivv8MNu/MSy3zS/FmWxe3imlnr1OKYkkb1S4GpsHjAeejSQZN7GCec1zzgohqCwk2VL1FeNmm5dUrLANCYw15qblzUC84LllQis49q8sL15+4erL+18x84OPH9j8ewQ9kmv/QXaMZv+rBmtEFipcV46R2/qCf9JVpwv5/5Icxt8OYFeWeNE/VXbkp4JutUBK0+PREPHpWs64wBuT1+fK6A/es/bUK6z3hB3Ew4v1dKRr5eZrCWeuz1zhOcQmFAvJyZqJyEYxT6+t6xBmVmpXyZUS/n4YhYWZfS3zVty995vWrJx7dNiVnZXrC/K5ppJi/2XCqK+/ZM9JsBnJmj5Is/1jR8ARcAQcAUfAEXAEti8CLlhsX/z97o6AI+AIVCNgoQL4kQnpivgA2QaJwXtIFzwo8JiA5OBHMAQTP6KJ884xtmuccyDp2CUMmcsrx0NWIHhAWOJpUEskToUesZBB1NXC1UBUGQkBdhACkAPgANlM+AaIIIiqfojcqeBVMhU6Y6LraLlVqlwwGLMWTsoEOfoXTwL+rrEwHRxjIhXjnl3VnAt5z1ywUGgcQw6XZNexEd9VBLTlsYBcZCxBlEPIEmKFf5twhpACuVVu4M5t86awdkKu2f0gOLn/rsJmL00EPD4O3ZQyJFYb49mpYIFXBAIooeMQWPD+gLxm3XiU+nLGKArnIQiBJ7v36+32tlBOhKTLCtMkL0kNLtS0R2QeaxHzEmEAepU2YdVJb616ENPYK2W4EbDjuDM9v7oJhhf9DKHNtSAH2UVNCJh6BQIZ8QRPtW/KGB8WOovwTw0vmwjsKCyVArlTxJXm5pzyU4T9pWKlrFwkfXKyaMllsmvCXGamUqaHhZySfVeiXN9AOSupaVZbU0EpLqKBUqWyWLksNoqwHCiWKkneojY9OVK8EVggulktP6TzEN62zkMSBicrafrJmV2DRxRKaHm0RB45lcQr6QJODcvFoOWZW4LuxR8M8uuXhMVZHbm2ULx3vIWzCf0N9tRhiXJW3F9pnc0z6n4JFuvjXNPuSuAdKqH3eIlU7kF/QepDAPNKWB0r1WLFpWl/IqBZaLKG9+UIL4hQwDOd+rL5gHliRDbPLIRQsAN31jEKc3fpj9d/rOcNs9dt2LNw2zVCmPXnYfXPctHtCDVbF11VoeySURxJ3ovXBG8hv4Vm/Z9STw3WsVs1/1gfRu3xMsL2jvqwOp5mNperPc24bjQasSKtCGs52J+V4svfDO8dpJKMlS/LECrwKuP5wt9Ooxq7aXg1xuhBMvK90Mf8TaY860m+o8EK9/qexL5ykMkr+Fvrkz0Ljli2esHxTyxbcEKhf3rHtEpf2JqVnj8zE65fL/865SqqFPLZnNYAsCoKy8Sz1IWLUQ9DP8ERcAQcAUfAEXAEJgECLlhMgk7wKjgCjoAjkCIA82MCAj80+ZELuYRAATnDrmaICghWPC8gHSHv+CGNWMH5kIicR+gTyJEk1I0MwtYSdnK8hUiaiuAbiUubwSAhbWUQO/zIZ28ppATEAJhAVPI5WEAqQ/p6mdoImGhVveOWvjVSi79vbCcs7xkL9L95VUC6JzubhxLt0iTNjDGIJnboQ7xDKDK+EAAQCiG2IP8IOTPuvAZV3WLeD4xrS8jLa5I8Pr1vh17nCIxdM2G4uwSKJL+GXjmHNkN68hlzpdqbAmGF9YDrVQuAVbcf9C24UgfWI4hwckz8p6w2nMnfpPe9XK94UjwpPOsJpFyvt3hZ4rmBNwAeEL+REa7llCEq9Hx9x7Xpi6d1Prv3IedpJ4Q1a8JhMhLqggH1HUys4DbE+YfUpo6IOowny/EzRDXG9VVG+SdCeU0oElQc9fWVF8qjYr5yj2SictwWSbEo5KI5EimmKcBXc29fkT4lN0mxXIrzlULMeB5Q4ouNvf3F1RIyupsLueLCedNs3U/IVWETKf/KusyBwZ/DWcGMsEnid5g8O7Yq4exgX+VD2DdeHZwUd+k5s5mejYNpD/wsWPOcdyehoOQvEUS5Jr2iNyV4fV2GOICwxzPmyZ69Ti7G2SY9k8KX6d8Q9dXPpbECZ56I0PH0MyI++QUokO/0NQVBkXHJMZZLpqeBYuKo6i/ymHrnlY+kXf2HuLhAA7VZ609Zfc98nqbRy1xmbtl4NY9Lvn9G4aEAe/2HFhzTrf5bodl7l/rnKb1HVLJ8JVvWSzNcIlQQq1fkQcOa9WL160k6D48TxgleV2tErNvfBXXbpbm1TYqJEIN5VKgSQxLwQ3ha8TcUAgGbGBDRGIusD4OVv9MXYMRmDwtLOKxYkQoUXJP+5nhEqbNlL00/O1OvPC/4O2Wwwvr8bol8i+Jcc295+q5Pdi06cdWyI948sCq/R667vzynWAlbM01B1BwpyU0+11qsRMX+gXCj1oUNrB9aM+zZWO1FuE360G/iCDgCjoAj4Ag4Ao5AIxBwwaIRKPo1HAFHwBEYPwL8uIRAtDwMkGX84GXHMaQiwoXtLGdnJiQqRJ/lr0CkgMzgO96z4/ya9BhICsLnYFvFfR9/1bf5FeyHOLhAQoARZAtEmWEIUcuOVQgDSEfDF7ICDMAuYdq8TA0EhsmBQegoI8Ppa/qX+WPJuHnP5xZ+ZaRhPTgO4htvJcLjQIgmxKOMucqOfAg/5uuaRuY2SOtL50BWMtapC0KEeYfQHkhK6tGq9k9PxJdYSZs3kcPk5GjS5xbyBNKNY1kfTOxjh3HiYSKCsCKycKS5GZhXtJnXu2SQe9+XQcRWF8QM6sl6BPFn59QclvzTwhchVrBTH6wh+v5DhpcEbbfCscfLLpZBliM23I63RqzZHrYn6yB9xtxHqGAXNYLTYOXX+uLK9J7gzRqBEDVa75MhblH3q0Skbi5kN0qxWC9RYmM2DNdk5FZRKkYFeVkUlGI7I5QziozWp38H+q6kP96X6sSuvoGSIkkFCgYTI2KU5V1TaW0pKH934mcTp+Qp47UQrQya4o1BiwSL7syi4BsaIbcocNjLwpYEqy1KQnBrRa3cL88UrpTOrPzGZUHzsjuD/gWHBr2Ljg+aVtx7c/OK+y7UEazBkLC2FiOQlxf8/bfiO576AsmELak0hDHjcayefZyLQI3wdLLszTKejVZMrOCeb5AxBsD4Mc3N7bbeV4sVqsss6VASoJK6tWhyTM8oOUoljnOxQrmpP9eq93o1b5mnzAHqz5xnHiUk+P8sv6Us0WJTeKhQ8y5WyKI4eKe+fc2WPfnXf6mfg3Ba0ByvkCciVysLt0qAqPhJGd5NiDp4EzBHR7oODHa7cX+eChcmEAwrFAxyQxOwGTf8PcB6x3pO+KWtxn3VNRBC8WhlHCdhoEaytmu+0T/mMcNGE5DmlfsiEJrXGGJFvfBseMDxPEFs2z3O5B6OCu0Pr9/zeSuWHv7Wpr4ZHfOK3aW2vlJptrwpctPamrq1usfyqJje31cJlO+mMm16YWDthkpFggX35u+gXLq2j3XOjbsv/QKOgCPgCDgCjoAj4AiMBQEXLMaCmp/jCDgCjkBjETAiwshISPhkB6YMwo0fsJaDAVKBH56QNhB1kIXs/obcMLIGgo4fvJAOfAaxwXnmwZG8WqidxjZlwq9mBAQ3sl3mtA+sIGp5j0ADRpA9CDv8G6LWPFHAlOTb2pS+KQxQI0pNUnC7ZLUHQPVtNhMwgxDxjajSznoNo1itb223OXhU4z4kCZbu1IeAYu4h9iECMC87ZSSMRsCwcQapNVHkdkI4y2iPCTBGYpqIyTHTNQZZO6gnbbNY+XxHMSEHAo3vzMMCUsvWmNGMmcQzQoYYQfsRb2oFC65Hbgp2DDMfLe/EYNibwIhYQL1JckvYKdY3RBEr1J85fWL6wbNEDZ4ZtgaZ6KEgUiicmfp3t67APd8qG0qswCsAohYMINxZH7CGrQ2DgUqoFpGJCA79Spq+XnJEMqYkTtCvs6RPNMn7YnmYiedHxVi788OiQCkH2YzUqHh2uRz3asd+pbUp09zWUpjT0pxbNSNXLCz4/QXlRXd/wzxzEAt4DnTHkqxEWGfU8zdkFga7R48HcxQGKshUU/5pZTPqyahzUy9oR34y0sOoFLQ+edPDfbsfs2vX/i8pV5pnXrn7FW9GYGJcJmEGzaoSOiNUMX/MMwKxjPEyaKmzS97WfcYsZC87403Ir73Ow/oAAQtymDUfTIe831B1acR3c2a2ZkQwt6ifZynY167yotlFsb2O0GDPKoFJszKYlDNR2B+EsTo2KCnKVp8GH5iu0pzmWY8nF73AXKMQdo7x2S+sntE54It4x/Pv7werc1b9HOqXX6RAZxoHYrp1ZEUhpeLkOcn4R+hhowPzYEqVQcYMpD3rIWvFC2T8LUAILTYuWGHccoyV7+jNt2R4e5k327BrgcQKflMzzxBEEFjxAGOsMk6fW3NP7lXrYcG4BXv6+VaFT7tlYO7+a5c+51/itfOPaVoXTpuWGajsrjHSHAZhm/o839Vd3K0cVXolXMRNWgOKpXiGclh0S/AayOdyq5oKmWXdvUXaF2qd8dBQVZ3sbx0BR8ARcAQcAUdg8iPggsXk7yOvoSPgCOygCNQk24bMgT6AYIFg6pDxg5kY6pBAiBCQWBA1iBT8AIeQ4Ye2hb+B4LhBxs5ACB7IS36sQr5ZskjQnKpiBXWv9q4gXAbkF2IFBAHfQRhAvlhSZggHi/kPZhCnRmAPJiZwn0YUE6Ks3tZPtrvfSJCx7h5tRB13mGvUEX6qcR0LxvQfpC/knYkGfEY4Nnbe0p8WWi2eiBwH6T1s/DDXbTxb+DPmPOOaPBatwsBECMYWoaEgy1gDqCvvWVsg61hnEBdYY8hjkVyvTvz4wEK0WPtqiEFwTcLUyNiVTBineqFOztfnv5RBuCZEa/pK2+oVrstxCBwQiJC2EHqfrXt0GOwnIvYz4YzgTyJhNyhW/4pMR9I+S2hb7zTW1m/LCOXFfRB1aYd54QxWt0Z/Hg0Uy/2Zptx6kdqrlVhoYS6XLYqY7FHAsmf6FeaJfhUgszKK/qKcFaGUi/Z8IdMfBtmBMIi6s0H0TCEo9rb3rCju88DXg5kPXk64G9ZFhB4LBUi4q3aheqLyU5wWL1M+D9G5iBg59b68LrYo8lIJsoq6H4sK117tdXqCnBd3RXvPuOt7C3v3fM6s/gXPCvoXPuvO4ux9VhfWPkY4rsFIXXa2m9CGZwSeBXUJ8UHC+VAv5l8S7kzGGs518KCoVyD3yTjCDvafyyDzhyWcG92pdj3ylIRh0BSGmXblVW/X4FosF5iDRTozb3NhNlwrwUBoxzn1uxJqx7tWgqhVosUzIp4Zw4h3iAkQ4TzL8f5hHUrWNEJcCbcefYKIytrE8/9fZXgQcI+/Fq0CiFMZjY6yArAhi6l/W2Rv0agHV+Yac/PaFLOBKuFpoiCaiOuCD2MFzAgZhmcPwiV/G2AU2sncwAj9hNfF/6T4sb7zNwR/NyU4S5AYrJiYZiE8O3QgnmHIgMyqwTw5TEjmuuS0+LgMwYh7rll94r/0rD/ijdl1Ucv03nJ+t76e4h7qsIUK/zanr1jKS5iYkQkz81S5MJctrdMg6y3kw5ntLYU1ijG3plgsR1I1e6a1FwYkbHCvsosWg/ahf+EIOAKOgCPgCDgCkxABFywmYad4lRwBR2CnQ4AfkxAq1aEf+JEMSUfhhzekC+T8STLEC4gJfiAfLoN0pHA8BCoEIqQQa7wJHUaukmh7LOTtZOmUJNSJjB/1kKy01RKUG6GFkAFekKNgVxXUJNm9yPeWtHki2lUdhgLcjfjmPeQThZ2fSSgekcpJ37unxUR0xbiuaWPNwt3YLlx2MZvAOJFziWszTrnsekTuAAAgAElEQVQXJLqNpUSMSD9jHkC8sYt9AR4WxMRPv7MQWIBgAoCFl2L8MV8sjBrX2yxOjBI1rs24JjEt681HZeShqC1EwSdE1P2M97TeQ92K69K2B2WsfaxzEJAHyIgHv2lmqSUhK0Fr8NK4LzhNNPCv1LJFQgjPs9rCnKPtnbIr0msjWOAdQhu2R9gUsChqIehWg9fEUfw0oaD02XzSWlQqocZfpEhQmUyuIMo7UiaCMM4LwVWFbPHRXKk3nLGhM5oTr+1t61s20Prgr/fKlHpfq/OfJaNfyS0CGY3gA4G9j87tQKgwGSGSZJWEDDIqN0VNok9SMt0S6AaC3StPBNdnlmvL9m5HH1FpnvH8oG3uUY/+4x1XK4n2UIIA88WIYSOJ63TNoB8x/hHfEcIw1vY3pW2pPomxzTxgfF0vu1bGmNluMfwRK2ZMa84NDFTa5DYzrSmfmVMsV3ZXX04vNOWWDwyUd1GSdb5rywVxUzYXtiibRasS68yT70VOob1Wy8tmlYb5oxofzFdw2CqvCt4WEi0sHFenjoFwJwTRh+uiKkRzR2tRUM9gFY0MzZ15Wm3eqpXiRToH8RES/WYR9askWmyPeTGaMWLH2iYBC0FmGxlYQxC5qjcpmJDHZ9+W4cnFWEG4xHsVwWKo9d3ulQhPMsRaNpRwPuNUCG9VWGOqc41wnx/ImKe8Z7xuXHXKB4OejhMzGwvzMmvWdoelYn9hY29JAnTUKqFrVv9AZW6lHBeisDKzEodRLqehL68KndukiTg3n88OKCRUTl48Ci0WdCsRtzJyV+zvzLHg6uc4Ao6AI+AIOAKOgCOwzRFwwWKbQ+43dAQcAUdgCwTsRy8/WCGpMFub+dHLDj1IQIgKC6uCUMHuUQgFEo/yAxnC7XQZlBO7MvmhTbgWfrhD5FhCzYkkWLdV1ybkqkoS6iBtP94mEDp3yCAK2NULPhb7nhBZHTIIWgg0cJgoDwvb3Qn2GH1q5DOECP0L+U09jEAWZ5UIF0aSb8bShYxtNay2vE+6c5n+YrwxB+lXdq2bt9K2mEvcw8QJxoolDTcPKghgyEkM4Q4xjrUiEekYOxpX1QIa50OYMV9YNxA2bXyOqD2DeJKwyxsimZ3K/yUjJ0RtwbPj/2QfkbF+PZG2Z7jd77aWUV/IPUK6PKHe2AtklOFhk/yh1U5eAcsyc4OXK8H0YAWx4hIZpDY70sGtU9a9vZIxkzdExHa5kM9ph3SwrCKxQqSkeMZ4Ju9zmbhcKkcbykH8dFCOmpSMW+xx1J8pllfMCFbs2lLe2LXbyj8dMHfNnftMX/tgd6HU1R7EEYnGEXZY7+h/EGGX+ZYlRZ68HxWJFlmtVgqrtVURros1at6YmxF0R6XmX1Wapp2hgyCAWYN5HvFsGqxAsDPuEItZn+uWIZIls5YjvvCs43mISF/tOWCJtllXvyRDuGd8seYzP7ZrKeQzmZ5yWVJT0C4SeR+t8rupL3epDJR2q0TBNAkS/YpMOFMztllZSJZpzuakTjVlYwmQmeCxsrbUE0pK3zMPmKvVO/M3ty0dv8xD1oE/yG7RQLlRZ52lJw7h1BAd7NmZnKcE64lFzAJm70AwK+7VmImTsfNvsiSHlkQLhCDOH3Subquk3EN0JuOcMcAIZg0EB7yKGC8fpLl1zsVzhZBwt8jwuKLwOpxYwXFJGD7ZMenxzDmEQsYfwmq9wvpDAUvu8yfZr2SIFU/KuvBUuuOCDyYeNMueXhv29pUK8rxq0howQ7LUPlEgbVJhxCRu9VcqGj9xZfZAMS635HMkbF9ewlsrDGe3NOVXBYVcX6lSqWRL4RqNq9Xy5JqosIWDNNc/dgQcAUfAEXAEHAFHYOwIuGAxduz8TEfAEXAEGoGA7Xxmtx9EIiKDhTNit52Fg2C9hlaAhOcHOIQ3Xha7yCAf+SHKeRBDkAv8YIdY5Uc1n0NeDkcMNqI92+IakC62OxwSFBKLuPxgwiuFzxAuwHBPGbhSIPAgdS00VKPrawLUpj3fmwgNCDvoIIrFk6c/+Yz+t75KdlrLEs+LRlfMrzd6BEQCVkQAWhxzLgDJviny+7YpJnRZ6CkjvBgfjBO8iBApWT8Ye0q8LIVCpKfeJwl602radazWlpsDwplrJWGQhgoJNVxzU4GHtYaE2Yin75edUnMeO5DZyfx2GesXhXOCYQjPiITaOoxweBeoZTNFrB8u+vZfRLYfLF0mCWmUWRx0KLr7UAUvEDwrFBAnIQxp+8D2EiuqKhp39QwMTG9rWiuxIi9iWwl0Fas+jOc058L5+aiEeNHcUkbXjEuVXHPfzKgrP3vDQ4V5a+/aff76e45s6XpqTr7U3SqxYriu+uv3qe+ZdtevkaS9Tjktssr/QTiprUsYHCe6+9Z8fs1dmaC4MQqaWb8Yl4ghQwkW9C+CH3hDEI9IGNNx1WHYWLfJQfCyOjWz3E2Qvjz7SCAN+TtUgveRYzS+I8NVa3vz2UymJZfLzJE3xXwJF62aqZH6eUY2E8+UpLiyVIk3Ee1KtC2yeZ08K/Qsi2cLKYUTCgs6ryuOtac+TuYAOA6akyMdy4g4XYnXRUXPwEoiFD1H/YdnylYld5wWAB2hIGRJkWjBOvMp3Z/zmM94XNwto8+3m8eKVbxG3DIhgmcufw8wAUxII3/OF2SDbU5gjSKElgm/jNWhJhB/ezAuuR5/b+wnQ0zjvPfIanyUtoL6Gn1C+Dn6m1B818oQ1nq0/oFrUuSxFP/+nuVhuRxl+4uSJ7UeZDJhQblPcsVi3Kzx0aP9DS1KfiNxUl4VEjH7gvI0jSl9FK3LZbNdhUJ2YzaTnaGarta/K4V8JZRgsVWF/ANHwBFwBBwBR8ARcAQmKwIuWEzWnvF6OQKOwM6EgBGGkIYQBfyq5EcshB7xuCHfIQsgvztk7DiFmIe0gEDlRzqiBTsKIY4gL7mO7RRM4jBv4jGndDgoGxMQXvy4N0GGz02YYQe8hc7hPUQXuEGqgal5ViQ4p6CMlECz+w/1aoIFx3Bde85SVwgO+g7PCogP6oRYQX8bkWc7YDfHzh7JTf2YiUMgFS2i7UBqm5hZPY5oKIKbhYKCaGMXNASd5V4gzBhznTlhogVrDO8ZX+bJw7gzoZPPQpJAjwfJVLRAWMV74RMyvMRMRLRLIyng5QDBh8cEJCjtGFIESnMkFCvfUmz/tZr/LWp3GPw8Xh8sz8wOXlAvcfTmtgwEq6MVwbe1m/y+sEmhkSLNwaZEqNhWwtOQsKZeFvHGnoGu9ramcnupqzKjf8WssFzKKrzLrDgqzy7n2+L2TKU/07su7ts4UDpk6c9fNKP3yf1ylYGgqdId5Mu98ssYUXN4RvDMYM3ZlGQ8Cn4hsroSrwsGomXBaiXk/m7dCockD45/Gka9S4NsE8G48No45o6nNt4PyTpII/kcQpd74tGDaDRcYZyyNrJ241kBMYxXx2CFcFck//6tDOFiW+ch2apehIPSh0noNZHNczRWFyiqV7smWiRRYr08L8pKwN0q74m8nhQlOVDkJExks9lgQDvmZ4VSNpry2RmSqHoVJqxFJPVjlThCiACbrQj4QTxUenU0xPg69fHvdJ8unfkP9UDMaKZWCJykJ5ZywSQ9prBhR+gcQqslmx5kPEMRSTeT68N1ZKO+H6R9rGk8Yxkr5l0KNs+T4VVRryBocSxhw5akWOK9xXqwlVghodQ81Ow+rGd4sXLPE2V18axzY9Y6BCDWO3AEbe5bV3xas743UBinfP9AKau1fIZm52yNo3xFg0A+N9O1xOf1+QqNDcI/NSm/TVY5K/rjKBP1KcBck1QwhYKarnOaW5pyld4B+ev8Nbxgo7rFr+MIOAKOgCPgCDgCjsCEIeCCxYRB6xd2BBwBR2DECBiJCOnIj0rIAIv5zb8JMcAPZMIbsDv4+TJ2j0IKQvRBL7Bznx/WkIEQmogdkBsWMAUGc1xk5IhbM7EHGlFj3giEdgGrjhQLyFJ2CLOLkTBYkAMIPoQIASMEA7CxUEwTseXQBBP2qyJKIJpQqCf3p38Qoqgfx2KIGAhOEFyY7YhHU0lO3kH6L4Vi8r7UC3m0HcSKWoAsZJwJWcwD1gvWAcYRBBhksJGkiBZK9Bsy70m+bcSe5bfgOpxv1ui1geuzq/6PsnMH6W0SYjPuIe6eESFpO8fr1oV+0THMjYIkEObQYs2S/UWj7i2efqtwN3ZPEfAkFq7EG4O+sE/n9QQZiRdB4TPbVqyok7TX1rJNIX6uPaa1lG1u62lZ2NTXPHf3cr79sFKmaU4l37YgKPXv2p+feU9zWJrW1tV5eqbUN7O1vD4RKXJKepAs7SPzrEAsIJcI3md4fiF4I2A8LqqWdagiTIuyd2okEb4LUaNacDokjMuvXrDm47cvn/vvLVGmNRcHGYW/GTK6Hn3zFxnXZxybt1u9YWHkMEIFnnF4E75PRuLkeoVQiBfIGDPMAfOca/R4HuT2w36cyWYzQSYb9mUkJ4l5LmpC4iYzU84yFVWyS4JFG+lJtGO+X58VNF9bpVVoU3ymUChkppXKcVcxqsxuKmRv7y/GvRIuRvvMAu+y/hLg7wiSkPPsfFdtzUmyTl4L5gt+nRFSFnOHFSJOSHk2RXxUxtyDaOe6I1LIhkVpbAfYmsbfPHg5vDAdMyS5PqXmkpbzio9/LEN0YfwzfhJBrXhZgBfXVrDoA8t1wbObvCA80xfLCAF18jBVRxD5WVovvGPZeNIpG4mnXuJFJxELx6o5Ei/mZMJ4dj6XbctKi9ZEZaxsiAOJFPqbQROnWdMQgVjh5cJVypMS4G2h7xZu6Kk8VSpFxXmzlSpl+/bZ2Hraz3IEHAFHwBFwBByBnRIBFyx2ym73RjsCjsAkQ8B2PPNqO+wtNAE7RzFECSMZLacFO/wshBTvIeQ5hh/jiBVpwI9gRxErqrsNEgHiBBKFeNHsmITAgFSARIH8hyCAlID8QrjolCFmIGqYYDFRQ4H6WegMnrW8J3QJdWa3MLuNIS8QoQ6SESqHPmMMUD/qDYFr5FSmKsfFFnX2HBcT1YWT4rrMYcwINxOyGFO8Z5wz3xHkTBgjNAokHmKXNnNvJhUZgwicNhcQ9QidYyGv6pK8n7z89lBkmYFR9xh5CGwGK/Wy4JpcH9Kbc14/CJrf0eeIsJB6hHtirasOy2IeS8Tmx0OJub6HZvo5eiXs1J5JHos6FyepdCRUkjA3pWAXeWK8IF4Z/J/C3ZykWbaXyMmbUvxKqffGIFVs+McW6sheWbtowp75Sv8hM7uf6J/Wt2xtKdvSX8kU5mjP/VFhVN5LEYEOicIcu61RLyVWSHmRUpMRvHhWhPUFi2t0XURdyP+bZbbDm8+5P4QqYfOKGiUhn4SzJAiFSV8QCqhe4uC3zd54+cpKdvaSddNefXcxv/tDcai0G4OHemLdI3QhzydyBQwWtItrMHZ5BrJ+QghDwA4mVtAxtIMxnNLrg4dKangvjuKC2hVPJplCrIGn8FAVxe3pJcyPxIesuq8s1wrl4g611kdNOnIW7lGCM6/wP/NFOuMJuFq9PE+TuTfapEwNqRDVVM3WD8JlEQoN0Q+MCcu21e/ADH6J3EArC6nfo07VhOlfCs5WXQnL9S+ya2WIFtTFvKO2pUhE/VkPKIyrY2UdMnJI1CuMKwp1tTnAe565lNq6m3AGVmwW4bltmx8QYPGsGK7wdxr5KZhHCLeIFIxV1uxhw2o9smRNMHNac0aCVqTxo3vHRQlbfZFqquFE3edLp2yWZ84y1X5AHTFLlW4vRbH0sUy2WCwWtNeht6U1LwetSCJYqFBR8sPw4gg4Ao6AI+AIOAKOwBRBwAWLKdJRXk1HwBHYoRGwkFD8OIYaYG2GZjMPCX7cWiJJ2xloXhmQThBelmSSYyH8+DxJkrkDEtrgBUZ4TkCvQFZBuiEC8IMccYf3YMDuc8gyjmWXr2Fpu3yHItrGMuiMSKJ+1AOxxDxmEEsgPkxIgsgjcS1hVehfYmnTr4gUEHWQG7SLccB5XMeIDicextI7U/cc8ygyAp+5bWHQGOOdMkg5+5wxzxicJ9KKzxlTkFyMHwQx5sw6rQ1PaQdvMZ/LNTU1ZfKf+9Gd2swblLXDOyxHUUZEWVlihYkmI06OkHqkFCUyQHxfJCNvxX/L2KFcW16pD8hNcKXsszIIRfMyYv5AXjMHIAlfIoNkh8SGhN+6lINS+bYgH9tee1pPeJsBxfDfhAV1uEH2eRlz7EmJF6sbLVpUhZIBP/qNOQzJSh0QLVm3Wc8JeQQpaoTo0dlKf3sYlW5QfgO5yGT2ipOUJKHIbe2rzubxtpKbiDSsxPsKwUJds6VggecKbcSbAoKU5wPeEghfjBe+T547aneiRlWF3GFPPWIqSZffITub76tLGPXNbx64L9NauP1B1e3Q1v7buBcEdr2C8Mru/mfLWBMhzbcoujcNpK/ZHQ8+1JFd7H8zyDX5+E4Z45pnJWT8ZMhZUV3dxANAYkO7vCUiKU24VIRyuEBIzMsFqijxokvzj5wWjPeiNAx1bFgKK2EprkQt+jRUSJ/eMMj2q5Nb5c2i/MsRc3grz4Z6nmFVlUmETuHM3L82xY5k02fKlMEiCaG0qaRPMMJCZfFbUM0ifBI3hYiapju/Uf8iN8SvZZDx4P6ExntC/ms8TeSzidqxHjB3EGg7ZDw/ES9Pqmpv7VvmGbkseOZyDXBg3FTMe67Ku4J+oz/424K/G7gH6w7jc6iwZNX3/FF6D+7DXAJB7jdcjozqa4R9A+UkbCUKpV42SG9YrUh/M+VpwcBQZKh4vpYCFEzGmY6RBoYHjjJta3LP1lirtDblyq0zmmZlw2Cp8lpMZN8MAb9/5Qg4Ao6AI+AIOAKOwOgRcMFi9Jj5GY6AI+AINASBVEhI0ijogha6CTLCwrZANLEblR/nkDiEfLHd0BA6kE8mdlhIIerG+UYyNqSuk+giRvYb8QYRAQkA8Q8pRvgSSDHIE0QLsIV8gMAFS3CCOITAg5gz4acRTTTxg7pBPlIvyBzq05H+G48KCBbqilcFnhRGZuItQv1pE2QM/4ZQfVwGQcWx1J/+bbTQ0oj2+zXGgUC1l0Kdy5AQu1YwYEwwDhjHCFsUjiGoCwQ4RoGkgywzzx2OX078c3Z25/OZgijUPXr7SxIqFLImjnsqMbHQg4poL0v2HYwxvwXjHyEOQe7DMkjO6sJ6BgHJ36OvkiFKvCltD59B5jOXED7Y3Q0pieBAXP16paj8Fh+THa6rvowVMglp89f9zOYxwHW4JvH9WVfvFGHJ/NoUAKdOGSYpeJAKFKwnloeI9QbszbuKexMKrlNGWBk8q7g/x9E2PCDoM4j6UN4TrF9rN3lOqKuTTfeqGqJFGC7T5+slUrCWcS1wxWMEzMzTjhBJeN6wHrFuMAZ4zpRHQCqzfv4pPYfrP6cakkxclIfH0rmtfX85p5Sd/+CM7l+uEBl+sY7prZMHgDHEM8xEYvo8KTqH+lBfyGHC67AuI0QcKfun6nvWvMcrhzZfJ4MMrpsHgHOGIfKHuMW4v0pC+ohAXl8uV9qVznydNsvPDfPBUs2zJtHLyjkgkULhobRlvl1y1OpskOkVF51T5yvOV6ZXOSyW6JjVSra8Rpm7V3X3DJQGBspFcp6MpXYpOd8j3C3JNNgxzv4qWNRcOKtRGqr35KG0ydtig+boJrkEkQAPgt/L8B6gL7o0DxDBxlS/YdpkYwUvK6QUCs9Q1pWhCvOcfDrkruBchDXWlGqxgnlrCbURJg6QIU50yFif6iV7t3vS1k1h3TaJhIiznTLGPc9u1mb+FqCMRjCIlSRbThUhaFc0/TfIcWK6RMzdKlE4P5agrAo3aw1fIPGrUt70V0FZxxWle0X5bDhNeVBKStzdWyqVe5T2prxyTc9ow4lZG/3VEXAEHAFHwBFwBByBbY6ACxbbHHK/oSPgCDgCWyGQEBvJz81NhCNkEe8t3jDihP3QTXZiykyw4Mc0RBTnmXjBsRNBGEyWrqN9EAQY7YdcMC8KyD9+4CMSQJBBCEKG8UMd8hASD7KG78C8kTjZTmrb/YrIBKFofcTOcOoBoczucPqSfeDsQGbHOAQm9YZMoV4QJxyzj4xr2w7pZGdoanrxsjMgYIJBKlzYWmGeVIwrxgfjgjGF6GXEHHOCHeisK6wpRZFakKYrxX+3ilCdLreKXgkVzZpRMOPauqtYNZnQ1pR4jGIFZDGhnJhrCAHsxkaU+JgMUp5i8eGtC9lhT+JkCHbCRB2afnG1XtkNXt+rYtNBKzVLPhXOVMqAA4JLKo8ENysc1P8MEWW/Olku+TSI74+4wpwFz2qpIxYRWy9sjK1D4Mp5CJGQoohDEPHEymLdgRRGjMTDwnKOsC4xtyHzEScpx6evvNB2BEutD/FcIUm8/Q4JFqtFakMSc63fyfBIMUnGBCzqT39bMnZIZBN7q24x5FvO5dofkIFPlXeMQhtFvRItlrfkKqtyYTxAO2jPKvW3efkl4Q3viksLlB849f6JN0joWJ96VDBWaQPhfAjxhZDLuYSCev4QNYOgZg0HD/BJ8rqMRJhIE2Fvcemxju0RgGgbEcQtx21xJt4gcvlx5RaYJYcZOVuQtiLaSx4TOQkSvdlc5hklUO6WZ9PubGZQ9m1yE8RFkdYtLfm+XC7b1VTI9S+cx3AaXyHZvPqA8QDeJkwxv/ACNBFx800ykqzYVhGzqlApC14YJaR+6n+RiAesQes1V/DgikYjXAySVJs6MMfAkjHE/GI947PnDjNOOBcPHQQ35ibXQFjpM1EtFRl5xhJKksI9yJsCNngCvUHGvB2qkOydDQaMZwRC5j6h7ViHkw0mIxAIB7u+hkO8Wh46CB+EEGtXKwZkG5QThQzt68hrUSrFWeXiXqZQUO0aOyWNo9U6VnpX9pnevuLKrp7ieq3npX33nBPe8dTG4IhF00cjnAzTfP/aEXAEHAFHwBFwBByBiUHABYuJwdWv6gg4Ao7AaBEwMskISMiuNJhJEtIDigACmwJBYDuBLXyUkQ+bok2r7KBJmi1cAwQEO6PBxIgvPqMgCPAdAgEEBbsxOQ4iAgIBMoFjkj2JeLg0ECsjAizGNq/sGua+kJYQG/QdZAbiBAQRuy8RVkxwYkcmfQhRQr2pJ6SKhYSCDGI3ONfkHCcfBMKOXkS2WhPpc/OwMcGNMcKYIG46AoGFyUEMg+FEAOAcyHJtyA2kUUSrtHtXfhXhRrhIWVYklyZDMCDPir5KZZMIOl5C18hBEZKMW/IpXCZ7fzqmB+s25u95VV/WCyVVe+45auEK7ZOeJTrzUe0E/4tWBghtYs6zG3yo8h59CWF+oYz1gvmJKECh3hZ33khoW3NYp5nHkLV8h/iAcV/6guMg/Vm3CImE4ELbeI84Yx50iJSWg8TqidcYxv3xvuCarF1ci/ckK4dshmy1EDecmxD4MvO0s+uN9pVrsFYx8P5ZdoHMhITlmahnVSm3aFpT8TGtYeE7VS2Nl4g6gQn5S/Amy7X13TSrp+V4tSHqy0Ybl89b91VEKjBjjCLSEnYHj5lqsWawun41bR/rJWt78qyjVM2PeufSNxTbCW/zJqPzaGf1Glp3PR3GA2qw+iYeLTL6Z31TU7a1XIoOaS0U2hW9Z8ZAv/o2DHpELM9Vgu2sph8pzwkDpCTKYSmbDbtbwvzTTbnc8umt+Z6WQpaQUA1Z75mXmpOImiShRvgijNGb0n5gLmxRQj29crJYK0pF6MeMSsJEFYPzU39OuxYEPv3TI0EAobR/lIS99RWvPD9NTMA7iTHCnDlfNpR4Sd2ZM9QJQ0jZoDYnHgaqVxKuKzXec01CnyES8rcBAtxrajGo82+8gBjnzHnGPf2MaMHcH49Qwa1sDmstjjZK7Aor5SijJCgrNEqS0JbFcnlAf7sgMC/U0RpGGYX5C9oq5Yo8MjIDusBAS3NBwkZYmNbWVJgzo9XyjYygaX6II+AIOAKOgCPgCDgC2xcBFyy2L/5+d0fAEXAEknjkKnAV/Ajlx7MREqzR/Nt26psowfG2wx7iZXPYlvTchhAak7BrqkMuQXax35NXiw1PlSFtIRDYiQlJgdADYYFYAI6QHuxWtDAO4NtoLwuDzgg/BAn6lnAveIIQoqJDBnGHmEG4FfqQPqWe7MrulEEWsssTUYN6Mx4gNSFDEGO4JrGrE0+RHTBXieHor0KghjC1Ob55rot4ZfxAVht5DdlnO/0tfBzEOOOI8zYk8c43JT8wS7DWvbaKkd+ATuCazL1fyvBCIAwNY3u85Qe6AMQoIsNjojibwpYkiTRrA/OH+Y/gd+owN3qhvscoEO94Y1FHBMSfylgrIEnBimtC/uHdhZcAHlLMVwwqF48JQkAhOOJNAoHL/Ge3N21HrGD+0z/M/SSnSHpNPmP96pSx5v0hfU/7WD+4/wMyxCjEKY4ncfhE9JkunbSTcFOQswgz7Do/MBN1L8pGa2cW87sGpRzNif9V/wEnxteLZJ+WrZ3ZdeUBA4X90MT6CqUnu2Z0/wLxCHzoG8QbRJmRiBUQ63jAEHoIUpm2b1676wkKmhOJl0d6XPWz1Z4lzAN7z3FGlo/7GUrYJt0f7JK8RFIaZmzsintyOYXz6i8VRC53y9MiF5aCvaVBNCn8z0Amm10hzydlUg+nK4/MOrleLJXIsTrMBOvkktHV0pwvnXHkbg17XqWiBWIc6wPPR8REci7Qd8yZrQrhoXKyCk9Z1STWEzfWCFTotV20qvy9jHH/JRnX5Vm3VgIB7ylD4WpioHlUcDxzhWcf4j0iAjlVeEYOVRBnr5XhgcOzkr8TeouXBZHqYRsJGHdcB5GBDSAIZwgWhKDju6EKaw3jEHzoXwRhxDPzfCUfzmYhbZhrDfo1QnHqTQceXRojSyRUhJW4Mk1jZBf9mwzaivoU9Et43pDRYMnnFEhOoaKU30Ih/eLufDa3Qp45eNOt6u0tDUxrrcghxNkAACAASURBVMTuXTHWHvHzHAFHwBFwBBwBR2BbI+CCxbZG3O/nCDgCjsDgCPBj3sgIC1dkhDpkFD+O+dzyLlSHgNpRPSqq0TJyifZDNEBYQaCxAxPyD8KD5xokKMdCJPKKKABxCMFn4Zh4D4lisaUbOS6pB31jZAa7N81bAjIEctO8Q2gDdeMc6kP9IVKoH23iM76DUIHYhHCmTQgxvDePnCSTa/rdFm1xIaORXTt5r5USXLarnvWC8QBpb8Qj/7ZY/9UhxcbtRTEKVJgTEKKfkUE8E0aIzyC7hwu9Un0b2sX8gChEXEAIWZeGuunLnLtpd7IISjwSICw/JSM3AoLfW0dQX4QIhBUrnMdcJPcF8xUPh2+nX0JYYniBQPrikQAJzxrVIbMAOsxhyFcIVeYt3i4IH2DAvOea3AOBAq8DvmeXOIKECSGsBfRxdTi7cZPrtGOYkEokUGfnOPUFixdno66gtf8O+VX0y7rkoqMM0XERUcbyiyixeNipYfhANlq3WybqWzaz68ez86Vn3p7ixG1HUrjn12X037Uy8KwW6be4Rhr2CZzseWD41BvnkMJGkG/hfTFez6K0UuYNxRycLzJZaY+z2iEf4dC0sFmJKUqZqFWSoTwugorycW/M57MDypk80Nqcf1K76lcEmXhtPp/rntne1D9zekviIdDIkua16FP/Mv4Ymwhjn5ThafTSuvfS6pGhp/UkTnJbgJyeRgrBBurHSDr7TiqfvVMzkWsy53n2sv6Yp2CYO0GEOyP9r+EwebYzv/gUcQ8BEc9InuWcN5RYwfhgjF6he5fi3mBZ+WaN12LQK28rzmc+0h/MQQRB5ipjlY0NbBI4OW0rOJjHRG3zWTcJM4WQwjnMUbzGrG2NDtXI2OWafXq8d8sNbrUm2iNqhKLCqf7Kwi5BYp4ErbVRFGSU30TrRLw+n8su10DZWMhnupW/IlnzZ01vqXT14HThxRFwBBwBR8ARcAQcgamBgO0kmhq19Vo6Ao6AI7ADI7CJb06K7TQ00oUfrBAetgs6IcRFRDdsp+VUgDXFB2oE8gG6BKHiOBkEFkQHJCFkmu2q5oc6hOZbZIQgYQczO5MRKXhl1zPnKnwCv//HV6r6jwtRHwhV6gi5Qb2pD7tE2fWJqMIuY8g4wsNAxkCcQExC4EKm0J4/y9gBSox3hA92rNI+SCXaY8SdeXFstcvaBYvx9etUPLuKtKX6to4wJk3ISNaOBpGyI4KoKkZ9dX0gJQnDQvx8DLIQ2hMysDZEkt3nj3rz77IOGTuiCd3Efu/VIl+32tlclQwbshPyE2Ly72QWamZE9a9z0D1pfZm/1Bl8mev1CvPTQtbZ94RNIkkva8+1MuY1awLrAxixNiFc2tpB39Fvddeq4ZKCj7WRdp76zwQAEmJ/MA6yL+tuOzlY3/7yqGXg7szsjZdJuOg2UTk9LROsn3ZWsHrm28SwloJdV12gY+9Ve0b06ELMhYS+VMZazdjolIHlVhcwwSUVIOgL+42TrJFDhXRK5wuiUeINkWI8biGvRgyBBN9NnhVPKRdFTjvgdxfZ3NbSlF2gms4WcB2bFJMw8ZhRCJ8HJXCskFdFt4SLZTOnNffqs9JE7pBPk6CDAZ48eBchIr5EduKQ40cjMxJlH+GLxFNOf63E6XYAdTvB5X6u/16okburRvMGvd6b6UjEikpmrvAW8S7RpiSPkyZJd4RwQ9yjHq+oui9XtLCYtdX5tO7xkHCcG/cHv42eDDZGDwULJFowh5bIEBoloCXPfdqGtxV/R9Au1gXzuOS65m1SfQ8+e5+MNQmBgroxfztlSbi4UYa9GhLO6i/TMcTff2xymCNvCsTRg/TnYkHvWyRKLJKnXCiLsplMpPBPxaZCHk+eTjldLNFrn8bWM82F3OrXnLR3wwWvETfED3QEHAFHwBFwBBwBR2CUCLiHxSgB88MdAUfAEZgoBKqI5WRXHbkVqu5lJMq4ifWJqv82uq7tEockgMCHyIJw4Mc8u6zxXthXBhkB4UVYCEK7QE5C/nEsxJd5KhiJ2+jqQ4BYwltejShAoLDd0vBThIthhzWEJ7HuIWB5NrMblF2gp8lIBsx5iC4IHrQb0hYClJ2djBPEERO0dvYx0ui+nBLXq4nhX+ttwxipbEuBYgjQrG6MV7wfIBWZp1fKmKuMbxIvMw8QJjvSsc8Y/4UMYQ8hkjkMaYhwwFwPahP3QmKnRCLeFswhBALEPsK6mBDAevFiGa+jKQgtGGW4MDK1YoWFtCPeP2Hs+DfrEu2CkDeMknBFE0WGjqaxaQJ11jHw/mQQZi9W4uj3ZOKeZ2cUDygtW2yEUgQbCRXloFB6KigWOvDCEOaDLk+ITRCzrOP/T0b/sm4j5EA6g5FhU7fqqfDAmm470+t6ndWenHoncX873rwtxhVmKw0LFRJiTXVjnC9XPoJQiZCbtQteYzBuLWaD7mwYtvWXIyUvj2fp74Cl09ua1/T0FZeGQfyMPC7wnkPASJ4hJE2uVyRkjKY7tzo2nTv2DGGOEYKLufiXtD8GD9slxDOS2rAEQV0l0ixLknMXlRvnqeBseV8QcuneMBs8ES4Ibpdg0arQbc0SNHolZtyv2XiQZIA9dQxzsZ6YWK+BiPu36enaGa0IHotXBE9GTweLJFq0qQ4IoDxHr5DhVcF16WPyc9SKodbf4MJmgery2k0tStYqxhaiBy1jLI5rfFTfZIgcLNwbwYT5UJQwQQiohxVJdL4sVGioSBNrmoSJDRIsuvV9SR91K4vFmmIpWpkrh+uV96RLgsWIVMKatvs/HQFHwBFwBBwBR8AR2G4IuGCx3aD3GzsCjoAjMDQCNbv+G/bDeIrjnhB4VT/geQ+5aQQH4Z8gEyABISkI+QCxwGd4JyBYsEMRhm0ivQyNlbPcAYgN7L7mlb6kDpBBEJTUmc8hU/C8QFiBMIKg65AhwvBvCFXIFkSaq2SQtNXhTHjPc93ELb31srMgMExS4MkqYjEXYGCZrxByENaIjYR5QgTolF2Szg3EPUKwUCyEEnOGeRAPE9II4QLCrkvCBfHnEUgQBLk/14TUJFQU4V62RWHuI8DQL+yoZ52AfK1N1Dup+i0VLVg771L4p+Vt/bd8uZjvuDlXXv3sOMxtTWiLnS7mFwVlZWuOxE7HIVzwoE1ivUNMwquMtYw1EQ8LwnrxHWU4PMx7x4SH4Y6v7WvGgwkeWXIINELkS4UUnkOMccbhNOW0GIiicF25EpdaW/MrC0qY3DdQ2r+Qz3aKiF5RLFZIvt3TpjwzZZkEiW1JOIObCUSIiCQ7/2jaJ98bcoLQAwgYyPAYhW7XCJfXxSH67hANhTP1lLpLr8yDZ4TI4TqGvCcjLWWd/1uNhpnR2uBO5dNo0yrQKqFiV13rCH3O+sCzkhrwzOeZiDfmSMtP0r76lV4ZgxaSEbECz8aG/z023PqtMWR/S0QSJWL9fdindpajStwfB/Fu+iSOMlGPxIn1GludCilWyuYyG3t6i92FfK7yyJI1o50LI8XKj3MEHAFHwBFwBBwBR2BCEHDBYkJg9Ys6Ao6AI+AITBACkEmQHITXwIiPbWFT2KGMxwFkF2QkQgA7LDke8hORAGEDgxiFAJjIEAlGEEA0cR9EE+oAMUmdiHXPDnGElPNkhKvhuYxBjBDGgjYScgYCF/IFgtbIEhM6aCO4IGpYIt5BY7zrGC+OwDZHYBhBIdIObwvtBiFOcBnmLJ4Jlsya+QLpa2b5AUZFxKXeCn0SLrgH6wDrBUQ53hfMJeYnIsjfpiCxTkDD8sq8bUQhOTVzH48q1jDCQCUku+qVlIkO8TTWRqSiBfh0rm8/q2v1rPOnVTLtt3UsfeMf2/puQbRAWErykURhU1DOzkmEimy0Icl1MUghXwjEMB5krHVgg5CEt8WIBKlUFKAv0z3+w4ob9apiQgfjgnWYxNnj8kwywYPr6HqWe4T1uV2745+pRJV8r7IsKDzUukolzkbZeGUmE2h3fKVJgkXyjFIon20pVlTjQj0JSYi3BQIbXg4k5sbrALF9D6G8UbNjsPBtybWy9X2XyJFBYbyMrESa+/InUN6MpZGedBpeK6Ilwdp4bfB8fV5UXRApyGuFZ5bJJUPlvai+78/0Dzw8/iT7Yfqe75Fb8DJhPNYNRzayyo/7KAsJR5/0a2xskNil/NqhJlW4NA6ifLnCP4O18rRYpbFVysZBSXlPSstWdTVEeBt3C/wCjoAj4Ag4Ao6AI+AIjAIBFyxGAZYf6gg4Ao6AI7BdEUhyd8ggsCDmESUgqCBUIBoWyizkEiQDBAOEDz/0CVZBSAg+JwY1u7pNrDCvjXE1bpBcEeTC5v4wdexY5b6IFuwop67UH1EiiU+d1pd6sROXf7PLmO84hs84F4KHuOKQKBAzkGu2M522EO6Ge40oHMq4Gu0nOwKNQ4DxytjHmOOM9+q/U+t5Do1KrKiuaupxMZDmuCBZLyFfmJOQsrbWQKoyZ1lbWGOGK9TxalmHDNK+VuDAu4Pd29+REVOf+Y3HFPdt+K7t4So71u/TRM3xHU99qT8T9YYKC7UhEw18VyGffqRcFfQZuUmyEireFYdNJyo0VLe+XynRolOfE94JQQLBCFIZkpk1HNwulyEeIeLYeBhNH9uaNx6Cn36gDeat0ZDnQ9oeBAvEZZ5NiHHcq79UjvIynlWr9bzoXbGmW9GhgrJEi3gS7Iy3Z6558P1A9cQLBs8XnktnyF431rE00vMUVmqDbEaoGSXBYm9FIdtbfw3co9fThCLi/Wg8NGpvi0jx3rQ/eL4y/hDO7Flc6/k00mo37LhU+CJJvAlyiCc5eVuQaHt5mM3gmcakKfUXy736yyfJV9QID6GGNcIv5Ag4Ao6AI+AIOAKOwCgQcMFiFGD5oY6AI+AIOALbHQEjovjRDoECUcEPc0g/9nGeLoMIQ5hYJIP8IjQUxArPPI6DaOF7yEKI0ST+/QQW6mpkpMWrt3jpkJokN4XYRGSgfhR2KrOjlc+oJ+QEoTkID8VuVpKRQnhCtHJt2slOdEgL8+KoxmoCm+eXdgTGj0AdDwzmzVZJtMd/p7pX4F4IJOSRsXXhOr2HTH9BegbfIZRa2DYIZkLO8YoQgdBxoYz1BJERkZLPOB7xkWS/N6fzFC8O5i7tIyQUhOhULL1RpvWxKGietmTXbzx5wBPHsE6xJrNudXW1nfrhDdPOfL+8LGKFjbpb4sZNKS6sUYhAeM0QdgcMbQ2zneRjwaNRIi1EtYWGCvHeaADxW+35wXOA9ZpnGJhZId/AQJk01VU5ichvMEzIoLFgtcU5w3hAVVIPKMY2Xi/m3TdHsg5jmP4+UGx5m/6NyFc/3GJ1auvhapwG50qSeXcmKM1IqHkhp3wYFvjw0Bo/GrwsEfGHKuREIXE8BWGC8Irfl3EufyMwFhGUmKPUuFFjargWj+h7Ey44WOPCPHZi5UahvonQarlTRnRBP8gRcAQcAUfAEXAEHIFJioALFpO0Y7xajoAj4Ag4AlshYCIFO1Mh+BEdiCdtxCDkA1RGNVnyHP2bH/WEXIGEInY9JAQeCfzA5zmYwQ2iJmdIw+BPPS+4hYVpsvpZvgmIS0JAQY5aKBIIIYgT6s7uY8JGJUk3ZYS4gOgiJAcGDpbUl3sgdHAPz2fRsF70C+2oCKQhoiwUE3MNwdPEPryV7pYhOPAeQZB49oiFeAoQKoc1ByGjI33PXMQrgznKmgTBS+H7ahGG60HLThnPiuoxkCZ/pu6ikTMn9Rf2v2f53A8+tmD1x1inIOSDp3f5LGGh2KmeyZeXXa/k3CTsrg7HB1kPcW9kPqeNxqOiukp27njOt+vR/7St0XmOqslvew8Gdp9acrwRbanFaKz/NhGF8yH06WdCMHbKEPdmC7GyZJ43qDUfrnuT6tTWQ9RCuSiCWDORJ2YsOU+5L5InYWzSjskIW16DTwnpRmFu4eVTWwib+A0Z8/Yo2XdljE82ATBvmct4WiXeCUNUcZt/NUhSbvNCqh4/CBnUL6m/nTfRgtc2B8Rv6Ag4Ao6AI+AIOAI7PAIuWOzwXewNdAQcAUdgh0HAQnRYmAaILnbq4pXAbt1DZZD1EGLskkbI4Ec7YgXkIh4YxLfGw4JzIRKT0EkTJVbUQR5ShZ271JG6Yuzs7JAhUlBfPoMIgjwlZAp1hXxh1zahOJ4r4zqcR7spXJOwV+xShjwFI57xWQklgdo3nhAp6S38xRHY4RGoJmVpLDvKmX+WG4d5y2cIn3hGIHoy9yiIEyZA8Gr5FEyQgHblWERHI+l3BEDNC2bG8jkfDBYe/rHNGN7x1DSw+oOWtSN7W45aJg8LiGQSpJOzJExDSzUEgwZ4QFTXo1ZYaEgdqy5SO85qhZFJRZbXaXy12MKzBiEvoycO80H9rY0EleQZ9yY9qZri3mRuzA1n6DlXDorxumB1OC/YVZ8HykERhJILlJ89iDQ68KKgxAqShnCxWc4b3s/BwityuokVv9B75iqejAgsPFuZj3hZ8Pm9MuYlz03+FqgvhTS698dwveGSco/hkn6KI+AIOAKOgCPgCDgCkxoBFywmdfd45RwBR8ARcASqEDDKgp2Q7IiEKDlBxr5LCBOeaezsJRQUnhfspmTHZRJPPT0eYoIwLXum30NWNHoX7XCdZrs3qS9tYrcq1imDVEFgoe5Hy0i4DW2DcEG7aReCBNdAoHl+et6uekWguVZG6BoS2EL9QMJUNjmQhJOdBBsON//eEZgwBIYIyZTsYk6TYSM2WAg5Pq9eO/pSb42t6pjmyeBcSqNyIkwYFqO8MN5heJx0yCCBE8pZHhi0E5FVa5MU07BltQSKzd4kjRQrRlnfkR7O82WEPgHDX3IHJpzpU54z9DvPWZ49T2iUF0T/3xmXggHlnHgy7gpmZ0rBi+INeh51B8vC7uBkHXFUmA9WxiuDXaKeYF+FemrRlXqU9ams/83Y7Oc0PLzVR+DtgcB4a2oIi2xgwBORMYlIQX15nvL3QuL5ONjcHd2t/WhHwBFwBBwBR8ARcAQcgUYh4IJFo5D06zgCjoAj4AhMNAIW5ghPBIgwRAoTLiDyCd0C+YAYwU5ednoeJyN/BcQEnhWQjTNl7PjcnHR7OxD6kJ0IESTbxRAoIPsQWBAf8AQ5QAYRyGfUm/aSrPZKGSTROTLi42OEWmF3KPHD95Gx65mcF5CkFnLEBQuB4cURGAsCVYJG9Twa0ZyqIUNHdM5Y6rgtzzli0XRECW7JOsb6ZaRwukc+2WHP+suudnJ3ILROpWKC1A7RX+MFfpgcF2CUeBfJc4Znz0ZJPaFsmWTyfLir3sfBKoV4eixsD+brQZ7XE/l2iRe7ROuD5nitxk5/cIieYAUJHBFeGTrens/H6Ho8238t45m4vwyvyrfKyAvDcx1B/1uyv8gQJBCaEE/4u4B6EfbJMmjYhoEeFynGOyr8fEfAEXAEHAFHwBFwBCYOARcsJg5bv7Ij4Ag4Ao5A4xGAbICEIIcFRP61MkI9IVxgEBcQ9EaO4W1B2CiIDXZVsvOSHZcQLBBsCBnbJLFvmsvCECGnBW2B7IPYg1yBUCFWPqIDdeN7wlbhScF7xAeOIbwFbUR4gZiB2OE4SEPECrxI7HvOsVwYdm9/dQQcAUegUQiwfqFcsC5Xr6V4svEda/G9Eji2yTrbqEbpOjwjPJTeKAFNPWcSkUfiRU94ehDrNQmPljkjeb9RIaEyPPEU/umBZOT0SLQYCK7XO7wgELh4viPQ8yzDeGbjuUEoJ77neowrxhciRYcMUQPvRO7N95aHJPHMTAXHKZkvZpRd4Ic7Ao6AI+AIOAKOgCOwQyDggsUO0Y3eCEfAEXAEdhoE8LKApKDwCgkGwY8wgVcF/yZfxW0yiA08EtjxS/gHvDIgPHg1oQBSBHLfdnNuSyBt5y73RkyBZEFAgZhBsEBcIQEo9ePf7BylviQLpT08w/HK4Dy8LA6UkZAbceb+9HMwAYtVaWJxJ+C2ZQ/7vRyBHR8B1lLIY9Yk1icLmYVQzHesYUkS7ilY3LtiHJ1mYb/IWWKXScOC1QoH3QqbxnPa8lRxOM93no1fTT/nOYcRPpFxdanMwjyZB4XlBrHnufffOPrPT3UEHAFHwBFwBBwBR2B7IuCCxfZE3+/tCDgCjoAjMBoEjMwwrwILEbVUF0GcIFQSZP1JshfKzIMBTwzCSEGm4Y2BoIE3AsSaxZUfTT0acmzqcYGOAMkCAQO5Qr0gbnhFqECAYdcoCbXJb4F3xYkyPCo4vlNGeKuz07ZzHUJKIXr8Ma0oYaV43q/WvXo9l0VDus8v4gg4ApsQYJ1lFzy74hFerbCOsYbxamGiphpmCeHd4ITeUw2DbVXfWhHDPHLs1fLFWC4r/s34GnWItm3VIL+PI+AIOAKOgCPgCDgCjsDYEdjWiUbHXlM/0xFwBBwBR2CnRkBkO+03DwuIe8QH8554nt7/VkaS6tNltrP3Cb1PwlHISEoNiU/OCHZmQuLzHpKttL2JfPJopHUi1BMhoiAAqTuhrk6WnZG+fzL9nGAae6dtO0ivCDPsOgUD2oWAgyjDjlTOwUMj2em8vdtKHbw4Ao7AjoMASbYV9ilZpNOE24TnO0LG+nqdfbfjtNhb4gg4Ao6AI+AIOAKOgCPgCDgCE4WAe1hMFLJ+XUfAEXAEHIFGIwChT9gRwh6R6wEyfw8ZHgYIFIgWR8rwWIDw53gItKdllpQajwpyQvA94ZIIuzSZwiQRygKRAUHGPEMQJXhPolG+v062WHaq7Pi0/mBBOVjGexKTniZDpCDhLTjwzK/epZqe4i+OgCPgCIwPgRpBgvWV9YbcA89MBbHio5fcUg+AZL10D4vxjQ0/2xFwBBwBR8ARcAQcAUfAERgtAi5YjBYxP94RcAQcAUdgeyFgHgiEdsKzgiSbEPd4IJgA8Qe9h5zfU3aADC8EmChyPJD7AS8LPA4ekBHGhOtEk8TjgHrTRkQV4r4T5grhAQHiBhm5N94lQ6RAxCCvBYXvaQtCjnla8PmxMhKSIspwzbnp8X3y5iiqzZNJqEmr5i+OgCMwlRGQdwXVZz0mlA8i63o+k2gx1ZrlXuhTrce8vo6AI+AIOAKOgCPgCDgCOwwCLljsMF3pDXEEHAFHYKdAAIGBXbvkpOAZdowMUh8hAk8KEkzDjBECCW8EiPrjZIgcJPFEBCBBJ0mpOYe42SHhmCaRaEGd8LKA8EOIQHwhPBT5OQgXhYdIdcGDAjGDJLeWkJzvOR+sSEgOXnfJYBPxRplMba5pjv/TEXAEpjgCiKisuYiwU1UYTQRk966Y4iPRq+8IOAKOgCPgCDgCjoAjMCURcMFiSnabV9oRcAQcgZ0HgarcFex4ZecuYaE6ZBD4hIaCGIPkR6jAywAPBMImEQYKsYLP8cYgx8WBMhJaczweB5BpPZNErLBOrU4iSs4JdikjOrw0bW915+OJgScFBQEGQYa2gROeJCQlnS8Dq2tkiBiG41QlEqvb7+8dAUdg8iHA2sJ6hDhavZ5NvpqmNZIwUa9uU6LukxZUr5gj4Ag4Ao6AI+AIOAKOgCMwRgRcsBgjcH6aI+AIOAKOwLZBQGICN5JukSSlRpzglR28lpviML0nweufZRD0/PsQGcQ9CV8h7yGedpfhhYCg0SkjVBKfcy2OnSzFdiXTltVp/cnTgeDCd0tlR6eVtTgr5OPAc4Tk3DfJEGUQOZ6bYgAOu8rAD6+LDTI8UJyQmyy97vVwBHYMBCx0H2sqgoUXR8ARcAQcAUfAEXAEHAFHwBFwBEaFgAsWo4LLD3YEHAFHwBHYjghAhOFBAEmPQLFQBgGPBwH5HMjfwDF4XUDIPyJbkR7DZ8+WIVIUZHhpWLJu1JDtHhIqFWYM3kh1QmhBTEFYoD23ys5M201oLD4j5BVhoshxQbgnBIsTZE/JEGgIFQUOeJjwnnNs17OLFYa2vzoCjkAjEWBdQrBg7fLiCDgCjoAj4Ag4Ao6AI+AIOAKOwKgQcMFiVHD5wY6AI+AIOALbGQFIfLwkIN4Jc0RuB8QHiH2ECAreBoRSQtQgBwT5IPBWwMsAAYPvIPx5ReCoTLKQUAYxYVUI4URoFXJQUGdydFBvcHieDMEGTxPEB763QlvxxOAVbwtw4BhyXGCQiQOE25qkba9qir91BByBKYQA6wxCxWaxYgom3J5CcHtVHQFHwBFwBBwBR8ARcAQcgR0PARcsdrw+9RY5Ao6AI7BDIVCVwwKSHS8CBAkECAj9Ttlusj1khETC6wKB4nEZybhJSA1Bf6QMQp9k3JD3iByQ/jwHJ+su4OrQUHiW4EnxQNq2l6Rt4XPahXjzkAxPCo67Wsb5eJ6skyHoIOAg2FBoP54WCCJeHAFHwBFoNALuwdVoRP16joAj4Ag4Ao6AI+AIOAKOwE6CgAsWO0lHezMdAUfAEdgBELDcFXhV7CPDuwABA4HCcjSQdBshA0Ke4yHkCQNFGCkECsJA4aGAaGG5KyYzsWaJsWkHYgPtPFSG1wX/RmzZU3aA7Pey62XnyhBoEHBo670yQmJxLRJxcw5YeHEEHAFHoKEIpN4Uk3lNbWh7/WKOgCPgCDgCjoAj4Ag4Ao6AI9B4BFywaDymfkVHwBFwBByBiUMAEQKRYrkMweIJGcmk+YywSZD45GogrwUE/QtkiBN4ISBQWFgkjqeYIDBxNR7jlauSjSMwEBPe8m/wb0QahAnajMcJggQeFLQRcQNMSK59iewO2RkyQkRhYJhkMvfiCDgCjoAj4Ag4Ao6AI+AIOAKOgCPgCDgCjsBkQsAFi8nUG14XR8ARcAQcga0QqCLuLTY64gN5GWbJIOjxFiB/xWMyhAi8LPiOkEfHp6+ES4LcJ6wUYgakPseSbXuy7wZGVCEEFgXhgrBQ/PtgGcINIaBoK99Rficj6TbeFI+mbeYzRA6OI0SWFYSLyd7+qur6W0fAEXAEHAFHwBFwBBwBR8AResaxXgAAIABJREFUcAQcAUfAEdiREXDBYkfuXW+bI+AIOAI7HgIQ9XgYEPIJkYI8FRREirkyPCwg6vmefA6Q/RyPsIHnBZ4IFHI/QN5bLozJjJTlsuCVdiDYIET8IMVgb73uJbtPdpNsPxneJ7SR3BYIFOTuWJ3igWhD4XouVkzmnve6OQKOgCPgCDgCjoAj4Ag4Ao6AI+AIOAI7GQIuWOxkHe7NdQQcAUdgCiNgxD0iBGIDBDwCBR4WeEvgNUGOCiPkIfEh7BEqOAbhAs8MQkQhakD8TxXCnnoirpjIYF4mB6Vtw7uE0FCdsg2y56VtByM8MMh5wfm027wqoingXTKFh6tX3RHYcRFoa582fddFe3aUS6XSk52PPVIpl1lfvTgCjoAj4Ag4Ao6AI+AIOAKOgCMwbgRcsBg3hH4BR8ARcAQcgW2EgIkLeBlYeCMTMSDp+RzPChJsQ8ojXBA+6UQZIgW5HBA4CA2VEP9TgbCvColVHRoKyBEtECBIrL1OhiCxUMaznZBQtJNQWItSbPC4sETjnD9p83dso/Hkt3EEHIFRIiCdYsYHPvqZL73orFe8JpfLJ+Hlerq7Nn7/W1/94tc++/H/LEvBGOUl/XBHwBFwBBwBR8ARcAQcAUfAEXAEtkDABQsfEI6AI+AIOAJTDQGIdsQIwh7xys5eclbgUcFnrTJCICFi4FnxsAyBg3wPkPsQ+5Z4eqp4WNBHVldLmE2bSKLN550ycnMgSJBsGw8UsEC0QNSg7ZbjIvFAmQpiDfX04gg4ApMDAa0Z4WcuvOSKgw8/+tjPffTD/3rLn667urm1te20l5x9zlve8c8f2Gvx/ge+9/w3vHJy1NZr4Qg4Ao6AI+AIOAKOgCPgCDgCjoAj4Ag4Ao6AI+AITCACcRwHVZbR+xbZLNkc2SGy18rOlp0pe7ZsD9ls2T6yY2X7yWbI8rKcDHJ/ypSqtod6j4FBe9qmVr3Ol82U7SY7SnaCbH/ZPFlzaoX0XBM9pkz7vaKOgCOwfRF4welnveKOpzbGLzzzFa+urcnLX/emt/HdGS9/9eu3by397o6AI+AIOAKOgCPgCDgCjoAjMNURcMJiqveg198RcAQcgZ0EAQj7qsLzC+8JjOTbGIm3ESFIvk34I7wKetL3HEfYJHI6WC6IKe1lgPCQtpe2UabJAAmPE/DgPe3n3wbelAmFtZMMa2+mIzBlEPjMRd/78f4HH3b4mScchgi8lXfaN3981fXNcrk494yTjpoyjfKKOgKOgCPgCDgCjoAj4Ag4Ao7ApENgSu0unXToeYUcAUfAEXAEthcCkGWENiJeOrkcCI9E0mnCIRECifeERYLU599PyBAwNsdX3wFCIln+DgQJjBBYJNdGpKDNGGGgCKFlybqnRN6O7TWo/L6OgCMwOAIHP+vIYx598L576okVnPW7X1z5w/0OPPiwpuYWwtF5cQQcAUfAEXAEHAFHwBFwBBwBR2BMCHgOizHB5ic5Ao6AI+AITAIEbIcvhDyEPZ4TCBcQ9ngdIE6YMA9xv0OR9paMO20X4bJqdzybF2Xy+Q4g0EyCIedVcAR2XgRmzZ4zt6IyGAJXfv87X7/1zzdcO9Dfh4jsxRFwBBwBR8ARcAQcAUfAEXAEHIExIeCCxZhg85McAUfAEXAEtjUCKUFfe1t4ehMijEhDnECo4N8WNonzEk+DHZW4r9OuqZRQfFsPJ7+fI+AIjBKBjRvWr5s3f8HCwU6TTtH7yAP33j3Ky/rhjoAj4Ag4Ao6AI+AIOAKOgCPgCGyBgIeE8gHhCDgCjoAjMKURQMhIyfrq0EcmXljoqIqOiXZUsWJKd6BX3hFwBKYEAo899MB9iw84+NCMypSosFfSEXAEHAFHwBFwBBwBR8ARcASmJAL+g2NKdptX2hFwBBwBR6AWARMuECXqmSPmCDgCjoAjMHYEbr7xuqtbWlvbDj/6+BPGfhU/0xFwBBwBR8ARcAQcAUfAEXAEHIGhEXDBwkeII+AIOAKOgCPgCDgCjoAj4AgMicB1v/v1zzng+aef9QqHyhFwBBwBR8ARcAQcAUfAEXAEHAFHwBFwBBwBR8ARcAQcAUfAEXAEHIHthsAPf3/TPb/6832do63AXOW+mD133vzRnufHOwKOgCPgCDgCjoAj4Ag4Ao7AzodAdudrsrfYEXAEHAFHwBFwBBwBR8ARcARGi0D7tOkzTj3jZa+87aYb/rj06SdHJFwoRF942W9uuL25paX1lhuvv2a09/TjHQFHwBFwBBwBR8ARcAQcAUfAEXAEHAFHwBFwBBwBR8ARcAQcAUfAEdgCgTlz5+9yyxNrip/8ynd+MFJoDjvq2Gff8dTG+AUeSmqkkPlxjoAj4Ag4Ao6AI+AIOAKOgCPgCDgCjoAj4Ag4Ao6AI+AIOAKOgCMwHAIf//K3LkO0IMzTcMfy/fn/9IGPIFjMmjN33kiO92McAUfAEXAEHAFHwBFwBBwBR2DnRsCTbu/c/e+tdwQcAUfAEXAEHAFHwBFwBEaMwA+/+42v5HL5/Mtf96a3jeSkxfsfeAjho9atWb1quOPbFHNquGPqfZ/N5XKEnhrLuX6OI+AIOAKOgCPgCDgCjoAj4Ag4Ao6AI+AIOAKOgCPgCDgCjoAj4AhMUQSuvPa2B3990/1LMiq1TUA4+Nf/+MTn/+/iH//6c9/4/k+uvbtz9R/ueGzFp7928Y8wPDTe/I73vL/2vJee87o33vz46gETLWbMnDX7/f/1qf/9/q+vv/3z37z8Z3tJ+ag9Z/H+Bx3y5e/95Kpbn1hbuvaeJWueffLzX1h9DHX578997TuHHH7UsUNB3dbePq0R53GNTDabff9/f/qLJ5/64pdWX5OQWJ++8JIrXveWv3vXSLr9jJe/+vXf/dnVN93wwNKNJDrnmic+/4VnjORcP8YRcAQcAUfAEXAEHAFHwBGYygi4h8VU7j2vuyPgCDgCjoAj4Ag4Ao6AI7CNEfjxpd++aMFuu+9xwvNOO7321iTXPvCww4+KVRAMZsyaPae3t6d74e577LnHXvvsu9c++x0wZ94uC2rPO/iwI4/OylUiiiqVRR17L77sqj/d+Zrzzv+H5pbWVsj/5552+pnV5xz97JNOufjn1/ylY+9997/0m1/5Qn9fb++/fezzX6k+BqECIWQoeD76hYsuvvDyX17diPO4xqFHHH3ca1Xvag+UV7/xb9+BWIFo8b7//OQXTnvpy181WJ0QPP7nf79+CbZh3do1X/z4f3zwhmuu+hXXfO5pZ5y1jbvab+cIOAKOgCPgCDgCjoAj4Ag4Ao6AI+AIOAKOgCPgCDgCjoAj4AhMXgRmzp4zF6+Gz1z0vR8PVcsjjnn2ieSvqPU2qHfO5RIovvOT39+IZwUeBdfc9cSqY0947vM5FtGjOuTTrrvv0fHHe59c+4Pf3ngXx3PMa9/89n/kXtP1gV3/rf/43n/Dw6OeJwjHIBxwzkc++cWLqus01vO4xhv+9p3v4Zp/c/4//gv/PvhZRx4DVp/9+qVXnn72q869/ckNEWLEYLghaHAMIocdgzjDNV/8snNeN3lHhdfMEXAEHAFHwBFwBBwBR8ARcAQcAUfAEXAEHAFHwBFwBBwBR8ARaBACTXKPeMd7P/RfHYv3O2C4SxKK6S+PreqfJoVgsGPPfevfvxuivZ5HRfU5JOSGpH/7ez54wae++t0fEt5pn/0OPHiw63LvPz24rGu3RXvuZccQZop7VYd34rgvffeKX9W7Dp4MhLbinNqQUWM9j/vgscE1d99zr324x2W/ueGOS391/W35fKHA97/8871PXHj5L7bw6LD6IdCAwzvf9+8fra7zP7zvI/9zW+e6slJ8zBiuX/x7R8ARcAQcAUfAEXAEHAFHYKoj4CGhpnoPev0dAUfAEXAEHAFHwBFwBByBcSJQKDQ1/e+3Lv/5uW99x7sz4da5KWov/7tfXPlDzhkqr8Ihhx997LKnn1qyZtWK5UNV78jjTjgZD4qmpqbmU19y9jkfetfb3vDYww/cV++c40963mnkqrjoC5/472eeWvKEHbP/IYcdQXLvnu7uLj7Dq+KwI485/oF777y93nVOl7dCxz777v/w/ffcde+dt91sx4z1PDv/ANVjyeOPPvz0kicee4USk5Nn44J//rvzSqVikWOUHzxfrz6KfNV2waf/7xuPPnT/vRd+7hP/VX3Mc0457cUP3HvX7d1dGzeMs5v9dEfAEXAEHAFHwBFwBBwBR2DSI+CCxaTvIq+gI+AIOAKOgCPgCDgCjoAjMLEIQJYfcsQxx739tWee+vgjD94/3N3+/Mc/XMUxx554ygsGO/bI455z8l23/eXG4a5F3gelrqiQb+IXP/r+d/90ze9+Pdg5b/y7d793/do1q7//ra990Y7BI+TU01/2yl/86NLv2md773vAQSTwfuSB++6uvZZSZeTO/6cPfITPf/2TH15a/f1Yz+MahabmZnJ03HLjddcg5ii01Icu+/aFX3rkwfvu4Xu8LOYqfwe5KWrr9Ipzz/tbQl399/vfdb6JGxwzZ+78XRBB7rj5zzcMh6N/7wg4Ao6AI+AIOAKOgCPgCDgCjoAj4Ag4Ao6AI+AIOAKOgCPgCExpBCyXw4vOOue1o2kIuSYIeVTvHMh3QiNV52IY7NqEYOLYvzy6sm+XhbvtPthx8xfsutttS9ZX3vWB//iYHUNYKMIsXXH1zffhpWCfn/Wq15/HNfdavP+BtddDHOA7rDb01FjP4x4HHXbE0VzzzFed+6Zz3vCWt19331PrqnNqUBe+r64/5+Fd8rPr73zkG1f85rraunItziFh92j6xo91BBwBR8ARcAQcAUfAEXAEpioC7mExVXvO6+0IOAKOgCPgCDgCjoAj4Ag0AIG3v+cDFxCC6aqf/eiy0VwOT4w99lq8b71zDj/m+BP4/I6bb7x+uGvKGeJQjvm5vCtWLHvm6cGOP+6kU04lZNMvf3z5JXhJvPL1bz7/8t/eeCfHv+P1L39RX29vj527z/4HHoynwpOdjz1SfT1FZMq/7R//9UN8pghL62u9ScZ6Htfb/+DDDuf1gbvvvO31b3vne779lc9/UrdYV10n3j/+6EMPVNeJsFqLOvZefOnXv/z52raf8LzTTuezO28d3lNlOJz9e0fAEXAEHAFHwBFwBBwBR2AqIOCCxVToJa+jI+AIOAKOgCPgCDgCjoAjMAEIkGMBL4OfXnbxN0d7+dXKTYFXAyJA7bmHHnns8eRcICfDUNedMXPW7LnzFyzkmMsVPmmoY8l1sWb1yhWESPrpdXc8/OGPf+FrN177+6te9+ITj6wVOmjT051PPFYpl8vV1zzr1a8/b/bcufNXr1y+jNwVsUr192M9j2vsd+Ahhw309/WRcJt2Xfatr24OW8X3hJvi9eH7772r+p4vftmrXkeYq2t++8ufVn8Ors8++QUvJFfHcHlARtt3frwj4Ag4Ao6AI+AIOAKOgCMwWRFwwWKy9ozXyxFwBBwBR8ARcAQcAUfAEZhgBA45/KhjucV9d99x62hv1dzS0holpVKpPZeE13ffdvOfawWB2uMWH3Bw4l3xwD133ma5Hgarx+FHH38COR0++oWLLkageNurzjjlfX//pldXezHYuYSKqvWuIIcE3hU/uuRbX5sxa/ace26/+abae431PK6z30GHPOvxRx66/7Xnnf8PF1/0pc/29vR0V19f6S0Sr48nHvmrhwXhoE445dQXX/eH3/yCPB7Vx5/wvFNfTEipu9y7YrRD0493BBwBR8ARcAQcAUfAEZjCCLhgMYU7z6vuCDgCjoAj4Ag4Ao6AI+AIjAeBWXPnzef8tfJcGO119ujYZ/GqFcuWIllUn0vyacj7e++89ebhrrn/wYcmYZSu+tkVlw93LPkt7rvr9lv+5sznHffWV7745NtuuuGPg50zT/kupGk8Wf39K9/w5rcjVFx/9VW/RLy4+/ZbthIsxnoe90F8kVNE4cDDjjjqB9+58P9q60a4qcceeuC+6qTae+y1z77U6bY/b92WF575ytcg+NQTVobDyr93BBwBR8ARcAQcAUfAEXAEpioCLlhM1Z7zejsCjoAj4Ag4Ao6AI+AIOALjRKBfiR+4xOw5m4SLkZbZEjoUAulZeFHUnrP3vvsfSDij+5XLYbjrHXDws47gmKt/8/Mrhzq2UGhqIvzULTdedw2hnIY6tkmuH23t7dPWrFyx3I5ra582/fx3v//fL/3ml7+wYOFui/j8qc7HH62+zljP4xokBMcbYl+JFj+6+Btf7enu7qq+Nnjsuffi/R68967b/397dwGeVf3/f/ynYBDqV0VAQjoGbGOjRzdSSiitghKKIAIiIClIS3d3t3R3b2OMMWCw0ThihHTo/7zA4/9wuLfdKxzy3HVxwe7zycc5t9fl530+n7f1c3OHSdDhgwesn6dMlSatweupHRiOAiuRuXIdAQQQQAABBBBAAIHnVYCAxfN65xg3AggggAACCCCAAAIxFDCPJzKTOzvbnI49UuJrJcC21zECFo9yNdgTWjtqW/koFDiwBw/sZd80ckLos/v37t6NbIyJkyRJqjK3bt3450imJq1+7PznX3/+OXnk4H4Zsz7OJWFsDnkiwXd066mtzH8nDn/w4P79WZPGPJG7Qte1k0JBC3tOj1TGGVSOxtKifbfe586cOnHv7p079pwXkc2f6wgggAACCCCAAAIIPM8CBCye57vH2BFAAAEEEEAAAQQQiIHAnh1bNigfRO2GzVqkz5w1uzNNZcvplvvzr1u1C/T389lq5F6w10mVJl16fWZNFJ09l7uHdkhYy+pYpgzGbgztmois31s3/3i0Y0G7ICIr+5pxJJXKGGv9t/W3+q735Tethvfp3vGmkQlceSquXb0SpgTZ1raiW09tKHm5/t64atliJfS2j1HHQemz4KOHD1mvJU76xhv63Yhz3Dc/d8uTv5CO1LptJMHQLhUFQXTt5QQJEkQ2d64jgAACCCCAAAIIIPC8CxCweN7vIONHAAEEEEAAAQQQQCCaAkr0/PMP3371+uuvJxo/b8WmfF7FSkbUVE53z3wjpy9a/fDBwwfdf2j+pT1/hepq54X+TpQ46aOdDpWq16o/c8UW7zwFixS3tq1ghXYdKOF2ZMNXAmsFAswjlMzyOvqpYfPW7b8wAijmZ1roN/9tnNL0Tt+Rk+ccDTzot2Tu9En6/A3j7KYLRpDG3md066kdMyCxaNaU8Y7mooTb+tyYwlnr9WtXw8L0e6q0j4M876V4P1Wf4ZNmDerZ6QcFLvy8d+9Qjgvdm36jpsyNzInrCCCAAAIIIIAAAgg87wKP/meCHwQQQAABBBBAAAEEEHgxBXZsXr+6ZcNPq/QcPHbq2DnLNmjHw/oVSxcEHtzvE3bp4gUj/pAwTboMmcpU+rhmlRp1Prtj7Fxo3/yL2kcCDux3JHYyOOioPm/btffAyxcvhNZp2LTFtg1rVmzfuHaltbx2Eeh3v327dzgjv3LJ/FnaKaEAhfr2yF+oSM16jZoqd0R3I+hitnHd2D6hHRSffvbVN581bdlWQYDWX9WtpgTWKvPSyy+/bKSYuG7vM7r11E6GzNlcToUcD9q1deNaR3PJlPXxDourYZcvWa8bybY3aVw/dO87ZP2KJQsaNG7ReuPqZYuNnRgByovxhzGoqUvW7zSG/HL/bu1bOeNEGQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEnmsB7Txo1rpDtxU7A074nr7+l/3PrqDQW3rLX0cqRTRR7ZqYvGjtdtX3OXXtzz4jJs4yTnJKbK/zfaee/Rdt8j6sxNLOwCnR92/b/I6Z4/I+ceXBoAmzFru4unva67fs0L2Pym09dOaqV/HS5a3Xfxk6fvq+kLD7OtoqturNWL55b/GyFauGN49JC9dsW7PvyBO7K8yyjVu26yQnjbfnkHHTdPRTiXKVPtLvmmOfkZNmK2m4M0aUQQABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEDgPyWgoETR0uUrVapRu0HZytU+8chXqIiZlNrZiSrAoCObwiuft1DREmbuB2fbVN4L1StUrFQ5tR9ePe1IUEDC0UK/5jJw/MxF7yZLnsJeP7r1Ihu/jnVK8X7qNOGV0y6QLC653HRdO0bGzFq6zvvk1Yc16zdqGlnbXEcAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEYlUgV+48+ZfvPBii3RULN+x9IkF3rHZEYwgggAACCCCAAAIIxFMBkm7H0xvDsBBAAAEEEEAAAQQQQODFEajTqFnLiQtXb/Xds3PbyeBjRw85kYz8xdFhpggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIBCnAjo2q//oqfOUr6J+4+bfv/rqa6/tDbl8r+6XX38Xpx3TOAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCAggQ8yZMqyaOO+wI1+IRfzeRUrqc9cXHPn0ZFQufMVLIwSAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIBCnAhkyZ3NZ5xN0/rftB46nSZchk9lZ7YZNW2i3xeuJEiWO0wHQOAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCLzYAokSJ06ydOv+oHW+x35PnTZdBqtGv1FT5s5audXnxRZi9ggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIBDnAs1ad+imY5+Kl61Y1drZywkSJNh88FRY+54Dhsf5IOgAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEXmwBHQOl3BV2hfyFi5d6HMj4sMqLLcTsEUAAAQQQQAABBF5UgZdf1IkzbwQQQAABBBBAAAEEEEDgWQskTPjKKzoGKuhwgL+972p1Pv/q9q1bN3dt3bTuWY+L/hBAAAEEEEAAAQQQiA8CBCziw11gDAgggAACCCCAAAIIIPBCCDx8+ODBvbt37rz51v/etk7YxdXds1zlap8uXzh7+t07t2+/EBhMEgEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBP49gQFjps3fE3zprmeBwsVeT5QosVfx0uXX7DtydldQ6K006TJk+vdGRs8IIIAAAggggAACCCCAAAIIIIAAAggggAACCCDwwgikeD91mmU7/IOVr8L8433y6sOqn9T74oVBYKIIIIAAAggggAACCDgQeAkVBBBAAAEEEEAAAQQQQACBZyuQ9I0331LOChfX3J7XroRdXjpv+uRAfz+fZzsKekMAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQQAABBKIh8Nbb77wbjWrPpErKVGnSxkZHr72eKFH6zFmzx0Zb0W3jrf+9/U4Wl1xu6TNlyfaS8RPddqiHAAIIIIAAAggggAACCCCAAAIIIIAAAggggMB/TiCnu2c+39PX/ypetmLV+DY5zwKFi2ls+byKlYzp2PqMmDhrwoJVW2LaTlTrv5wgQYJqdT7/atbKrT4+p679qfnoz4zlm/cqiBLV9p5l+Wm/bdz9zQ+dejzLPukLAQQQQACBuBB4OS4apU0EEEAAAQQQQAABBBBAAAEEEIhdAVePvAXU4v17d+/Gbssxb61EucdBFAUuYtJartx58pevWrP2nVu3bsaknajWTZk6zQdTl6zf2bnv0LGh58+e7vFjyyatv6pb7VTI8aAcbh55s+dy84hqm8+q/JvGdhC5sRPkWYnTDwIIIIBAXAokjMvGaRsBBBBAAAEEEEAAAQQQQAABBGJHQEcUqaUAP5+9sdNi7LXikd+rqFpzy5O/UExa/bZdl19U/8Yf16/HpJ2o1E3zQfqM2tHxl/HTsHq5In77du8w62fIks2l+Q+de549dTIkKm0+y7LZcrrlVn/HjwQGPMt+6QsBBBBAAIG4EGCHRVyo0iYCCCCAAAIIIIAAAggggEC8E0iSNOkbtRs2bZEgYcJ/Xt57N1nyFOkyZs4a7wbrYEBZc7i6nz19MuTa1Sth8Wm8xmlJic0dCDF50z9voaIlChQtWUZzu3Xzxh/PYo56JoZOnrfsz4d/Pvzi47Je1mCF+s+dt2DhjauXLb504ffzz2I80ekjW07XxwGLo4cJWEQHkDoIIIAAAggggAACCCCAAAIIIIAAAggggMCzFihbudonyknQpFX7LupbOQsWbNgT0H3gqEnPeixR7U9j3RUUeqvvyMlzolo3rsvnL1y8lFyX7fAP1t8ZMmdziU6fUxav22HmjWjTpffA6LQR1Tpd+g0bt/vYhdvmLgVrfRfX3HlknjZ9xsxRbfdZlu8xaMyUfSFh91955dVXn2W/9IUAAggggEBcCLDDIi5UaRMBBBBAAAEEEEAAAQQQQCDeCWxavXzJmZMhxxs1/7598pSpUn9cq0EjLa7PnjR6WLwbrG1AGY1xKvHzoQO+++LbWD0LeD3KW7Fg+sQx+tvNM1/BqI7Rq0SZCjpO6vBBP1/VvXlGJu8VAAAgAElEQVQj7o+EUn9Ksj16UJ/uRwIO7LeO+dVXX3ut24ARE8YY106fCD4W1fk8y/IubrnznAgOOnL//r17z7Jf+kIAAQQQQCAuBAhYxIUqbSKAAAIIIIAAAggggAACCMQ7AS3ojh3St4cW/tt17ztE+RKWzpsx+VRI8DHlMYh3A7YMKLuru6d+jY8BC498hYrcuX371tK5MyZrjNHJY9Gsdcdufxo/c6aMG6E2bt6I+yOhWv3Uo9/J4GNHp44ZOsB+73/qM3j01bDLl6aMHtI/Pj8XOo4rQ6as2Y8eOugXn8fJ2BBAAAEEEHBWgKTbzkpRDgEEEEAAAQQQQAABBBBA4LkW0LFK166EXb537+7d0hU/qqHJVK5eu8FHn9ZvqMXyCvld0l4MPX8uPk4yh6tHHiWFNgIW3vFpfAkTvvKKW54ChQ75+3pfvnQhVDtYlMciKmMsXLLsh64eeQusXbZoXui5M6cfByz+iNOk254FChdToKV980Z1Hj548MA63sYt23UqUKREmboVi+XRcxGVuTzrsjrKSs+1uTPlWfdPfwgggAACCMS2AAGL2BalPQQQQAABBBBAAAEEEEAAgXgnUKhYqXI/dOs7OEOWbC737t65owFqoVpv1/9+7uxpf9+9u+NrsEJjVT4F7QaI64X8qN44F2Pnh97y9/fZu0t1Dxh/l69SvZZ2sdw1tl040552VygYM25Ivx5mvoi43mFR76tvWim4snbZwrnWMdas36jply3adGxUo0KxsEsXLzgz/n+zTE53z3zq3whY+Pyb46BvBBBAAAEEYkuAI6FiS5J2EEAAAQQQQAABBBBAAAEE4qWA8hEMnTJv2SkjF8FnVUsVPGP849bNmzcSJEyYUG/Qz506bmSg//5Y37mQp2CR4jncPPLGFEVv0GfP5e4R4OezN6ZtxXZ97VRQmwe89+zU3wr8yFWBDGf6KlKqXEXtyNiw6rdFQYcD/BMlTpxE9e7cvnnTmfrRKZPi/dRpSpStWHXOlLEjrDsoKlb7tF67n/sN/fGbhrXj49FbjuYaX3feROe+UAcBBBBAAAEEEEAAAQQQQAABBBBAAAEEEHghBMyFcB33szfk8r2sOVzdZyzfvNfn1LU/q35S74vYRvi49mdf+p6+/tdGv5CLMW07c7YcudRW7YZNW0SnrWTJU77/TrL3kkenbmR1Bk+cs1RjUx8qq+CDftcOhsjq6vq03zbu1j3Ikj2nq36vUa9hE9XPX7h4KWfqR6dM0+87dN0TfOnum2/9722zvo4F03MRm89CXLqb416wYU/A4s0+R6Lj8G/X0c6cDzJkyvJvj4P+EUAAAQQQQAABBBBAAAEEEEAAAQQQQACBZy7whrFCvfvYhdtKtqzOU6ZKk3at99Fz3ieuPDCPIoqtQTX6tk0HLbxPXLh6a0zb1GK62nL1zFcwqm29ZPws3bo/6Ju2P/0c1bqRlVfbmw+eClu2wz/YLKucFjLuPXzizMjqa3eF5tVv1JR/jmVSoOPRXI2cFpHVj871l42fFTsDTgwYO32BWb9Jq/Zd9oWE3a9UvVb96LTpqE5cupv9acHf++TVh78MHT89tsb9LNvp2n/4+AkLVm15ln3SFwIIIIAAAggggAACCCCAAAIIIIAAAgggEC8EtFhdtnK1T1555dVXzQEpaXGHX34dkThJkqSxOUgtWGfK6pLT2ld02+/Ya+BILai/+trrr0e1Dbc8+QspAFD6w6rVo1o3svLaFaG2ew4ZN81advKitdsVJImsvnZXaME9Y5bsOcyyX7Zo21FtaldJZPWjc71A0ZJl1H7J8pU/fjdZ8hSDJ85esi3w7DWvEmUqRKe98OrEpbvZpwJYMdl5E5vzjWpbOqZN7j/+3H9oVOtSHgEEEEDgvy1ADov/9v1ldggggAACCCCAAAIIIIAAAn8LKF/B2mWL5t2/f++eiXIk4MD+3j+1aa6cFrEJpSTSx48GBlj7im77Od3z5DOaOmAmC49KOwWLliqr8j57dsR4p4e93zwFCxfXZ/v37dpuvXbAZ89O7VgxTlx6J7yxFi5Z9kMdH7VqyfxZwUGHD5nlXnvttUdBmdvGDYnKPJ0tW6VGnc+uXb0SpoDSgo17DxU3cllcvnghNG26jJliI7hkjiMu3c0+sud099C/D/ru2+3s/ONLuVzGDpokSd94My6ey/gyR8aBAAIIIBA9AQIW0XOjFgIIIIAAAggggAACCCCAAAIOBbTwHZXjmyLaOaE30bPmyOUesH/fnuhwZ87mkuuckWX8yuVLMc6lYe/fI79XUX3mt/fJgIXf3wm4c7p75gtvzMoj8fDBgwejB/bqZi3zmnHOkX6/c/v2rejMN6I6ci5h7KxYt3zxfAVLQoKOBG7bsGbF1bDLl9r3HDB8ypL1O//3zrvJImpD17V7ImXqNB9EVC4u3c1+s+dy87h37+7dIwH++6Ni5ewcotKmvawCQkq+Hl4b5g6ag0481wpsRHcsOqIsunWphwACCCCAAAIIIIAAAggggAACCCCAAAIIxAuBlxMkSPBjjwHDipWpUNk6IB2tpPwHdRo1axneQBs0/ra1jurRcVPhldFi7lctfvhpnU/QeZWdtXKrj6PFcuVy0HVrMmgdZdSsdYduygFQtHT5StY+tFD8Q7e+g0dMW7hy0IRZizcdOHFpve/x0AFjps3Xnz4jJ81u+M33P8YGsvJ/bAk4fUV9Wtt7L8X7qTRmJTh31I92V+h6l37DxtmvK3Cga1E5okv3aMikub8NmzJ/uZm821G/xct+WEVtOzr+SW3oeKpfx81YGJ5Nw+at2+toLrWhP3oOlEdC5WPL/e13k72nHCsT5q/c/HWbjt0juk9KGq9jtVTm3fdSpNTRYcqZ8m27Lr+Et1skojmE11fFap/Wm7p0w65tgeeuK/+HvhfKP+KovHbV6L5uP3z+j93HL97RM26W+7hWg0Yjpi9apUTtizZ5H1aydfO5VB4T3Xv7fVdSbrWjZ0bt6Hv5WdOWbacawSXNVTtk7ONQGc1zzb4jZ3VPB46fucjukc+rWMmfeg8eHZGvxmJ/tmPje0MbCCCAAAIRC4Qb7QYOAQQQQAABBBBAAAEEEEAAgRdVQIGC2l80+TZlqtRpt6xbtUwOn37W+Bvlu9C/Fbi4dCH0vI6YshtdCP39nD5L80H6jDpyyn5duyYGT5qztGDRkmU3rPpt0bUrYZer1/2i8WdNWrQZ2qdbB2v5nMZOAP3u//exP7nzFSw8aPysxQpu6NipqkZC7qa1q5Tet3PrJpXTArqLW+48t27c+EOLrW+9/c67xgaL4PfTfJDuFWPVVnUuhYaej+l9TZMuQ6ZkyVO+rx0KatPa3sXQ8+d+P3vmlDl2e19ft/mpu3YGjB3c96lE4MaJUI+OhHJmh4Xenv+p96BRH9f+7EuzDx0l1e7rzz91ND8tbt+88cf1vdu3bLBf1z1esXDO9Mo163ymQJP9vrm4unu2+LFrr8MHD/huXL1scakKlavpGTh0wHffxOG/9o4Nd91bLeAr+KDxeRYoXGz10oVzrEdmmePWorx2cSycNXV8+sxZs4+bs2yD7rWONvPIV6iIscnn1UE9O/1gnWdkc7CbqI8eg8ZMUcBC93mY8WxmypY9p74XRrztFX1mrZPc+LKMn7dik56L3+bPmOKSK7fn10ay9+WLZk8/f+b0Se1MUb1bN/74Q0Gt68bRXClTp/1Az+VLRn6ZxEmSPpVHRgEofV/0jMlYgan8hYuX0jOdPEXKVJ80+LLZ5rUrlprj0DMxYOy0+cXKfFhF382//u+vv8pXqVGrXNXqtZYvmP1PrpUvvm7Vzv7cWueSPZe7h+bS4dtGdbeuX708pt8X6iOAAAIIIIAAAggggAACCCCAAAIIIIAAAtEWqN+4+fd6i76BEURQIzreSG/X623tDz/+pK7eDv9l6PjpjjrQQrbqaiHZ0fXuA0dNUv0KH9WsY17X4ujuYxdu24+H6j184syth85cVfBBi7d6c332qm2+SlSdNYeru/rpO3LyHEf9aOFa1+27RKKNYqmoHR9qW2+yO2qvz4iJs7Szw37NtNEuEEf1eg2bMGNvyOV/coyEN1YtTOtNfY1hzKyl67K45HLTm/8b9gdfaN6uc09H9fTGvcYVXpvaraL2Wrbv1ttepl33fkN0TQvtupYoceIkcndkGx13LcLvPBp6U/dXAQEFu/S86bnQ3OzjyWBEKzSeGvUaNtFuhcWbfY6ojsYlg11BobcUcLDWi8ocVE/l9ZwqUGe2k7dQ0RLq1/rs6pruh3Z7aBeGFvv1mZmUvVSFKtWs49DuIj3rrTv/MiCyZ1HPyZ7gS3eNWMYbSpDufeLKg3pffdNK3wfN1TxCzGynbdc+gzS+anU+/0qfqZx2GWkuZhmNdceR32+Et0vKiJ28PHftzgPanZEyVZq0kY2R6wgggAACCCCAAAIIIIAAAggggAACCCCAQJwK9BwybpoWPrWTQAu/ChLMXLHV2zxaZvnOgyFjjbfaHQ1CR/JsCzx7zdFxMuaCvX1RXG+fm8ERa5vLdvgHj5q5ZI3eLl+yxffooo37At80zt0xy2iRW8f1OBpH3S+//k5zMN/Yj02wrgNGTFDb2hXgqF0tBut66rTpMpjXtRC8YMOeAC3Kv5PsveSO6ulIJl2PbKyd+gwZo/Z1rI/aVXkFKvSZFpvt9bXor2t62z68tjUmldGxRfYyCo4ogBDZuHQ9qu4KbOl52egXctE8RkyBKy3Oazx6Zuz9lqn0cU1d6z966rzNB0+FpTKiFWaZ4VMXrNA17XSw1ovKHBRAUbDCHvzRs61xGWkl3rK23ejbNh3UZ9nK1T4xPzePM9NRXNayZqCtfNWatSPznL9+98Fxc5dvrPV5k+b2IJ+9rnveAl4qY+6CMq8reNO6S69fzd/1XdNYlcfEUf/aUaLrcoxsfFxHAAEEEIh9AZJux74pLSKAAAIIIIAAAggggAACCDznAkpofDL42NEzJ0OOVzfe1laS4K6tm31x//69R2//62ib8KaohNsHffftsR85o6Nt2nbrMzj0/NkzY4f07WGtf8BIVD1t7LB/FlV1TQvoWvD39927+9t2XX8xXu5P06ZJ/RrXr129YtbVcTrGKUfXHI0lV+68+XUUz+WLob/H9u3Inbdg4Xt379wJ2O+z11Hbmo8+tyYfr1SjdgPtDJk5ceSQsEsXLziqpyOh1G5E49Ub/9pZoCN+enX8/us/jR+9tf/hx5/WVb0dm9Y9FXDwKl66/J8PHz7csXnd6vDaNhOTGy/uP3U0kY4vUh/mDouIxhcVd2Pd/3+DJ8xeor0Azep+VNY8iqqisYtHgTIlJt+9bdN6e3/aYaHPiperWLVn+++aKrG6WebGjevX9e8bf1x74rlwdg7auaCA1LEjhw6OHfTksV1eJcpWCDzo52N95pS3olHzNh22b1y70npEWra/d1oEBQb4W8dvBgr8ffY4DLSZZXXsWaasLjl1JFaL9l17TR41uN+qJfPD3SHTqmOPfrqHQ3p1+SdHi4JB2oURFHjwnyCWe54CXnoWjgYGPBXYknnj737srDEsmDFpbGx/b2gPAQQQQCByAQIWkRtRAgEEEEAAAQQQQAABBBBA4AUS0NvtGTJlzb53x5aNCjJ82aLtT7Mnjx0edPjxwqt2WSQz8gwo94SdRQueWrA+4PN4wd76o1wLOmJmRP8enZzJ0aA31FVf+Sh0TNCIfj06WfMZqC0top8KORbk6PZ4FvAq5ue9e0ds3zotJKfPlCWb8mqYARx7H0cC/Pcr8GAsDhfSNS0af9O2Uw8FW6aMGtI/vDEZ3K/fjSBgobfj23XvO0R9d2vb/EszKKRjuszdHHscLPAXKFqyTICfz14jtnM1vL7V1oMHmtHdu/Yyu7dtXKfP7EnOY+quY8XSZcyctdN3jRuYwQo9Q9qxoLaVI8NRQCpjlscBi707tm6051FJmvTNNzUH+zPm7ByUT0U7Nnr82LKJ9f4q2bsCeb57dm6zzrtG/UZNdWTTyAE9u5if634rJ4vP7u1brMEUXVdujksXfj9v/9xuaQY2lI/i8sULoaN/7dU1vHun50K7faaMHtJfeTzMckr8rrwlm1YvN4JCj3/cjbIKRjoKjFWqXqu+nm2Zk7sitv/LQXsIIICAcwIELJxzohQCCCCAAAIIIIAAAggggMALIqBkxlo0VtCh6qf1vkiS9I03xg7u80+CaPOYqNMngo/ZSbQTI3GSJEn373s6UKCgg4Icq5csmO0MZS4jYKFFdCWLPm68Dj5j4qh/zuFX/SwuOR/lNjh66KCfvT0tOKd4P3Ua++KyM/1GVkZvqKuMFqPDK6uFf+NF/L06pkdllBNEARYtKIe3I0TlHu+wuOtwh4WCMzoK6s6dO7c7GsmQ1Yfq6F41+futeHmZCcrNsSnApLwSu7ZuWBvR3NS+8hs4Gt/6lUsXKthR01icj6iNqLiXq1L9UwVA5k4dN3LTmv+/oK5F87TpM2ZWPwd89jrchZAhc9ZHAYvRA3t1s49HAaWzJ08E2z93Zg46xuzR8Ut7dmz1t/XtVbJMBV3fv/fJgIXymaisgivqU8eXmcnD+3Rq+619HJ75vYo681zq6CjV1XMzrG/3jo4CSWbbGoMCEItmTRlvftb0+w5ddbxT/64/trIGqnK4eeY1g4/WseneN2vd8ZHnri0b1prPV2TfB64jgAACCMSuAAGL2PWkNQQQQAABBBBAAAEEEEAAgedcwMwjEHhgv3e9r5p/r6NorMcwZcrmklNTDD52JNA+Vb3prUVz80gk87p2S2Qw3opfOm/G5IgWXq3tueZ+HLDQon/fzj+00DE21utmMuajh/yfCliYuSV8jYXn2L4dekNdbfrsjrhtLWJny+GaWwGeht+0bq9joGZNHDU0ovFEtMOiTsOmLZTIuX/Xdt8ZJyD9syBfo27DJlrg146Cs6dPhth3UehNfS2i79qyMcKAhZkbRG//28eotmdPHjPcxTV3Hu3WCG8OzrorqNWmS6+BJ44HHfn1558eJXbXj3b3fN36p+7m7ojAg/t97H0paJAuY5asIUFHAu1BBZX9IEOmLEcP//8jkMz6zsyhSKlyFWU5c/zIp5KiFy5Z9kO1ZQ3GvZ8mbTrtEFm+cM6jBPTKfTFn9Y79+byKlmzTuG51e2AgecpUqVVHAZHInkvda5WR0foVSxZEVL5Q8dLltqxbtUz3XuMfMW3hymatO3Qb2b9n5yVzp08y68o9Zeo0Hxhf3YP29j6qVb+hmQskLnYmRTZfriOAAAIIPBYgYMGTgAACCCCAAAIIIIAAAggggIBFIKuRoFnn6WihXefzz540epgVSHkY9LujnQ1uHvkKajeE/S39khWqVFOdNb8tnOsMthalc+bOk08JpdctXzzf0QKvcby/m/I3KNeAvU1Xz/wFNQZH15zpP6IyCqAot0Jki7paTNfuh4HjZy7SkUETR/za+/atWzcjals7LHQmk72MEoc3MxbyA/39fBT0Ma8r+fPXbTp2V46Cc2dOnjj297Fd1vp5ChYprmOC/Bwc02Utp/ut33VckKMxThsz7FcdL9Tom+/bhzcHZ92btGrfRYv3g3/p3M56NFGDJt+21oL+5rXLl6qPY4cPPZH/QZ+lSJU6rQIwu7dvfiq3heagvBiOnk3VjWwOFT76pM7VsMuXNlp2fKiedh8UKla6nAJC1pwoOt5J128bwBMWrNoyZvZv6/XdqVepRL5dxmlVTz+X+QrqM799u7ZH9hwagcFcKjPHCBTZ88FY62oHhgINum89Bo2ZsniT9+Ecbh55W39Vt9q4of16Wsvqu6vv1sngoCPWzzU/HcOlnDX6PLydLZGNmesIIIAAAjEXIGARc0NaQAABBBBAAAEEEEAAAQQQ+A8JZM2Ry91YzzykI5ymjRs+0HomvqZppLfIqbP99Ya7fdpazN+/9+nF2AJFSpTW29/msTmRcaU3OtFivAIDOg7HUfmsLq7up0KOBznKh+FmJP7WLo+IFnojG4Oj6zo2SUfqKPFyZMEHv78Tb+tN+Qu/nzs7b9rE0ZH1+errr79unPT06Kgn68/nzVq2VdBjSO8uP1rn9HWbn7q//W6y90YZ+Q1k5uieeBYsXEzHe8kyov7NN/qVf8NROd2/uVPGjcxv3Etzd4u9nDPuGq+eLV/jaKXNa1c8CkzoRwvvSl6tz4287Kc0T+0usPfxQYbMWfSZo7nm8ypWUteMpO+7ozoHLeQXLlGmwpb1q5bZd/MUNo6D0g4UP9tRZ0q+rn66Dxw1SQGYrq2/blj7w6KeCto56l8+em6MGNtTu4Ks5RVAMI69yq7v2crF82ZGdN/c/x6DkWumY4nylT6aMHxAr8qF3TJtXL1ssb1e6rTpM+gzfW+s1z6u3aDR/4wbs33T2lXq87ARGIvsWeU6AggggEDcCBCwiBtXWkUAAQQQQAABBBBAAAEEEHhOBTIbC+zGeumrLm4eeeZOGTvCPg0dCXX8SGCAPeG0cgfoOJ79trfHtfiqIIiOUNKOCGdYcnnkya9yyxfNme4oV4aSgesonsNG4MDeno4VUn8H9+/b40xfUSmjRX293e/MUVM6Wun3c2dOq/3xQwf84ijJ8VNjNyZ2/+/cFOY1HeNTo16jpgrA7N76OPm1fvR2f23jmCjtWgkzsjJrN4p2AFjb1A4PN8/8hRwFkex9K7eCgj+Ojlkyy86cOHqoFvM/rtWgUXTdP/2s8TdKSj1ucN8eZhsKFnQbMGLiK6++8qqO/8qey91DOxm0W8Hej3lskaOjq5QTQ3Uc5VCJbA56dt96+513vY04ir3PclVq1HqUH8RnzxM5NZQnRTsy2japX+OjormzaPeLPdhhbcvVCFgE+vt6R1RG5TNmzZ5D35vdWzetM/K0h0X0jKZ4P1UaXR/Y46e25fNlSzNywC9dtBPGUZ3kKd9Prc/Pnz19yryu70vj79p11k4qBY0eJYx3kHg9Kt8TyiKAAAIIRF+AgEX07aiJAAIIIIAAAggggAACCCDwHxPQW+J6k1wL8/OnTRh988aNP6xT1CJqeIECvT2usn62HRap0n6QXvXO2RbTI6JTzgtd1xgclcuULXtOLcYH+j+d4yCjkStD/R0ycnDE9u1RPgi16b0r/ITb1j6NQME2vc2+ePbUCc6MRQmy7TshSn1YtbqCFvNnTBxjtqFjj34eNHpy6Lmzp3u2/66puTvCMD5h7UfHe2lnhj2IZB+LAkB6O19HMUW0WK0ggY46KlamQmV7G866V65Z5zMFVqxHJinwotwYQ3p1+fFIwIH9xslFrudOn3piLmZ/Rkwhmf6tQIF1DAqYKQfFtg1rVkQUHApvDgrUqb0gW/4LLeK75HL3VFDFflSScWLau8onooTezgTjdJ+ceS6z53Tz0Fg2rPptUWTPjcagMnOnjh9p3w1lr/vOe8lT6Pm6diXssnlNCeGTJH3jjaljh/2aLYdbbkcBwsjGwHUEEEAAgdgTIGARe5a0hAACCCCAAAIIIIAAAggg8JwLZDYWijWFB8Zb/rMmjXkid4U+11voCgY4yg3hnqeA1+VLF0KtCaFVR0cA6e+LDpI5h8eVK3fe/FpYPrjf2+EuiSzZc7mprnI32NswFs4f5dgIDjp8KLZvR053z3x6036/cWyRM2336dy2xecfl/Gy70YJr66OnDI2MDxxdFPRUuUraTF885rHxycpUNN31JQ5xsvyadt/27COjmrSfdE14+SpRzs6zB+P/IWK6m1++84Ae/8Vq9eqbyxavzl78tjhkc1LuzWUK0K7JKxlnXHPkDmbi5FuIeOm1cuXmEdb6RinNp17/bp1/erlM4xk1wrOKGeHuTvFPh5jQ8Cjfm/fvvlEPpCaxi4UBXysOT7Cm4ujORipMdKpfOj5c2es9Vq079b7nPFQKwhiz43xphEtcHY3goKBOubMmedSO0w0hh2b1q2K7H5oDCpz34ldEbI1TqS6YbaZzNhyoWO4xg/t/2gHkBJyhxrncUXWJ9cRQAABBOJOgIBF3NnSMgIIIIAAAggggAACCCCAwHMmkDlbjkeJfjeuWrbY0ZE7Og5K14OPPh0M0HE3OrbIPmW9ma7PEhlHKdmvpc+UJZsWp62f623/LEZCbR2HE14OCjOHwrEjgU8l3E6VJl16tWdNjqwF4ESJEyeJ6e1QwEL5CSI7psfsR2+y23cCRDSGBEbEwp7DIoe7Z17t0jDiEldk2aHHgOGFipUq92uPjm1Mb+NoorRq157s3CNfoSJHjaCOjjoyk2rb+9dCeuvOvwzYZCSath8dpXujHTXWOi8ZR08pgGI/1sgZ9xzuHnnVlv/fOSYyGZnT+4+ZNt84ouhk51ZNPtO1FEbWbUdzMcdgztEaMFFy+AZNW7Q5cezoYe2wsI7X2TkkNnYZqJ7V3y1P/kI6XkxJtbUzQoE8lVHQSH8ba/9/GPGTJwI34d1f7TSyP5c63krHStnrZMvpmlv33Jnggcag+mYgJ6LnS8c/WY/Zat9zwPAwI8ioQJGZ38KZPmP6PaI+AggggED4AgQseDoQQAABBBBAAAEEEEAAAQQQ+FvADEgsmjVlvCMUJdzW58bmh7PW63qz3dUjXwFzIdp67fSJkOP6XTkXrJ/r99mrtvl+VKt+Q+vnWiDWLo59O7duCu/GqIwWXi8ar8Pby2iXgj5LlDhpUv1dydg9MHPFFu88BYsUj8mN1mJvRuOsIp/dzh0HFZ2+FJAwNlg8scNCRyAp6KFrnfoMGVOzwZfNdFTWLCOfhNmHEeN5Tf++dfOPJ47wMnZYFAnw89k7ds7yDcMmz1umYJB1XFrMHzxx9hJj0ftGzx+/a2ofc8deA0dOXrR2+zvJ3kuua3ojv3rdzxv7ee/eYd814oz7P8c5Xbl8KVtOt9zj563YpHm1+OKTymYQyJzLzb8X4u1jOsc4uzEAAAmsSURBVBl87Kg+M49wUu6OrgNGTNBRZoN7dW5nP5rJ2Tlcuxr2KFdEqrSPA17vGckh+gyfNGtQz04/KHChOSvwozH3GzVlrspoLNrdYnXVePTMaUzWsSsYZX0udTzUrFXbfOo0atbSPkfNTbkunHmG7B5mHQWregwaM0W7JszP7hjbK8x/K/F5aeO4sV9/7thG91LHjOnaBdsOE2fGQBkEEEAAAQQQQAABBBBAAAEEEEAAAQQQQCDWBaYu3bBryRbfo+auCHsH/UdPned7+vpf7yZLnsJ6TTsl9HnLDt37zFyx1due42DE9EWrdF1vdHsVL13+yxZtO+4KCr21zvfY71oEt7alpMwqqwXt8Ca4YX/whU0HTjyRw8AsW+GjmnVUv/fwiTPbdu0zyPvElQdDjcX68ObkLGION4+8ard81Zq1na0T1XI7jvx+49dxMxZa6y3auC9wX0jY/d+2+R1T/wPHz1xkvuFvlmvYvHV7XRs2Zf5yc/Fcb+/rs5r1GzVVG/r36JlL1n748Sd19add935DtgWevfbb9gPH02fOmt3RWKt8Uvdz1Vu4Ye8h9bsl4PSVnUdDb2o3jb28M+7ljeTVam/FzoATuv9qSwvr1raU1HzzwVNhWw+dueooV4aCYxv9Qi6u3nv4jBbdR85YvFpt2gMEZpvOzkEBBJ9T1/6csGDVlrpffv3dyl2HTspIOSzUvp5ZfTd0H8xns3jZD6voWs/BY6fquVbwQVaOxqMAiNrXd6xJq/Zd9AzLwTwyzRyvAgyqr7wezjw/CqLsCb50d8byzXuVdLxSjdoNRs1cskZtzFm9fb9ymJjtaHz6fMDY6Qs0lp8Hjp5sXlMAUdfyFylR2pl+KYMAAggggAACCCCAAAIIIIAAAggggAACCMSpgBY9i5etWDW8TiYtXLNtzb4jT+yuUFmdzb/7+MU7WvBUcMJ8W9tsR8cKaYFZ180/U5es32nmXrD29+PP/YdqMVULvI7GocCDFqwXbfI+7Oi6dmdoV4D6UTt9RkycpUXwmMJpIXhvyOV79gBLTNu11l/vezxU47V+VqpClWr6XAvcCghpfvY+Nb8R0xau3H3swm1zN4QZQFCgRc6zVm71sfqb7dnvlbVtWZv3Q3MfM2vpOjPBt30Mzrhrl4rGqUDFlMXrdpjJ1e1tlShX6SMFU9p06T3Qka8CLgrimPe4S79h48wdHvbyUZlD45btOumZeRSEGDJumgJDGot+V+Crz8hJs5Xrw+xDbWuHitV1+rJNe0pX/KiGo3Hr6C2zrAJ7jo7pUtBBc7PujIjsGWvQpEUb6xhW7j506vNm3/1g31Gj79Qm/5OXVVaBMeuxWmnTZ8z8KJhhHNEVWX9cRwABBBBAAAEEEEAAAQQQQAABBBBAAAEE/nUBvc3t6Mx9DUx5JcwcGI4GqhwSWvzVwr+Lq7tneJNRTgUdvRTRZI38yBnCC2iY9bRwb327PKZ4ypPgnreAV0zbiai+dhvIOLp9WBfttTtAQQbrorXuj2d+r6IKIEVlx4kclbDZmXHFlruCBRGN0Uh1kU6L++Hl5rCP1dk56Lkyc6TomCkFabxPXn2onSrhzd/FNXcejUWL/pEZKbj3P+OYr/DKaWeM2oqsHft1OWhHivK12HfgWMuqb+UOcdS+Aj8RzTOqY6I8AggggAACCCCAAAIIIIAAAggggAACCCCAAAL/px0MOhIIiugJ5MqdJ//ynQdDzCOxotcKtRBAAAEEEIiaAEm3o+ZFaQQQQAABBBBAAAEEEEAAAQQQiOcCesM+W07X3IEH/Xzi+VDj5fCU62HiwtVbfffs3Kak1of89zuVADteToZBIYAAAggggAACCCCAAAIIIIAAAggggAACCCDwbwno6KdHiZuNpNT/1hiex351bJQSyytfRf3Gzb/XcVo6VktJuJ/H+TBmBBBAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQT+VYFK1WvVV8DCLU/+Qv/qQJ6jzpWYfNHGfYFK6J7Pq1hJDV25KeSYO1/Bws/RVBgqAggggMBzLJDwOR47Q0cAAQQQQAABBBBAAAEEEEAAAQSeEsiaw9X9z4cPHxpnGfnBE7lAhszZXMbNXbbh9u3btxpULVXwzMmQ46qlJOtyPHzQzzfyViiBAAIIIIBAzAUIWMTckBYQQAABBBBAAAEEEEAAAQQQQCAeCWRxyeV2IjjoyB1jAT4eDSteDiVR4sRJhkyas/T/XnrppWa1q5Q5e/pkiDlQz/xeRY8GHjyAY7y8dQwKAQQQ+E8KkHT7P3lbmRQCCCCAAAIIIIAAAggggAACL65Aluw5XI8E+O9/cQWcn/nnzb77IW36jJl7tGvZxBqsUOLyAkVLlvHz3r3D+dYoiQACCCCAQMwECFjEzI/aCCCAAAIIIIAAAggggAACCCAQjwTefOt/bydLnvJ9joNy7qZUqlGnwYljRw9vXrtiqbVG3oJFisty5+b1q51riVIIIIAAAgjEXICARcwNaQEBBBBAAAEEEEAAAQQQQAABBOKJQObsOV01FB1lFE+GFG+HkTDhK6+kTpsuQ9DhAH/7IKvV+fyr27du3dy1ddO6eDsBBoYAAggg8J8TIGDxn7ulTAgBBBBAAAEEEEAAAQQQQACBF1cgy98Bi6DAAAIWkTwGDx8+eHDv7p072klhLeri6u5ZrnK1T5cvnD39rpHA4sV9mpg5AggggAACCCCAAAIIIIAAAggggAACCCCAAALRFOjUZ8iYjX4hF6NZ/YWrNmDMtPl7gi/d9SxQuNjriRIl9ipeuvyafUfO7goKvZUmXYZMLxwIE0YAAQQQQAABBBBAAAEEEEAAAQQQQAABBBBAIDYEpi/btGfsnGUbYqOtF6GNFO+nTrNsh3+w7+nrf5l/vE9efVj1k3pfvAjzZ44IIIAAAvFLIGH8Gg6jQQABBBBAAAEEEEAAAQQQQAABBKIn8HKCBAmyZM/hunDmlHHRa+HFqxV6/uyZ2uULeyhnhYtrbs9rV8IuL503fXKgv5/Pi6fBjBFAAAEEEEAAAQQQQAABBBBAAAEEEEAAAQQQiAWBt99N9p52C2TN4eoeC83RBAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggAACCCCAAAIIIIAAAggggMCLJvD/AEZzzx0bBJeBAAAAAElFTkSuQmCC"},{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO2dd5gcxbW33+6enGdzDlrtrtIqrHIOIJLIILBJxmDA/mxz7euAA9jY+GLsaxvHa4PxBWN8MdkiipyEUM5Zm3OenZynvz9aWhCspBFISLD1Pk8/0k53VVf3dP/m1KlTpySdTrdVVdVKBAKB4DBIklQnKYoSSiaT5pPdGIFAcOqiKEpYPtmNEAgEnw6EWAgEgrQQYiEQCNJCiIVAIEgLIRYCgSAthFgIBIK0EGIhEAjSQoiFQCBICyEWAoEgLYRYCASCtBBiIRAI0kKIhUAgSAshFgKBIC2EWAgEgrQQYiEQCNJCiIVAIEgLIRYCgSAthFgIBIK0EGIhEAjSQoiFQCBIC93JboDg2LBYbej1elRUouEw0Wj0ZDdJMEIQYnEKYzBZmTF/CTPnLmDMhIk4nQ7isSjBQABZp8NmsyPLEi11e3jntRd58dl/EwoL8RCcGMRSAKcgNnc2V9/0TRaftogNq17l3TdfZ+f2LQwOeEip6iHH6vRGRo+t4bRzL2HRovnc+Z2b2Lx150lqueCziqIoYRRFCQGq2E6NbcLMJeojL7+rfu7KK1WjQXdMZYsrJ6qPvbpGzcl0nPTrENtna1MUJaTIsvxDVVX1CE46ZeOm8bNf3Ml3r7+Md1atJplMHVN530A3xoxiRuXZ8ET1/OHBxzAmfezcufsEtVgwUpBlOSF8FqcQX/3+z7j71q/T3NpxTOUkWcHhdCIBiXiMzIwsbvrOFTzzz/u4/JobePGl1z9UJhaNEAqFjlPLBSMBIRanCnon1cV23l2/7ZiL5hRX8r0f/wRJ0v6WdQYmTZqIXZ8gt3wct//mzx8qs3/zKv70+z983FYLRhLCZ3FqbJLBpT7z5mpVOg51ZZZNUO+9/34V9OqKN1af9GsT26d/UxQlJIKyThHU2CDb6/q48IJzPnZdOTkFdHd3YM7IJzjQfRxaJxCAcHCeQmxc8zb/77b/pmbcaDrbWvB4PB+pntLxkynNMNMdUCnKtvDaK68d55YKRhrCwXmKMdjTxleWn8Vp51/G13/0a/Jys2hp3E9rYwM93Z309/bR39vN4EAvvT09+H2+Yesx6BUS8RSTps5gy7o1AOiMVm7+/o956A//RU+/95O8LMFnBCEWpxjJRIyXnnyIl558CIPRTElFJSVlo8jNL2D0uBpmZCwmMycXd0YmVquVtsZ9PP/EP3nlpZeH6kgkUiiKzJwFC7jrq78D4JwrbmLGnHm0bp/PY088O8yZJSrHT6SvowmP5z0xsdrsBAP+4RsryVgsZkLB4LC7TVYX5150Ec899hDhaPyI1200WbDZrfT39h75BglOHsLB+endZEWnVtZMVX/z4DPqjTdeN/R59fTT1fsefUb964P/GPps+Y3fUV/csF99fvVW9em3N6k1Y0cfUtdNP/yN+ucHH1UfffFN1WExqIBqyypSH3/5LVUnoTryK9Sf3nXnIWWWXn6Tesv3b1EB9dwv3KwuXTLnkP23/uFh9Z/PvqWeu+x0FUlWv3b7b9XnVm9VayeNO+S4S770n+oTr65R7330BfVP9913XJy8Yju+m3BwfspJJRPs376Rn3zvm5x+/sVDn3c01zOudhZP/uO+oc8eu/e/2bhtN7d/9fM88fRKKipHDe0z2nM4+7TpfO0Ll9HmiZKX5QTgjIuu4M2n/4+ECrn5xdjM1vedXeLSz1/Fk//3dwDKR1UhoQztLRo7naocHc8++zJGs4mzP/8ViuwJfvf7PzFr1tyh4+accwWnz53EVefM5ytXXshdd9yBemDf4jOXHce7Jfi4CLH4DJCZnYdvoH/ob39PM/vrGti6ZcvQZ9XTFlPsSLJp224KCorobG8f2nfxF75MoKeTCXPOIksXor6tF8Vg4fKrv8DGNe8AkJWbjz80OFSmatoiyjIV6pq7tP15h+6/6IpreebRf2DPciHJNq79wuXcdfttmE02/OEAcMCP8t3vc99v/4twNM5513yds5YuAGDM9NO48qrLT8DdEnxUhFicisg6LrziWjIzXEc9tKB8DLfe8V/c/+f3B1ilePrJJ7nquhsAMFpd3PLjO/jtHT8kkVSxWq1EgmEAyifM4IJzFmMvm8TXv34D3//aDSRT8IX/+BH5mQ7UZAqQOP2c8ykurtDqszj47m0/IRHT/BC2zHxmzpxOyYH946YvYfr4YlaseJbMzFzOveI6nvrb3Qz6w+j0RlQ1CcB13/oJxXkZhAJ+dEYL51+8nFQiiawz8p8//BF//tXPj9MNFRwPxKzTUxFJ5tLrbuaSyy6nv7OJrRvX09zYQF9vD6qqYrY6KCotZ8qs+RTkuvnzXT9mzdr1h1ShM1r59QOP423bS3H1FN586m88cP+DAJx9xVc5f+ks3lmzifMvXc5P/+NaSqYs5eLzlvDcihWMn76QXFuKx1a8wg03XEtrl4eUtxVH6RR6G7YyasJ0nn/wd1QvXI45PkBx9URefPJhLr3qi6x643WmzpjOD79yFY0tHdx1/zOML3Vw6RmLiSZSVE1dyE9/eht1TV1Y8PHCa+u4/ktfIJZUUNUEr/7fPcQzq6nMhp/++Kcn4eYLhkNRlLAQi1MYSZIprRzLhElTKCmvwGazIUkQj0Zoa6pn+6Z17Nm9G/UD09YPouiN1M6ci7+vnT179r6/ZuadcT6FeZm8sfJpunv6ABg3dS6TJ0+iq6WON199mWRKZfS4yThtRjatX4vR7GDqrNm0N+yhqakZRW9k6ux5dDfvo7m5lcKyKsrLS9iy7h0CByyX4ooxSPEALS1tQ2evqpmKw6Jn07q1pFSVnIJiUrEwp196A9XlhYybOIYvXbIMf0jk5jhVEFPUxXZKbVd85VZ11Y4GtWZc5Ulvi9gO3cRoiOCUQdYZmbVwIQ/98S6279p/spsjGAYhFoJTgktv+BYTqsvx9Pcf/WDBSUGIheCkY8ss5LJLlvHwQw8hS+KRPFUR34zgpHPh1TfywsP34AtGkJBOdnMEh0GIheDkIulYdu4yVjz+ODrFQDx15DkkgpOHEAvBSaV4zFT8rdvp84YwORyE3hcFKji1EGIhOKmMnVTLtk3rAMjNzaO3UyTrOVURYiE4qWTnZdPT3gpIVFZVUF/XcLKbJDgMQiwEJ5XBgUFyC4uZvOBcYt276fdHTnaTBIdBhHsLTipWVw53/vE+LEqCO2/5Oo0t7UcvJPjEEXNDBAJBWiiKEhbdEIFAkBZCLAQCQVoIsRAIBGkhxEIgEKSFEAuBQJAWQiwEAkFaCLEQCARpIauqKgRDIBAcEVVVFVlVVZFAQCAQHBFVVUVaIoFAkB5CLAQCQVoIsRAIBGkhxEIgEKSFEAvBiESShF//WBFicRjKK6uZs+h0KseMP9lNOe4oOh21M+cet/om1k4/bnWdSBSdjuVXX8+Ss85j3pIzcWdmfegYu8PJmAmTTkLrTn10J7sBpyplFVW8vvIZCopLT+h5ZFkhlUqe0HN8kOmz55NMpY5LXZIkkZWbd1zqOlYURSGZTP/eZWRls3n9u9Tt2XXYY8pGV9HZ1no8mveZY0RYFrIs43JnHFOZZCKBwWiko7X5BLVKo3RUBQAGo/GEnucgkiQxpmYyXe3aC2GxWj9Wfe7MLAYHBob+nrt4KWaLlamzjp/l8n4MRiOSJCFJEu6s7GMqO7pqLK1NR87xmZ2Tx0BfT1r1OY/xmfq0MyLEQm8wYHe6jqnMlg1rmDR15tDf+UUlAJjMFgxGIyazBVmWMRhNOFxuAAwGI3kFRWmfQ5IknO4MJEkiJ6/gmNr3Uampnc7eHdsY6OvF7nBy3qVX4MrIxGK1odPpKCguxWK14TxwTS73gX16PVVjJwDaL3ReQRE6nZ6yikoa6/ZitdkBePfNV7HabGxauxqrzY7FZsPhcmMymY/LNdodLpAkjCYzDsexfafZuflMrJ3B1FlzkSQZnU5PUWk5E2tnICsKU2fNw52ZRSqVYtzEKWRm5RyxPnfGh7sxn2VGRDdErzeQmZ2DwWDEaDLh8w4SjUSIx2IkkgmAA39HsTucSLKMb9BDZrb2sCw4/WxSqSQWq42qsRNIJhPIskzd3t2MmziFotIy/vLrn3PaOeejqiorVzyeVrvMFguJRAKzxcLYmsmcc9Hl2B1OQsEAoVAAm82B3+elu7OdgM+Hd9BDKBQg4PMRDgWRJJmMrCztxXG6CIdCgEow4Mfv82r1BIND5zMYjVitdryDA8iyjKwoJBLatcycvxij0Uh5ZTWb172L0+Vmx5aNVFSNxWK1EgoG6O/rRVEULr/2RrZuWMuoyjEYjEZmzF2IyWRmxaMPMWvBEiZPm8WTD/+dmslTkRWFDe+uYs7C00ilUrz0zJMYjSZKyisIBgOkkkkUnY5UKoVOp8NssWIym7FabVhsdiLhEIqiEIvFiIRD5OYX8u5br2GzO7jmyzczONBPNBpBkRUMRhMBv5dYNEpnexvdne00N+zH098HQGd7K+tXvzV0P8orxzFz3iIeffA+Tj/7fDasWUX1+ImMHjMOVVWpGl/Dmrdew+5wIisKeoMBg8FIKpXCZneQlZ1DU/2+4/SUnvqMCLFQVXVIKDKyssktKCQeizHQ10s0EsHr9RAJhQCYNmcBr698BoBgIIDVZiOVTNLe2oQsyxQUl7DikYeYMHkqeQVFdHe2Ewz4KSotx2Z3sH3zBgCsNjuujEzsDifZuXnodHpcGZkYTSb0egPJZJL8wmIa6/YSjUSo27OTV577N4qioKoqAIpOj83uwOF0YbM7cGdmMqqyGpPFgixJgITf78XrGWCgv4+Az6e9LLEY0Uj4kP58Sflozr5wOS2N9ZRXVpGZncO2TevZs2MrA329ZOfksW3TOswWK43791JQXMLYCZN45fkVLD33Ivbs2EZBsWZdBXxedmzZSEnZKJacfT5//d0vmb3wNIrLRhEKBsjKzcPr6Wf0mPHc+7tfMKpyDBaLle1bNgIQjUao37ebvMJiykdXYbbasNntRMMR4ok4wYCfcDhELBZDVVPIig5ZlnFnZlFUWo7VaqO/p5u1b78+JMwqIB3890A3xWg0DV2/3mAgHosd8lyMmTCJV577N2oqRUpVsTuc7Ni8nklTZzLQ38fbr65EVTXxdbjcOBwu9AYDiqLgcLnJLyxGkmXU4+T/OdUZMWJhslhY986bRz3W+D7fgdlsJr+olI62ZqrHT+KtV144MOSm0tfbTe2MOTzxz/uZNmc+WTm5vPrC0wz09QIQDPgJBvwA7NmxddhzzV54Gj2dHRjNZuKxKKqqkkgkhvYnk0kGopG0+9BHIjM7h2efeJj2libsDieVY8dTUjaKlgN9eKfbTU9XB7n5hYyfXMuqV19i1oLFFJaU0dvdSV9vN+Mn1ZKTX8j2zRsYWzOZXVs3UbdnJ7FYlFg0wpgJkwgFA9Tv3UUkHKa5YT/JRILS8gpeeX4FPu97q42lUik6WpuP2Sek1xvo6mhDURSc7owhYQVNKED7vlUgHHrPqiofXUVLY/0hdYVDQbo62nC5M+nuaOf85VfywJ9/izszm3feeJlEXFtKMZlM4unvG7JQQBOkpedeNGKEAkCRJOk2QDnZDTmR6A16SstH01i396jHJhIJJkyZRkn5aNpbm2hpbGDG3IXU7d1FLBKmpbEei9VKV3sb4VCItpZGHE4XXe0tTJo2i3gsdshLcSSqx0+kfu8ukonEUNfoRDB11jz6erpoa24cukanK4NwOETNlGk01+9Hp9OjAnV7dmK2WGlvbaKopJyMzGzWvfMmC5eeg6e/j6ycXHILiujt6iTg8+Id9Gh1xuM4nC66Ozvw+QbxejxD1ls8HqdmyjRCweCQgH5UMrKyaW9tJpVK0dvdlXZ9ufmFVE+YSElZxdAIl9czoHVjYlFqZ86lo62F+n27sVhtVI4Zd0RnqCzLmC1Wero6Ptb1fFqQJCmFJElRNFH+zG46nU51ZWSe9HZ8cJNl+aS34Vi3OYtOP/I1KToVUCVZVqUTcH0Wq+2k34P3rlU56W34pDZJkmIjYjQkkUgwONB/TGWcTiclJSXY7fYT1CrNFP8kkAHdcQpYlOUjPzKKohmpJ8o8DwUDJ6Tej0LqGGI8PguMCLH4KGRmZrJo0SIuuOACTCbT0QsAOp2OvLw8Jk6cSEVFBQaD4QS3Mj10MiwpAP3H/LZlWT6q6MZj0aH/j6T+/EhgRPgsPgp6vZ6ZM2dSWFiIx+Ohs7PziMc7nU7mzZvHRRddxLRp00ilUvh8Prxe7yfUYtDGAz5MUoUcMxRaoTU47CFpoaoqPV1Hvg+CzyaSJKVGxGjIR2FgYACPx0Nubi6jR49m8+bNw3YbJEmisrKShQsXMnHiRAwGA11dXaRSKQYH03N0HglZgkwTZBghpUJvGLwxrSP5oWMVhVQyMcwe2NgH11RBH+B0gdMKq3ZAJDbs4UfFoINFk2DRZK2NvV749ztQfwz+PkmS0BtMJBKxI5r0kgTqcBcs+EQRYnEYEokEL7zwAsFgkGg0islkInQgFuMgsixTVVXFnDlz0Ol0BINBIpEIjY2NbNiwAZ/P95HOLUtQWwlXnQazq2FUBjiBRDf49sD6dljRCI83wuD7XvbDCYUswdyJsPxS+MVY6BrURCKRhJvuhi31wxYbFp0C06vhO5fBzLHw5lbY3w5jiuGNX8Njb8LPH9bE42i4s3KZMH0RbU37ady96ZBh0DHFcOVp2n0wGmDNLrjvBWjqSr+tguPLiBILSZLIyMhAp9Ph8XiIxY78s9rT08O2bdswmUzo9foP7TebzRQXF5NKpTCZTLz55pvs2LGD7u7uo9Z9OEblw1fPhy/OgmQH3PMivNUFkgIXz4NLlkLzozArF26ugd9th7/vg8Qwv7wSMLZUe7HPmArPvQN/fhie26NZKV88E576CVz3K3h9y9HbZjfDL2+Es2fAn5/WhKbP+56VU5AJN18EK++Cq34Ou1sOX5esKExfuIypC8+jvWkv3a31BP2aJTZltFbH29vhibehox/OnQWrfguf/xm8veOYb6vgeDAShk4PboqiqBMnTlS/9a1vqcuWLVPz8/PTKmO1Wocd5jQajeq4cePUmTNnqtXV1arJZPpY7assRL33q6iPfw71ngWo5fYPHzNnPOq2v6J+8UzUyZmor5+L+uxZqMXWQ4+zmVF/9kXUnsdR//INrW63EbUmz6YajOah406rRW36J+rpte8vLx0cLhv6rDgb9YWfo67+PWp10ZGv4/qzUev/oZ3zcMfIiqKeufxG9du/+pd6xdfvUE1Wuwqo2U7UDf+D+u3lqIp8aJkFE1EfvAXVbj75z9JI2yRJio0osQDUsrIy9dZbb1Xvuusu9fbbb1fLy8s/Vn2KoqjKRxhv1+l0qtPpVHU6LS7BqEc9fwrqDRNQFxegGuXDlx1XitrwD9RFk1ANMuo3alC3XYo6NxdVAnVMMepLv0B99/eos8aiypJWriAnW732hm+on7vpFtWVmTtU34Ia1P1/R509bujBOOR8GXZNKB69DTXLmd713XCOJmqTKg5/jCsrT62df45aUFatAqrZgHrft1D/+X3tfgxXxqBD1etO/nM00jZJkmIjbjTE5/MRjUYpKirCbDZjsVjo7u4mEBh+/F6StP7zBfMULlyUxeKJcaZWpjAboHMA4gn1kL720TAajVRUVHDxxRfzla98BY/HQ0dHB9FYkoAPtvfBrkFtBGOY1gCaP2BnM/ziBnhtKzxXBzs9cPdsmDIGbr4WtjbA1XdBY5f2bVc44GfzHYxediPlE2fS291J476dADT3QF073POfsHE/tL0vujzPDX/7tubjuOG3BmKyC5PZTiwW5khex60H/CC/vFHzaQzn+IyEAnS21OEf7CPLCX/8uuYPuem3h/d5JFMgRmQ/eSRJSo04sVBVlfb2durq6jAYDITDYQAGBweJH5gLAFr//PzZcN1Z8IWLxnPG8tuYf+73mDjrMgpLqjn7jLksmynhUlrwBlX6j+DLlCQJl8tFeXk51113HbfeeivXX389NTU1xGIx1q9fDxE/gQT448OVl6maUMuo6gn4fR5ikTANnWAzwy2fg0114EmCZTR87SqwtcEbL0MyoY2iXFUJd86ATd1R9lknkF9YxPaN79Kwb/fQOeo6tJf6vm/B5NGaSE6t0l5gbwCu/42Ogsq5LDrvaopGj8PT00nQN/Dhxg7dZ1i/F3Y0wr3fhAllsLcNBj5wn3QKLJwED3wHInG47A5o7U3rqxR8gkiSlJIkSYqqqnpqRA99wuh0OgoKCpAkiZ6eHsLhMBKwYCLcdHEWo8fOQnXMJn/scpKqHp1OR1ZWFqFQiEQiDskwicGN7Hr9Rzz7yi7+thIC4UPPYbPZqKmpYdasWSxevJhFixZhtVqRJIm+vj7uuOMO7r//fmIhzbKJDfOrabbauO6bPyWnaDQb3nmNlx7/K9FwEEmCL58L31oOBj00d8FvHof9u+GKCpiTBy4DbB+Af+yH19oht7iM2QtOY6C/l307tzHQ33dIVGSOC65ZChfNA6MeHnkDfvckoJhZcN41zFl6CeGgj5WP/IXta19J6z4XZsF3L4ezpmuWTteAZqkoMlQUQHE23Psc/HEFhKNHr+94Ix1YPkdVhclyOCRJio9osTiIJEmoqooswaUL4aplJRTNvgtz5kTy84tQFIXOzk70ej3Z2dkEAgEcDgder5eBgQFsxjh1b32fTWtW8ot/qfQd+PVUFIXa2lqmTp3K4sWL0el01NbW0tXVxVNPPcWrr77Knj17CAaPHCklKwpnXXQlUxeczfbNm3j1qfvxD743A9Jm1l7swYBmphsMRhKJBJKaRJYg/oF3oKS8ArvTRW93J0G/f9jJWPKB+K6U+t49qp4ynzlnLCeZiPPsQ3fT33Xk9HOSLOPKzAUVPH2d5Lq1kY6SHHDZNOtldzOs2wNdniN/R8cTRWfAas/GYs/EmVGAxZGFpEp4+1vx9rfh9XQQj4WOXtEIQojFB7h6KVxzQRW2MT/AnjcNVVUpKytDURTa29uJRqOEQiEaGhpYunQpZrOZQCBANBol4BugY/2P2L1xBbc9AB6/9oKNGzeO0tJSRo8eTSgUIhwOs3XrVhobGwmFQmn5O4x6yMowM2vGGNR4gMb6Rjr7E/hDWqxESoX4gRALs9XG5BkLUFWVrevfJjzMXApJlrnw8qvJzS/gledXHDEn5fvRG0wUlI8hHPDR096I5g05PDZHBpfe+D1MZitP/O0X9HYcYSz1E0DRGcjOr6D2zEpMtkz8veXIOhOKTgdIxEJ+BjsbCAz20N60Cf+gCOo4iCRJ8RHnszgcCyfCD/7jAlKFN1MxYQmZmZno9Xr0ej319fUYjUYKCwtJJpPYbDYSiQQulwuDwYDJZMJosuAuXowS2km+pYFV27WXeGBggP7+fjZv3szGjRvZtm0b3d3dh/hHhkOStCjL4mzt3+7+BDv2dNPSNkAylUIGLCZw2zUHbGWhJhzonZx92Y2MmzqPkM9De3PdhytXVYpKyljz1utcetX1bFj9dlqJb1PJBN7+LoL+9MwAWVGYtvA8sgpGEfAO0FKXXoCEwWRm7JQ5uDJz8A/2H1NS3sNhtroZO+18qqbPZ/zpg7iLu/H1KiSiThKJGIqiIyX1kVHSj8niwKQvwutpJxE/MWkDPm2MSAfncLhtcOfXKnCN/w4t3QlqamowGo2YzWZSqRQejwe3243NZiOZTJKZmYnJZMJwIGtSMBikubmZouJSXEWL0A08QXevn/oOzaEaDoeJRqMkk8m0LIkclzYq4LBAQyd0D0LiQFcingB/CPxh8IU0C6ajXwuOynJCjlPFlVVARnYeTXV7aGk4NO2brChk5hbQ192FJEvU7d3FojOWsWvbpuN+XxOJOOFQCIPJTMPuTfR1pmdZlIwaw8Vf/CajJ0wj5Ouls/3jWSQWWyY1sy/FnV9OStXTsU9Hxz4ZnVIFKR0SEgZrF1nlHagpE9UL2gkHUhAtwtPXivoJZ18/FRFicYArT4NzLroBe/FZTJ8+g2g0isFgQJIkPB4PeXl5RKNRBgYG8Pv92Gw2FEWhra0Nu92OwWDAZrOh1+uRFBO9vR7KLatZuR7ix/icuW1an76tF/a2plc+pUI0rg03dvQl2LdrJ4p3PU37tuHxHWrB5BSWc/6VX6W6ppa6XZtoqt/H6eecz7ZN64YyQx1P+jqbadi1kZ72hrRnoRqNBqrGTcbmcNC0dxsdLUfOyH0kJElm/MzzKBg7mtzqOlKpLpLRYiRyIKUbshziEfD3x1DVejKKVBx5YYIDKopaxGBfC0frcn3WEWIBWE3wvWsyKJz2Q4rKxtPS0sLq1asZM2YMoM0+TaVSBAIBDAYDiUQCi8WC2WwmGo1iPJCaXlVVYrEYFouFuJyFr/Ex+jwR6o4xkVIsro0W+ELgNMB4FxTZYJwbjApEEsOPmLyfeDyBSRpEJyfo/cBcNp3ewJjJs7A7s+hpb6K7vYWB/l4Wn3UeOw7kyDyIhJYHw6IDt/G9Ke7DhZYfHpV4LHJM09VDgQDtTXvZv2MDe3ds/lgiZnflMfuiEkqnNmHP9uLItmFxgL/XjSwrKHoDBrNKOPo82eW9mJ1RAv02QoMKSbWfZCibcCBEJPzR5vl8VhCzToHlC2H0+MUYHeWkUilSqRTTp08nkUigKMqQz6KyshKfz0dGRgZ9fX04nU7y8/NRVXVo8lhBQQGxWIys3DK6Kq/jytN+w9vbIXgM3d6UCgYFblwA3zoH8hwgJaGvBbytEAnDX/fAQ/shcIR3aMCvOUY/iLe/m+f/dQ+FZVU01e0BYP/unZx53iXoDQaS8RhFVjijCGbmQJEVCiyQYdLallRhaz+s6oJNvdAc0Ka9f3DEBcBotmKzuxjo6zwmsVDVFG3NH7YmjDJMz9aGgr1p6kduQTWuIh+qFMbTYad33yRMjsq44/wAABmPSURBVBiKTvPpq6kUAW87iVgmnbvGEgrup3hsCWoqhCvLSTi3C1dXMYP9YuGhEScWB62AgyyZDI7cGnQ6A5FIhEgkgvXAwjsH18OsqKhgYGAAl8uFJEmYTKahjFCSJGE2m6murga04dKuri5ipkksnOrCaR08RCwkSUKv1w8lxlFV9ZBRkXwH/PEGqBkHf30FWno1X8S5M6GwCv7yvzDRDU8sheUvg+8wL43JKFFeNQEcKs11uw9Z9ay7rZHutsZDjq9f/Ty/+vJFVO9/hAon7BuEl9rgwX3QGtBiIgByTFBqhzI7XFsN1S6IJbXJbC+3Q8v7Bl+mLVzG2ClzeefFR9m96Z1h2ynL2n080qpsMppl9dNpYNHD5emFd6DTm7C73QQGe3HlZ9NcP4141EC8V4eqqgeehSQ6vZnc0W5iIT9R/0RUNuEq8tDfFiaRTGB3ViLJyoj3XYwIsbBYLBQXF5Obm4vb7aa3t5f6+np6enpwWFXMzko8fj86nQ6Hw0F2djayLBMOh4nH41gsFnp6erBYLFit1qEXO5lMIssywWBQS4LrdAJgMBiIJQ1YXGWYjdp0TqfTSUFBAeXl5YwdO5bq6mocDgft7e08+eSTbNu2DX3Czx+uA08U5n9Lc2we5I//hovmwp03wB+fgmAH/HMJfP5VCHxgZnqmA+ZOK6Jk3k2MD8Z5/tEHUFNxers68Pt8Q8FHMjA1G64cDZeWbaBxyiX86flHeK0N+iIwnC1Q74N33xcObpBhYgZ8aQx8fQK80g53b4P2EERDQfQGM2VVE9mz5d0PWRcGo4l5Zy4nBax55SkioUOHeWWgxAa3T4P5+fBME/x0k5bPIx1MZgdmF0R9NXTujRKLRDC7fESDKVKJXEjJSLpuisfuIb8qRjKeorthN1tfKCCnPEYiOJ6oL4msBJGQRrjXYoSIhdVqpba2llmzZpFIJPD5fLjdbt555x0UeZBkPEifvw+TyURRUZGWObq3l0gkQm5uLl6vl3A4PJSqX/e+RXEOOj51Ot1Qvk6n00lGZhZSVAv00uv1LFiwgHnz5lFVVUV2djZut5vc3NwhoQl6ullS5OfNvZpFEfmAxZBIwmNvabknnrgd7n4MJA/8bSF86a33wsRnjYX7vg1re8ppMWeR4zQybuJkujta8A16sNod9He2MiVT5UtjYHEBPNkIi56G6Uo9a6iiN7ofs9VKLBrVIlWPQCwFG/pgwyrIN8O3J8FLy+De3fC39a8QiYTwDvQM2w0xmiyUVNVgc7hpb9zL/u3rtM9lWJAPN46FyZmwognOewH2DA4vYIcjkYgS9sm4ClpJRHPRGYyEvaDT20kmQZKBlBOVAP7+FPYsE7kVBkpr+9j+SiESJrIKi+mu24I64qVihKTVkySJvLw8dDodOp2O+vp6+vr6aG1t5cI5cVx548goPZ1gMEhGRgapVAqDwUBmZiaqqtLf309ubi52ux2fz4der0eWZVKpFKFQiEgkgtvtxmg0snv3bvLy8gj4BrAN/p17n/bj8UN2djYVFRWEw2H0ej2JRAKv18vOnTt584036GnaRPtgjKfWvTdMOhwDfnhhPdzzDfj7VnBF4buTIZSEMxZpcznueRZ++XAYi91NT3sTe7etZ/zEKUyfM59I/VrumhTgmiot/Pvm1bCiGQai0NrSxLKLL6enu4vPXf8NikdV0rhvV9oOxkBC67q81qFZGleMStLQ1MTm5t6hSND3E49FScYjpFIpGnZuwJ3ycWk53DUTLq+Atzrha+/AU03QEzn28YhEPEZGVgVqchbRoJ2KOavpatpLLFCETm9GVVNIkpH+ZhfxqIFEohtXrhF3gUrTliTu7CnEoyG8XY30doyclceGY8Q4OIPBIK+99hqrV69GlmVisRjhsLZil8cPgd7tWCvfuxXNzc3s3LmTs88+m0gkMmRFHKxLVVUyMzPp7u7G5XLhdruxWCyoqorNZkOSJOL+eryeLiIxLYv32rVraW1tHRpdUVWVVCpFNBqlv7+fRDye9svQ1AVX/hwe/RH88G8QS8D/fhcUF2x5BSK7YIm9l9Db95CSdMw0qywrm0nJ7t9z5S3fZP+al1n64CoGPjAPw+sZwGZ3YLU7yS4sI79kFJvefYOGvTuP6X7vGYRLX4bzSjUh+9IY+N+9mjj54tpLL0tgkFMM7n6bqsE13FkV47RC2NgL/70V1vSk3904PCq9nfvILhlHLD6A3hinbHKKwc5teFpL0etLQZIwmLIJ9jkxO7sY6AiSTEjYHLNBVQl5evB5OhnpQ6cwQrohwJDz8oM88y4U5b1JvHA/VWMnoaoqRUVFyLKMx+NBp9NRVlY2lH8zHo8PRRT6fD5yc3MxmUxDfozS0lK8Xi916/9Cf0uSgQPTLuLxOM3Nw6++JUugKAciMNNkwz4tG9VPrtGiOP97FTzxEkyywYwcWFasEk2FSaQ0H0jTqhXcu2OQtU/8hIuuu5nyKTCwZtWH6q3bswtSCVY+8XfcmTl0d7Sl36j3kVTh303wXAssK4Evj4VfzoLOIESTYNJBlglApScc47V2OHel5lg9tqHZI+MdaCfk7cVpLaNlWzNTzsnEYFJZ9+96vK3F2qiXTo+sgDPXiM4QxtebJBHzoyZ0RHwD9Pd89DiPzxIjfm6IUQ//+22wVlzP4uW/IZlMotPpGBwcxOPxUFZWhsFgIB6P4/V6cbvdQ92UVCpFd3c3yWSS4uLioZGN1W89T2TzNfzhqRRvbkuvHbpjEAtZPpAZJ5VCkrTkudHhprYf+PeD754ky3z1O7fxr/v/Ql9P9yH7ikrLmbVgCY//42+8t3poGkgSsnz4hMGyBFlGqHRCvgV6wtAfhc6QZkEMn7/j+FBePZ/isbPJqQwweVkTvr44W54Zj04pIRYNkkomkRUFR06AgglriPhc9DYpdO7IoK1uAx3NaeQc/Iwj5oagzdLUKTAhv5nMqisJhd8LtDIajVgsFnp7ezEajUM+i4NzQ2RZHor2NJlMdHV1sXnzZvp3/Rl/fwP3PqfVnw7D9emHIyuvmBnzl2IymfB7PSQSibTPMYSqsn3zeq656T/YuGbVIUPJsViMmfMWs3ndu6QjFCazhapxNcRjMSLh8GHLqEAwocVk7BrU4jN6IxBOnngDPxQcwG7LxmDzkVUaZtU/nJgt45EkGZ3egCzrkGSZeNiEI6ePhrUuBttkmndvoKtNJPwEzWchFhkCnlsL/X0DhDpfZWBgYMhikCRpyCl60FcxODhIOBwmEAgQiUSw2+1kZGTQ09ODx+PB17UJR+xNHnxZ8yUcT/QGE+OnL2LuOVey+Pyrcboyj7EGidLKGqYuOBe90cJrK5/h0quuO+SIeCyK1WpLu8axNVO4/uZbuOYr38SY5mJMnzSxSID6XW/QuTPFS7/TI6vlJGIRYpEAwcFeUsk4airFYEcjGx830LG7m22rX6arbecxZUH7rDNifBZHIhiB/3kaxs94kdza96I3D2bRslqt9PX1kZGRQWlp6VDmbrPZDEAoFCIYDBIcbMHU83tWbUuwOr1Z38dEIh6jt7MVT38fyZRKOBI+eqH3oSgK0xacyejx08jKyeaVf/+Dyupx1EyZzvbN6wEtdiSRTKSdCGbQ008sniAnvxinO4NI+NTMAxHw9bBr00pcGUXYXT7MVheyogdVRZIV4rEwAW83nr5mQkHPiA/AGg4hFgfYVAc/+/1KfvOrRUTleZhMTlKpFMFgEL1ej9PpxOv1YrfbaW1txWKxDAVhhUIhetp3MrDxu+zc28v/PH3E9JQfGVVNsWfT23j7u1HVJH7vsWWMSSYTtDfuoaisEr1OQVF0PPPEw3zjBz9l9/bNJBKaKRQ/hmUMWhvrePpfD+Bwugj4P8nV146dRDxCX3cdfd0Hpu0fiNCVkESWrDQY0T4LSZJwu92AtqjQ/tY49btXM2uCHbPFQe9ABFnRclqYzWZ8Ph+KouByuXA6naiqSm9PF2tf+i3+nT9jy65OfvUYhA4MSTqdTkpLSykqKiI7O5vc3NyhCFBVVT9SngZVVfEP9uEfPLaFng/S2dJAw54t1O/eSijoR1VVPAP9TJ+7kP27tf75xNrp7Ny6Ka2Ff1OpFJ1tLTQ17Dvgszi+KDIfcmoM89HHRHQ1jsaIibMYjoOBWgUFBQSDQfbv308ymeSF1V7av3YX377+VaZMmcRgeAwUzsWRUUp2djYDAwNYrVb6eztpq19HaP+vSbZu5Ol3tQjL+Pv8FE6nk9mzZ1NZWUl1dTWjRo0ayq7V2dnJww8/zKpVq2hvb/9Q39isg6osmD8Rqou1odXOXti+H/a1Q4v/w2HeR8Jh0XKLji5MsL+thfV74eA8yj07tnL6sgsxWyyEQyG6OtqxO1wM9vXgNMCEDKjJgGzzgdmnFqAA8svBbILdLQn+ZwXHPMP2cOS44PRaLWdnhgO+c4+2YJFTD6cXacOr2z/BNHwCjRE7dOp2uyktLUWSJEKhEHV1dYf80usVmDEG5k6AqWPMZJfMIqNgCs6sCpBkBrr3svGdf/P8m028s5MPTQUHsNvt1NbWsnTpUsaNG0dVVRV5eXm4XK4hv8fKlSu56aab6O3tRSdBngWumQaXnwGZ+bC/D1raYTAEZfkwazxkeKBrDTy5D55ohNVdh49NcFjgiiXw1Qu0JLnbGqE4R2Z0gcobW1V+/ICWTTu/sJhZC5bw1MN/Z+a8RVQZ/cyJbuS0wgMh3b3QGYXFM2HyPFDMQBzqNkOGGcwV8IO/w/88l/7IzgdRZPj8ErjtSm1ezL9eh5c3QmMnLMiD70+B/V74z3chIlwKnyiSJMVHpGVRUlJCdXU1drudhoYG2tvbP9QliCfhnZ3alp8ZZUrFG+S6X0dRtExVO5pgV/ORfRN+v5/Vq1ezZ88eMjMzqaiooLa2lsWLF1NcXExmZiY+n4/s7GxCnl5m5sLyRTBpMtz7NjzxFvR4QVJ0WKwOQkE/Lkucby+Hc2qhZy/cNUObF/LzzVp49MGetyxpv8w/+QL0++Hb98AbWyElGZkyayEFORYWFLzBK78c5P/9AV7d1IrVaqPYLnFZdjcXzxrDMys2csnL2i+5wQgPfBeyR8Ptj4MnoOXdeHsbxKNw3Uz43g0wuxBufwT2H+Oa0FYT/OyLmkVx85/gtS2alVZshXvmw+mFcPd2uGeXEIqTxYizLBwOB/PnzycvL49EIsGqVatoaGg47BCZoihUVFSQSCRoamoadiX1Y0FRFCwWCwUFBRQWFmIwGNi0aRP9vT3MqIZx5fDcmveyXUuSRE5RBXPOvIy6HevZue41VDXJLZfDhXPh4lthUTb8YAq80QG3rIWkDD+4Aq4+Hf77UXjwJQgcCF51uLO5+hv/hdli4fV//y+O4Ov87dsqv34IynMWcWFGF/Vt3fzLeAYP/PMRVLQ4lF/eCFMrtajRD67rYTCacWblUeLo4+4b/NRmwG33wb1rtNiKo+GwwM+u0/KgXnaHliHMoYdLyrVw8d0+HXdsM7K1M0RKDGWeFEZcUJYkSVRXV5OTk0NhYSFr165l3759R3Q0mkwmpk6dyqhRo2hrazskZFxRlKFIznQ5mFGrv7+fxsZGGhoatCxcenDZtVXJPe+bqa03mCgfW8vsMz9HQflY6ravJRTw8s5OqMiHa8+GO56Bf+yFM4rhq1Ng8Vlw+nS49hfw1KoPx3vklVZhNttIdWyjdLCJoiB8+SqweLv5Vd0EfvRCHRVT5rJ98wYMOu1FPmMqnHertgrbofdUZuqCZUxbeB4dvTF+91AzCaPKD66BSwthbws0f3ilgSHsFnjwFijMhOV3QHM3nFkE9y/WpqX/57sSLxnnU1B7JtFImMH+nsNXJjhhjLigLEmS8Hq9dHd38+KLL7J79+6jZtnW6/Xk5ORgMpmGJpMdxOFwUFNTw9y5c8nLyxtKlnMsHBSaaFybfh76wOSuRDxGe+NuutsbiUXCKIoOSZJRVbj1fuj3aiuhFxbAo36oPh/OGwX/ug+27nvPz69IkG2CyY4QE/ffx+fb7+YXuWtYlA/3rYVzfgwZk8LklqpE4gkCfi9uO9zxRbhgjvaL3zNM10JvMFJQVkVe0SiKRlUTS0rc+X+w4HuQrIQXboX/mndwHsh7yBKcOU1bGb21Fy65HXLRcnT8aR78cz/MWwEvd0i4CyopHTOVsVMXoCgjsud8SjDiuiEGgwG9Xk80Gh2KKzgSLpeLL3/5y/j9flauXEl9ff3QPqvVyvTp01m0aBHd3d2sW7eOzZs3f+yuynBY7W70RhNBn4d47OBa1poj9vufh/PnaPNcHngJVr4Gd07TEses7tKmd1c6INcMHSEtLd7qbtjSf2j/v3Y03HP7JBr374acpUwwPUfPINx4N+w7zHwySVYorayhZsYC9m1dw95t64b2Oa2az+SmRdCzE/78OrxUD65suPZMWFAD/3wG1q6DC4phVq6WW+Ovu6HlfesulVRNpHbe2bQ37GLDm8+JmIiTgFhkKA1cLhdXXXUVeXl5PPLII2zfvv2Q/W63m8suu4ypU6eSTCa599572bx58yfeTpNB+7U+aJlIaKnoLizTRKMnrOXJeHA/NB6hW1BdVcSc6iDF5ZXs3LyOlzZoyw68nw+mJlR0evQGI9Fw6EMvsgRMq4arTofL5oHNAEYJpFbo2AlxnzYr9vEG+L86aAsOE/UgSZgtdmLRMMmjJOMRnBiEWKRBdnY2N9xwA4qi8Oyzzw4rBLm5uVx11VXMnTsXSZK4+eabaW39dCZ4NVus2J1O/F4v4dCRl1U8VixGyLBAsRnMaLEkW/uhNwxRYSyc0kiSFB9RPouPgslkIhKJHLHL0t3dzdNPP01lZSWzZ8/mnHPOGUro+2kjHAoy2N9/3IUCNKunzQPvdmjZtJ5r0SwJIRSfDkbUaMhHwel0UlxczODgIFu2bDnsIsZ+/3u2/aZNm446ynIq82ltt+DEIUlSSnRDjoKiKJSXl5ORkcG2bduGzbZ1EIPBQFFREdFolPb29k+wlceHjKwcCoqK6e/tobP909mNEpwYhM8iTSRJQpKkEzLKcSpROqoSz0Affq82RipyOQgOInwWaXIwue5nndamekpHjcZqt7Ng6dmYzGbyi0owmswUl43CZLYgywoWq5aUWG8wYLFaycrJBaC4bBR6vfjd+awiIlwEAJSUj6alsQ5FUZAlmZaGesZMmEQ0EiEjMwuzxYrFaiM7N5+Bvh56ujrJKyyiqKScSDhEU/1+3BmZ9PV0E49/7LTcglMQYVkIAHAcSOQDEtl5+bS3NGE0mdm9fQuZ2bns2rZJG1Z1aEmBJk2bSXtLE6lUkt7uLswWCyaL5YSMoghODcRoiAAAi81OYXEpgwP9RMJhHC43/b09BAN+jCYzqVQKp8tNY91eJEki4PPiHfTQ1tJEMpnAZLFSVlFJ/b7daSXNEXy6EKMhguOCoijU1M4gEg6xZ8fWk90cwQlAODgFxwWT2YI7I5POtpaT3RTBCURYFgKB4KgIy0IgEKSNEAvBKUFmds5h84HIskLl2PHD7ps5fzFWmx2A6XMXYLM7DtlfUj6ahUvPRm8Y3nguHTUanV7/MVo+chBiITjpWKxWrv/6dzBbrEOf2Z2uof+7MjLwe7U1SST50EdWlmXyC4uRZJkx4ycRi72XPUhRdLjcGTTs3zu0FsoHyztdGSSOkADpg8ePZMTQqeCkE4/H2bphLYlEHHdGFjqdDovFSjwWo7i8ArvDhaqqJBIJ5i05k9amhqGI2py8ApAkMrNyCAYDtDU3YrHacLrcFJaUkptfSP2+3ZRXVqOmksxasJjm+v0UFJUQjUYoKhtFMpHA7nCiNxgwmcw43Rnavy43sxcsob2liYLCEpA4EIQWJhGPYzSZSKaRQOmzgCRJKSEWglOCWCxKSXkFBUUl2OxODCYjeYVFtDbWM2HKNHR6AwG/l1QqRU+XtkCJ052BougwWywYjSZikQgDfb1MnDqTqnET8PT3sWXDGirHTMBssdLf20PA78NisTJx6gx0Oh25+YXo9QbMZgsdrS2Uja7C4XJRUFRKLBolGNBmE1eNm0A0EqGguASjyUR2Xj6yrOD3ndqrsB0vRlwOTsGpTUFhCc2NdYRDQeKxGIqsEAoGCQX8BHxezGYr3Z3vzeYtKimjtameSDjMzq0bQYIxNZNIpZJ0tbehqirujEx6utqJRMLkFRbS3dFOUdkoLFYbne2ttDU3EotG8Qz0MWbCRMKhIHq9gVg8Rn9fDwP9vWTn5fPuW6+RV1DIzi0bAagaO4GuETYzV1gWglOGUFBbmT4SDiOBZuYnEwz09ZKIx/H7BsnMzsXT3wdoyY4DPi99Pd0kEomhWbKdbS0YDEYKi0sJBgN4PQM4nC4G+vpwOJ2YzGa2b15PJBwiN7+IPTu2UDqqkuaGOmYtWELj/j3o9QYG+vvIzsmjp7MDv2+QVCqF2WpDliTaW5sYHPhoS0h+GhERnILPLFXjaqjfu+uYEvlUj6vB4XKzfvVbJ7Bln05EnIXgM8tHWXjaYDIR8PuOfuAIRZJlOZJKpYwnuyECwXFFko68tqTgmJBlOSpLkvTZz+oiGHkIoTiuiNEQgUCQNkIsBAJBWgixEAgEaSHEQiAQpIUQC4FAkBZCLAQCQVoIsRAIBGkhxEIgEKSFEAuBQJAWQiwEAkFaCLEQCARpIcRCIBCkhRALgUCQFjpJkuoURRl9shsiEAhOXSRJqv//TQYyChKGA5sAAAAASUVORK5CYII="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydCcBNVdfH9Zb0Nr/NyZh5zEyGIg0KDUoTpUGSoURJEUJUpEgZQwgpkjQqQxSZ5zkkDSqNGtDwrd91t++6zrnD4xnuvc//ZHfvc88+++z9O+fss/dae62VI4c2ERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABEchiAkdk8fl1ehEQAREQAREQAREQAREQAREQAREQARHINgSOsO2EE086mXTcCSeeeOxxxx2f65j//jdnzpxHH3VUzpz/sY08+/bt3bvru293rlu9Yuk/f//9d7YBpIaKgAiIgAhkawJSWGTry6/Gi4AIiEDiEch/buGiufPkK3DkUUcdtfPrr3Z8tnHdGk3QEu86qUYiIAKZR6DtQ91679796y+jnu//ROadVWdKbwJ58hcstPOrL79AAJneZas8ERCBxCNQsVrNCx/q8dTAd954bcKeP//4o0iJ0mXzFSxUJPc5+fKfduaZZ6OYiLXWg5/u3W3Ys0/0iDV/RuRDidJ/xISpfN57W+MGGXEOlSkCIiACIiACEJDCQveBCIiACIhAQhCofmHdyzp069P/3CLFS4ZW6Kcfdn0/cfSwQQjq9u7dsychKqtKiIAIiEAmEahS48KLhk5880P6v1ol8568d8+ff2bSqXWadCRQvvL5NUdOeW/u0oWfzL3z2noXpGPRKkoERCABCRyd65hjBox6ZVq1WnUuiVQ902P8/vtvu3db1/4H/fxff+3b949t/1pyx7Gv18PtWm5cu2pFVja1RJlyFce//dHiX37+6ccLS+c7JSvronOLgAiIgAikNoGjUrt5ap0IiIAIiEAyEKjf6IamvQYMH0tdv/lqxxdrli9ZyGStcLGSpQsWKVaiZfuHu9eqe1n9Vk2uvoxJUjK0SXUUAREQgfQgUNP6PsrZvH7tKikr0oNo1pRRvc7F9TjzGWflPidraqCzioAIZCaBJ18YNdEpK77/9puvF8+fN3v96hXLPt+yeaONdbd/t/Obr3/+8YddKCgys16Hc64KVavX4vivd2z//HDK0bEiIAIiIAIiEI2AFBbRCGm/CIiACIhAhhI465w8+bo+9dxwTvJMry4Pjhs+qD/KCndSzOl7PTtsTKnzKlR+fOCIcW2bXRcQ3mkTAREQgexAAOsz2rl4/tzZ2aG9qdrGIsVLlaFtG0xgmaptVLtEQAT+nwDxKPjrX9uuq1u1tK23+SHZ+ZQpX6kqbdi8Yd3qZG+L6i8CIiACIpDYBP6T2NVT7URABERABFKdwF33duyC2fyrY0cMHjN0YL9QZQVtX7Jg3pzbr7201q7vv91Z86JLr7ioXsNrUp2J2icCIiACECCmT6GiJUrxfdWyxZ+KSvISwHc9tV+zYumi5G2Fai4CIhArgcnjRg4l74Y1K5engrKCtpQ6r2JlPrPaNVWs10D5REAEREAEkpeAFBbJe+1UcxEQARFIegJHH50r16UNG13P6rORg/r38WvQN1/u2P70Yw+3Z3+zlvc9mPQNVwNEQAREIAYC9a+98RaXDTciMRyiLAlI4PgTTjwpd558BaiaFBYJeIFUJRHIAAJlKlSuRrFLP/3kowwoPtOLPOnk/52SJ3/BQpx43arlSzK9AjqhCIiACIhAtiIghUW2utxqrAiIgAgkFoFipcqUQ5AT9Of7RaTavT/99UkE4C5bscr55+TNXzCxWqLaiIAIiED6EjjCtvqNbmzqSv1y+9Yt6XsGlZZZBIqVKluOc6GcN4XF4sw6r84jAiKQdQQYr3L2pQs/mZt1tUi/MxcvU66C68dMYbE0/UpWSSIgAiIgAiJwKAEpLHRXiIAIiIAIZBmBc4sUL8nJd1nkwWiV+Puvv/6a/9HM9//5+++/Tzjp5JOj5dd+ERABEUhmAtVrX1zPrcr/bfevv/z+22+7k7k92bnuxUuXLU/7t2/9bBPXMjuzUNtFIDsQOPKoo44qWaZcRdq6fNGCj1Ohza499GPWjf2cCm1SG0RABERABBKXgBQWiXttVDMREAERSHkCJ5p9OY10gQmjNfiJLh3aXFu3Sqn1CloaDZX2i4AIJDmBJs1bt3NN+OarHREt0JK8qSlf/RKl969MXrtymawrUv5qq4EikCNH0RKlz2Ns+9WO7dtiWZSTDMyKlz4v0I+tXr5kYTLUV3UUAREQARFIbgJHJXf1VXsREAEREIFkJvCXmU1Qf/MKFZPFxC8WtZCUzG1W3UVABEQgGgGsz86/4KJLXb6vd3zxebRjtD9xCRQvs1/Qt27lMvl9T9zLpJr5EFj2xQGjoJyW5W9L/5C1fN4TxcyHQNkKVQLxK1YtXbggVSCVLFs+YDGyetmiT1OlTWqHCIiACIhA4hKQwiJxr41qJgIiIAIpT+CrL7Zvo5G58+YrcNRROXP+9de+fSnfaDUwSwiYwOUcOzHClm9NyPJ7llRCJxWBGAk0u+e+B8m6588//mCV7tdfbpfCIkZ2iZbNLt+xBQsVLU691ipQbaJdHtUndgK8P4ta+q+lZZZQXGjzIeACbqeKNQIW0S7g9qpli6Ww0J0vAiIgAiKQ4QTkEirDEesEIiAC2ZEAq9EsHWPp6OzY/ljbbEH7AqtNc+Y8+uiCRYqViPU45ROBWAkEn8UjLX8ZS2UtlbTffMc/wfw8v/8J+R7r6ZRPBA6bQN4C5xZu0OjGW4h1sGDurBkU6JS7h124Csh0AuZGpfx/jjzySAJur1+tQLWZfgF0wvQicIQVRCpt6dT0KjRVyylboXLAwiJVFBZmXVGJ9uzdu2fPxrWrV6TqdVO7REAEREAEEoeAFBaJcy1UExEQgRQhEDSdp389y1J5+/uEFGlaujfj22+++pLgfRRcsVqNC9P9BCpQBPYTQHHIc4iQhVWi0bbjLQPxVXJFy6j9IpDeBO66t2MXBNwTRg15zhbnH0f5+EFP7/OovMwhUCIYeHfb5o3rf9u9+9f0OutJ/zvl1NPPPDt3tPKOsC1aHu3PXgRsXJorDQtqUPxzLzG+PTZ7EYuvtTybKJ7N6+lf61atWBrf0YmZu0zQxRXKin379u5NzFpmTK2Ci1eOCF3EEuImLWNOqlJFQAREQAQCAw5tIiACIiAC6U+ASd0plgpZCgictHkTmDfz/bfZU6P2JfXESAQyiEBBKxdlxbeW1phLqID/7fAtZAKKYIY8/2ZQfVSsCHgSyFewUJH6jW5oinXFuGGD+p+ZO09eMn71xefbhCw5CZQqWyGwMnnV8vRzo3LhJVdcOWPJxq+mf7JyS7VadS7xInPaGWedPeyV6TMXbvl+z7VNbm+RnPRU6/QmELQwPMnKjXdsyrgWN1DrLO1O73qlUnnOuuKzjevW4NYvFdpWvsr5NWlHqliMxHlNuPfPtuRci8Z5uLKLgAiIgAikhYAUFmmhpmNEQAREIDqBYywLgiZWdseyojt6iSma48N3pk2haVVqXlj3eIu+naLNVLOygECItRORQX+wtNZStPgVzu0F1hUaJ2XBdcvOp2z94KO9nHXFzz/9+ANCZ3h8/eWO7dmZSzK3vdR5FSpT//T0+97ukR5P4krx6KNz5brPvnvx6T/85SmVq19Qh/hQlavXqpPMDFX3dCXAew1lxfGR3CN6nJH3KHHGTrckq50IlyTV4lf8xzanhFmzYsmidL0bk6Mw4r6WtHSeJazntYmACIiACGQCAU3EMwGyTiECIpAtCbBCe7Ml/LxmK9PpeK/28kXz5+EaCsHLxVdcdW28xyu/CEQhgOIBoW8eS0Us8WxG2nB1gWCG51bPrm6vTCOA66BLGlzTGLdBWFcQbPu4448/AZ/hP3z/7c60VAQl8Jlnn8O9ry0LCHD98p1bmEDFOVanY6Da3HnzFXDN2fn1l1+EN417xwlN2bd4/rzZWdB8nTIxCSB8ZXEIbhLjUTzwbsRVIkG34zkuMSlkYK3KlK9cleLXrFiaEsL9wsVLlTnOXia0ae2KZYszEF2iFo3FrbO6lavQRL1KqpcIiEDKEZDCIuUuqRokAiKQIAQwAWdFN5un+5kEqWeWV+Mf295+fdLLVKTh9U1uy/IKqQKpRoBJNooKVsWxMhSXFpE2F7uCfIFn11xIpRoTtScBCbBqnngDL48Y9AzWFaecdtoZVNN0FV8TsDneKrMC/+W35iwaPumtWfEeq/zpQ6B46XIVWJ1sXmF+37R+zar0KdWUH0FB6OYNa1f37HjvIe6e9u75889N61av5Hyfzp31wesTx7yYXudWOUlPAKU97zeUDvH0Kz9b/m8s/eTejUlPIgMaQB/urKpSxX3SeRWrVgfVH7///tu2zzauzwBsiV4kzwqW87iEksIi0a+W6icCIpAyBKSwSJlLqYaIgAgkGAFWotW1dJElAvhqi0Bg2qSXR7O7QpXqtQoXK1lasEQgnQgwyeT5w9JptaUvLXkqLILuo1x+3GUwOdUmAplCoHrti+tVqVm77i7TTrw0ZEBfTnry/049jc9d36XNuqL2ZfWvIibG99/tRMioLQsIOMHl2lXLlhCAN72q0OPBNs2f7Prgvc2uqns+90x4uSi4brmybrWbr7igUqtbGtVLz3OnVxtUTpYRwHIQ14i4LI3VUgIlRylL9S3lt4RrKG0eBPIXKlLMDNtORriPQjEVIJWrXK0G7diwZuVyFhmlQpvS0IZf7RgWEZyZhmN1iAiIgAiIQBoISGGRBmg6RAREQARiIIDCglU4WFr8FkP+bJ1l6+YN65aZaygg3NDsrtbZGoYany4EQhQQxazACyyhqNhg1hKRVpQilMF9FMdoUpouV0KFRCPACnysK8g35One3X7/7bdAQNsTTjr5ZD5/+P47gsXHvRGYmYNWLlk4P+6DdUC6EDiw0jod3UFRsc+3bN44cdTQ59y94lVZgv2uW7V8yT9//x3Nqixd2qpCkobAKVbTfHHWFplBNUu4l+N+kgzBB2DZ8pXhlGPtyqWLU+XZO6/SfguLDWtXLo/zvkmV7Cj2UDgzRsSlmjYREAEREIFMIKDBRiZA1ilEQASyJQEUFqxAYwWb+toYboHXxr44hGxXNLqxKX6/YzhEWUQgGgGeP5QPBSyxqvT7KAfg1zuvJZQW0YJzRzu39otATAQaXndzsyIlSpfdumnDuikTXhrhDjrBlunyffcvP+OCJe7NCZmksIgbXbodUKpcxUDA7ZVLFy1It0JVkAgcHgHGVyyo2WEK/HiUWSy+mW1pjaV0sxY6vKYk3tFlylcKxK9YsfjTTxKvdvHX6LQzzjr7nLz5C3Lk5vVr082tXfw1ydIjsLjFQnetJY0Ns/RS6OQiIALZiYA0xNnpaqutIiACmUmAoIS482CQi9BJLjmi0J8xfeqrHbr26X/Kaaef0eDam2995aVhz2fmBdO5UpIAz+FGS7kt4Roqmr9u4ld8ZgnTf5I2EchQAhYb+dhWD3bpyUkG9On6UOiK3P8ed1zAneDu3b/8Em8ljrVjnZBp7cpsGSQ1XmTpnv/kU049zV2DNcuXLEz3E6hAEYiTgFkeOhdQWHEdzd9RrA7dGXh3/mkJl53bLWXHOAYx0S5VrlIVMjqXfOYZavfePXv2mEe4ff+aO6XQeETEuzjCLOyOPPI/Rx51VM6ciz75aNY7U18dH9OJLFOFqjUuKF66bPnxLw4eEH4Mbqns3/++/mrH9ngsPXgnHWnbb7t3B8ZATvHN943BuDix1O/U0888q2K1GhdQB9qFVVgsxyVoHsaSuET7wpKUdQl6kVQtERCB1CMghUXqXVO1SAREIDEIMLljFRsD9DS580iMZmReLfbt27v3dVtdfGfbBx65vlnzVumhsLAZ4FFM2n6xALap6nf33CLFS5Y8r3wl5r0fffDu9J9//GFX5l21hD/TqVbDwpZwf/GDpUgKCwQ5+CdmYkpw0T0J3zpVMOkJ3Hr3fQ+ccVbucxbPnzt7zox33gxtEEGz+Xvv3r1x34sFChUtTp+AO6lvvtqBkCXmLW+Bcwtf1/SOu0cOeroPwb/DD6TcwsVLlTF5VO4tm9av/ebLHQgwD9nIV7ZilfNPPe2MMxd+PGfm7l9/4bmKe8tlErRcuXIdY4YmP8Z6cI06l1xe57IGV5/8v1NO/earL7+YPnnCmPWrVyyLdvxd9z306GVXNrrh4dZ33BQeJPusc/Lkoy07TQL4/bfffB2trNLlKgYEl+SN9xpEK9tv/3+PPfa4v//+52+Cbsdaxtl58ua/6vqmt48dNqj/b3aRQo87Otcxx7DA2sKgfIWLqWhlcq2q1LjgojPPPifPFrMYWvrpxx9FO0b7M5UA7zksgHF5iED6qzjOzvuURTgcg8WitjAC3P9FS5Qqy8+MzUjxQDrF+pdYFRaMbweOnvTmccefcOLMd96c4voYnueHevQdWKtuvQa4G7TH9vcX+vXqOnbYc0/71SX/uYWLNr2rTfuL6jW8hkVD5Ftlbuw639u8ablK++NXMIbevH5NVAsLlOX3d+7V95qbmjWnjhxrupp9He5q0ogxajw8EigvrqCKWGIsKReLCXRhVBUREIHUJiCFRWpfX7VOBEQgawgwIcRk2FlVxCw4yJrqJs5ZX3t55NDbW93/EJO8ytUvqMOqrHhrh5CswXU33dq46Z0tzR1HFSZsCLomjBw8cNizT/aIpLhgRdjQidM++OmHXd+3ufXaK5joufOz+q1l+4e7X33jLXfYSrm/Rr/wzJMTRw8bFKl+1OWZFydMRXjIZO2zjetwpXBgu+Ka65u0aNepKxPE96ZNfuWprh3vRXETS5tZudv1qeeGE6jX5d9lUqWmDetU9RMgxlJuiuVhgonPbVxBESgyWoBRJqNFLSHgDayIttWnKYZEzUkUAqefeXbu2+5p15E+6ekej7QPrxd9Dr/FEjC5SfNW7Vo/2LUXgqE/LLABfQ/HIrCfvXLbAVdoFs7gb5SaA/p06zRnxtvTvFg8+uTAYfS/5q58yXvTXpsYmqfuFVdd265zz6fy5CtwLr+zcrdv94fahfeFl1/d+Gb6tgIWgJZ89EnNrr64umlPcKsRdUPwfkuLezs0tL48T/6ChThgx/ZtW559/NGOH779xmS/Amh3t37Pv4gAPjTPzXfecx999sAnuj8c6eQt7+/UzZY7H1mtVp1LnMKCPvb+zj37Fi99Xnl37Kz3pk9FmEdgXb/ynMJitYd1BfFFbrz97jYFCxctARsTKD6KUicqGJ8MrLRu3fHRXk64+OrYEYOf6PJAm1jK69z72cEoeL74fOtnb02eOJZjELy2fahb72ub3N6CFdesCn97yivjejx0bwsvZQjcb7itRZvWDz7a0+SnAVdmbCi9nnvysUdiqYfyZAoBXJSeYwnXh1GVbiE1QtmPsoJjGaMEgm4TK0rvyP+nVKLMeRUQ0tPPDR/wVE/7mpO/6cvtX04+jzyKX/b/zf94tswIYzf9W3h/G+mOwFETygry0OfzWbRkmfOGTpj2AdZd7lie35btH+nup7Cwfqjt/V169T366Fy5UFhuMisKFBi4tnrupdfecmVv+2zj+kgxczifGVOcMsTOT1/Je2uVucI7x94VjHHv7/J4v7kfvvdWqIVJptzx6XMS5nE8L8R/ya5Bx9OHpEoRAREQAREQAREQARHIOgKY2FuqaekBSzdaOjB5z7paJc+ZB45+dbox+7ffsHG+Qim/1jBZGj7prVkc79LS7T//476jcIhEAqGWyxtqBo8A69mRE98ILZfvocoCr3KZPLpjsBwJzdOs5X0PhpfnXMNEu1pMiues3v4Dx89b9+XPo6a8P2/Bpp2/8zfCxmjHp/p+hCiW/mOpsqWnLfW2dF2IO4xDENi+Iy01sNTBUiVLOYOBu1Mdl9qXRQR69B8yOtIze0OzFq3Z3/7Rx/tFq+LQiW9+SN7FW3/YR5/w6eZv/wjvX9zfi7bu2nvZldfd6Fcmx5O3+oV1LwvNc+/Djz3hVSblYZVBXtx/uD6cvvedBWs/d33wI737vxCtHewvVqpsubfnr9nm1Ycv+fynv6vUuPAiv3JQVLjjxr4569Nezw4b896i9Tvcbyhc/I5FSO/yVa99cT3y3dKibQdXf849Y8nGr1weFDeR2oOwj7yhfT+CSuoUzpHrla9gIRSscW0oClo90LlH6HvOlV24WEnc90TduEYcU/fyKxuRGavEcdNnL/S61iXKlKsYXiCLAh7rP3iUyz9pxvyVU+cs3eDuR1Z8R62EMmQKAbsm3OPXWrrV0gEFXLST8+601NgSfcDDlk7j/ah35MHkmt7V+n7uexaTRGN6uPvrX3vjLZyLZ42yChYuVgLlNL9N/2TVFqwlUDrc3rp9J7+xKm5Yyb9wy/d7UFw4JTnK9Glzl28K7QN4xiPVmWNHvz7jY46h/y5iVnjkR1nhxqdO+Xy4bc/s461Nx1liPHm+pQK69zP7Cuh8IiAC2ZWALCyy65VXu0VABDKawOl2AlaWsiINP+RpcoWR0ZVMxPJxC1Wr7mX161xa/yrcSuz8+ssdsdQTZcWLk9/9qJDZ42MZMezZJ3pMGT96OH54mUTe90iPJ5u1bPcgq8ycb97wcnFfwm9YObDKzO2/p8Mjj7EiltXLmMmzihVB0ZWNm9y2cN7sD/3q58pj/9oVSxe7fOdfcNGl1Ie/WX3LRJNA45T3Qt9ej0ZqL25JBr/8xvsIBhfMnTWjU+vbb2LF9IWXXN7w2ZGvTGOlbCy8skEeVqfjyoC4FKwIXR7FVzduMliVSBBSXPCwiu4om5gyVsIdAEFK+c7vuEbBjzF/88mqVVa0c05WorL6lHLYz+/OpQ9/k9flcSv1yMNvviv3tIo1te5YVt9jCYabpEFP9ejs1TpnDeZcQ0Ui0PbW665AMMTKXo5DgYFgv5O5NsItDxYLCJT+tmWvuCjy6wPpc92q3R/Nn5Q7JwpWrN/4+7VxI4diEVDqvAqVEcpT7qUNG10/bdLLowePn/o+ffDHs2a8g+UFfssRdNG34UYq2lWEi63QnSHjOH0AACAASURBVEEdzPX6NiwqcCPCkuTHnn5hJAqHltYf+1kjoHTmHG+/PullLCD4Tl/5wstT36O+Bc3aza8ORUuWPo999P+LPv5oJtYFTlk0/6OZ7/d+uN09rIJGicHvWJFQP6/yeD+UqVC5GvuchQWK737Dxr7Gu4Rz8H7avvWzTax+Rklwi7lkefyR+++Jxsjtp7zH+r0wkvuI33hXTps0blTNi+rVR6ldrsr5NfnNbjHfoO1n5c6Tl3cKxxMYnNXY8C9ZtnwlrEde6NfTLD8+mnlexarV/zFzmnWrli8Jrx+KLK4vlhdd77/ntvfenPwKSowx02YugHnVmnUunjpxzIuxtCsoAGfcRH94wBWa+r9Y6MWUB66MT3nXEMfCcwtTRPDO4v3HKn6UarzfsHrinfmL5cV1He87xrq4QqVsrFNdYr97X/KOpQ7s4/ryN67eOJby2HiP8s7dZoljuR+oK7/zDuU79zTndHmpE+d171fO4VxA/ptZ94+zqjoca6kgg6gf59e66BIyfTL7g3dxw9R/+MtTTjKLOiyTH2jR9FrnQo8xq1dhWOUxNsZKrt0dN15FOS7fd+b3Diu8fkPHvuZ+ixZEvM1DXR9noc+Pu77/rnnjy2vTf3Msbgm/+mL7toJFipU4wxQhO8ySK2rjEi8Dz8wVlnC5+lbiVU81EgEREIHUJCCFRWpeV7VKBEQg6wkwAWNyV8BSwK2HttgIYDKOAJ6J12VXXnvjmKEDo64uxsAeiwwEZUy07rn56ktD3S+9NGRAXyZmuHyqUqN2Xdx5eNWmVNkKlfgdYZUzfUfpcEfrDg8jYGrbrHH9T+fO+qDLEwOGIswqVqpMuUitKmVCH/YjlFw8f95sviOY6vHMkNEItAY/3bsbipV6V113U59BI8cjLKTdfnEoEAI99cJLr5Bn+aIFH9/brHED50LKTUpPN4fjsZFO+VzHWQtZ2bvVEj72Pf3sh1DAbzN+vXGVgdsa/Hs3sARPhCoIanDzRj5c7DCBrWBpgSX8viOQ4e91lrjW2yxdaamyJVyBrbDEuAt3U5wHYc1OS5stYYVFPlwOEPOGfdQBRQbKkT0mFEIgw++4JnCKjQMxOTJLIGPn1naYBHj2O5qP8f19wOPdEPB4FYmAmN9d8O1Ip7UwF3ucD3PKNUFxoO9ZsWTBJ/SJsVbZ5PkEFg1sP+7aFagXfeC9nbr34fvwAU/2fKHf4135jrsPl9e8+JV5ftyUd+mDUcDgCsi5/nAuraK5tqL/w5INZcWSBfPmtG9+8zVO6GY3/h/PmzIXhQXCcxTU4fE1ENoVKVE64D/+rSkTx7m6Ucb9d950NdYXUyaM9l35XLzUfpdPn21Yt+bcosVLPtSz73P8Pf21CWO6dbjndqdAsrLHorAg9giKZi/lD9YS1BEGFnB7EeVgkYGygvq0bXZd/ZVLFgZ8oTvXYBUsQG2s14lrjIVO/UY3BJQy+L1//OH7WlIXXDuxr3PvZwajBLnqgvK4ufPccH3FDhT03Ce9Bgwfi7ICN1X33ta4gXOLtXHtKvqvQ7aaF116Bcos2HS8p9n1Lg4Lf69duXQxCgvaF2u7LB99JO9V+m6E2ixY2GL9H/1xqBD6oCLV/8VMGL70B7yreNdt8jmSdw/v0AKWePdxHMo+rHZOtoRrqJqWeD+hPHDjDq4ZcaDcuwtFFWNg3qHh1k1D7TfuXxQVXu4aGUOjsODd97ollBoFLSE05v3IvYGyjXcx7kNx41grWM9P7JN3K4sVsNbiveqUGryrUWKku2uf0uUrV7WycyxZ8PEcPjNyq2yxYih/3sz33m7/aO+nCxQuWnzpwk/mMk6NFm8GizjXpw8z11WhygpX57mmKOY5ZtzJb4w5/dqDNTF9DftRFDtlhcvv3mEEIM9IJhlYNvc/9xr3oOZ0GQhaRYuACIhAKAEpLHQ/iIAIiED6E2DihVCRCRoDW1zTsDqNxEQJIRQTbz6ZMDmho5uweQYGTsYJOS5NChYpWuLJRx9sG6vfWqwYZrw19TWCvrJqNxaFxR2t2neqdH6t2igZwpUVXF7ObTKcTSgsEKh5KSxQJDhzdbcfn77d+z7/IhO2/j27PoSygvLWrFi6CIUF/uEj3T7OfcbHs95/xykWOnTr0/80UyrMfv+tN1BWuPJcOZTpp7C4/tbmrVi1i6DugbtvuS403oUtoGYilcOMS3x9qqf/rZ7QJSJIIeg9PPwEIqENINYFyginnODZRFCDlQYrr/3GTAHXMSEbQp1rwn5DiHpT8Le59olQJXTbZn8U8KCJYgThEArQkZZWWyJwML8jJMJ6hDr/an0Mygz8WdP3oAgJCGUsudgdAeFMFCsTjyqkz08+rkPo81xyfKkzq2uddQp/I3RilS2/IXQK7Ue5tgjWXOwXngOEZvS3lIOgk3shvF8lP4IY1wc7YWiG978IznHVgVL1lZeGP+9H2HSkgTaZTDyuQCrEzEHov+v7b3fGG8+G/pFzIvD61gTYWE/gZo7V/B++M22KU1aQ50TrrFzdL2147Q0I0bE4QEEc2ibnLsoMOyLGrzALilH00QjJ77v9+obhioDPt27eSF9Of8xq3XABGopcF7vjz7DYEgjjRzzX9/FId3PJsvvdHW1ct3oFdcGyBSu2bg+0uiM09hEKJlYlw+S/xx5/vJfCwllXfP7Zpg0orLF8Q6CHFQLxkUKVPaw+5rzxCPaJL+GUFbwjn+nV5UHXtv+ZqY377mdJ4/ZXDrrXmjfz/bdRnFMm902LGxvU/WLbFgS+vhvWGMS/IMOo5/s/ER40/lhjw74/ft8dj5CS5xHhMiv1uR4kFMUIpOn3UO7yyTNN3tAxVKTqHta+KP2XK9v1Hc7iDmE7fRD9Ff0W/RfCfMZ+7CMf+0jOeoDvtM0JRTmOfCT6A8qjv3P5XH8JB5fXMTkQtylEOM87A+UC5UUav7CfPhdlE/m5hhxL4v4KBGYOtoc2uc1ZSbh9keKo3B1ynNdX2skGiyZR8qJ4m2GJY6pbusESixQYA0yxhHIV5lh58X7AVehs++Reoq2wO6Tvj2fcTdwIYothhRWPkjhKuzx306eiMMWamD6x0c233YV1HZYV0ZQVFIgrqKNzHXMM74dRFtvH6yQowYlpwdiYMenWzRtYjOG5te/Sqx/94Zuvjn8Ja7TQTPTLWHLRZ36+ZRPX45At+HwxFuBe4r7jevA397CzePV9R8dznSKcn13O2jU8G2MwFGRYSmuMnZabVseIgAiIQBoISGGRBmg6RAREQARiIMDECDdQTNgRnDHoxoQe4ScDXvYxIGelNZ9M0EsG87FamwE6v7OSLOBqxgb0CCLZx2SXCRbnYALLIN65pnH73OQrsDIqmMdV202m+ZvJL5sz16euzl0Nk0Rn6s8Ej7KdEDRqoEVcHhFQFuHOU90euu9fm6y4CkT7/ODtNwIKC7c6M9Lkj5Wsd7XrGHCjhAuS8MDW7lwmM0FwmYPJk9f5QwOqIrwhz6133/sAgrFli+bPG//i4AHuuH9NesV3Atj6tQVhV6Fi+4V/c4PllatcrQbCSlbY9rTgpeHlRSqTlbwtO3R+jDz9ezzSgQDboefG7zt/b9m4fm00vtlkP9eZ1Zjc76wUd8/CIc23Z4t9CGKYiHJtnZuJLfYdYY0T2qQHugIehfgJpF3gTAREuOOh3yBv+GpU7u0JlnBBg3JkvCUUGzy3TrlBWypYWxEEco8gPKZPoa9wLq+YlPP8u/KdcjVcqO+UDKH9S6hihDJc/0HZ1BmBF8ch6II1G64h6FNwn4e7BfbR56E8gjv3OH0eQg4UQdQVtxXUk74U4RjXDOsUykEoRTBozs0x7lr+YN9ZHUp/yQpY7g3aj2CE830eLIf9bkWvc1liP6XfhnsiXOhQIorcSFYHe/bs4fr49ll+tUIZwr7VPq5AIrWmUPH9cQ9Ml7ISAdNNze9uSywE3Ej1eLBN89BjTTYXCIbNhqJg2qsvjw5XVrDPKYK3bPLvm3BrVLVWnYsRkj1sbqy8BO3Ux+T9fyAoP8mkg+HtCFX0nm7CvHivmlMwFzfTOFYMf2mmCh1b3no95w0v64jgqmOvANTkLRviDoog1N0tEDi/9+ncoXWosoLfjrLIu3yacDDwjoq2oVTALz35CHYeqqzgt3pXNXbKUXMXM+OAmxevcitWq3Ehv2Ohh9992tqxZbProykrOKZp8zb3404Kt19Dn3ki8G4K3YoGLRDjfCc5ASV9C4J7+gT6DxjRjxewRF/C4gHuAcZO/wsKPOkvYEgZbmxEn+PGOVxHvjvhvlOKupX3Li/jIPoW8tI/cG76JPZjneCEquynr0Nxh3UMfQcWfc4NIApvBOnUiRX/dS2VsEQfTN/DOI8+kP4J5RAuKTnfq5aICUNfjmKavsrFI6Gu9JVY53BP8QzynnDKEPpD3FTSd9BPIsDH//5S+2Sjr73UEm360X7nOXEKEsrmuL0mAP7L9lEv3hVu/IpVhuu7g8Ud+HjTvjUM/9H+dsw9duVYbj9GtFL1Osh+o41OmRGaBdZOOUabYI51I+8E3hfOBRXXjfchrPmN/ass0V7uO64xx8e1OXdQKyJYIsRVYITMjCXZvWbFkkUPdH/iGfrfxx5ofaeftV5oUYyrcSHKb8+byze/PowFO849IGNgv0VHvG9c342rwPBqN7BYG/yG9Qdu5mJgwPPB/ckzgoKS54dnkmvOd54vxgU8bzwf3KturkL53Mf0GW4/5QQWj1lyi1foK3jHM7ZzzzHn4NwcTznuuzuWe5nFK9w7X2XV4o8Y+CmLCIiACKQMASksUuZSqiEiIAIJRoBJNCupq1hyE0kmQJgUIyDAvQIuO5jAotRg8HyWRxsQUDJZZDKLANKtGuZ3Bu0M1hlUF7A02xIDasphYv+RJQR5TMYYfPMbg3wG/AzgCdTHQB13ERznVjQxAXf+gZn0M1nmePfOIF/EDWEKyoqfftj1/T1Nrr7US+ATqYDF8+fOZlUqgp7K1WvVwR+5X/57TIiPcgA/4W+8MpZV6J6bUy6Y9yjPd59z74SgBtcqnPvWlvc+gEDx8U7tWoZO1v536v4VrJF8g6OscAEMcTFF/lYPdOnJ53NPdH8Yv76uoq68SGVef+tdrXAxsnnD2tXTJ08YE95I58f84xA/xF4gbGLnhDIHCeFSZfIVslKPlZQFLCG8RygU6b7lnuceR2CxydI0S6ymY4L7niUmv+xjAozABqEPzxbPJhNehOPkRWjF8TzTKKtGW5ptiRWf7EewhfUDzzHPNArL6yzxLNIvUG6kjcm710YfEHr8zfY3KdKGoIbnn34BwR9te8USdUdgUyC4D2E+7WO1KsIszsWx9G0IhxD64L6FPg3hE9xwgUMAX9x90B9RNooT+p6Ay57g5ly+IJTEkoR7knJwm0VZbqX4CPtOf0m/hXAOlgjPeJZxA8L1ow2UQX0RFFIP2oeg0Sl4qS/XgHw8f9SLc28L5qVtlEn/yjFOEWxf02dDWcHzjgsffI1HKvXPP34LCHdYuRvP2fEjTv5oPse9ynQWFhtWr1iGi6U72zzwCPme7NrxXueeyR1HjAT3HWVE70fatwovE4sJVtfyu59LEfrvVh269CDPhJFDBvopndkfqR/Hwm7b5o3rcY1Szhi8N+21ibFyow64gSI/ygr6+27t77ndq48nHsgBSw5b4ex1jtLl9ruGQRFAjAqs6mZMf/3VqR7vqLPPycu4IMfOr77kvo+40bbOfQYMIdOcGW9P69utYyBmh9tw8UT8Cvf3p/NmB6wCvTaCYeOGi1XadS5rcDX3Ga68iHkSrR4wwM0i+Z7v27NLqLUfv6FAJ+gu12T5Yn9XMj7nYcyBezwEzvSjJMYi9JmMlVDM1rfE88EzfrEl+hnGCSgu2U/f6vp1+miedcqlf6Mf41jGZPRJ9GG1LdFvMPZB0M8+lAS4j6S/gzN1cq6PyMO7IPQ3+9N3u9pjD4oPF8QcYbvbGBdG21BucH6vmCx3ehxM3xeweLGNdyFtYjzIeADLPd5L9K8k4lJstDEBjAhYD3MUJLCij6TPxFUnlgv0k4wxt1nCYoJ3IPm4HpyDewm+vNvIR9/LNUNZgTKE/pj+Dd701eznvJzTWddxvfiba8q7hrz0KZw7VDBN3ej/KZ97hecKTpyDfNSDMsmH4oiyaDsbihv20fcT84FYLZ7WdsH8h3w4hUUa7ne/In1/R+nATlzgoQR//80pkz6Z8yFjlagbLtzIRD/79pRXDrjOCz+wSIlSZZ07qKUL/PuEG29v2ZZjGac7t4SuLCxBWrTr1JW/iR8XpXLw5lozJuE+5H5FScF9zvud54U+knECzyb9NeMF3uVYraK84z7m+rNYhfEDygXuQ/oFxoTcY9w/bpzHPck9y9iK+5Fz8SxyjLMg5DnhvmIMw71KH/CiPRfr7BmJW7Flx2oTAREQARGIkYAUFjGCUjYREAERiJMAkzUmkgx4mSgzCGcwziouZ/5/VUiZCDCZTIWvGmUQzcSYyQmJQTR53cZgmQE652GQzoSc8+GLm4koA2smYgz6OY6yELwyIWCgjlCPQT95mSQy+XYBEBmkM8ml7tTZrUwMOf2hXwkojbsKBBWtml592YY1K5mYxrWhJECYhxClYrWaF/opLDC/N7dRmP7nwG96JLdTCN/I9+svP3kGIHX+y/GdTr4mzVu3wxT+lZeGPR8uQEPQQ55ILk5YpUseAgxiqk87Kle/oA6+wgm2Ggrk7Dz5AuVhyv+rWV+Ew2LSiMKC30cPfvapUPck/Fb38isb1bYg5TCf/PKoYX6wg8oKhA1M7FgJysoxJnUn2j7uHa4zAjiEBtxHTATd/YqQwwnnEB4xaTyw0v9w/UEHFQ0IIALWK8Gy3Up+Z6bPM0QeZwXAd1cHvjs3P85FBc8P9z5McQHBPRwoy+obqrCBA88XXGZb4jkI+O+3fDxfOUJcgnAeVvIz0ee7ey6cVQG8OAf7nCsQ8rvVvK6NToEyyvY56yUmyzyvTIzhwH1BP8I14lpcZgkBDN9pEy4aEE5xb9Nmnmcm5CgcENJF2lw/4gRw5A08Sz4bbeC+8BKQRTlVYDdCovCN1Y4oTFHYOEEW7GgD9yNcYIKwCcESAgcEVTDnutBnYQ3FKlpYcQ04hvuUfQgt6L/cylmOQ4AWWF1sCWZcIwRs/IawysUIoSx3L9rXw99QJOC6A2Xs02YlFa1EW3BPH5zj1NPOQFAX81a+8n5FQiSf416FIYQ/14JRsM+8Ii29+Y5W96FcIYDsB+amL/yYKtUvvMj9hrLCyxVJlaCfdSwn/IK/1rv6upvoU1l9i8Dcr6HUD0E5+/2UxXM+eOdNhPoXXd6wERZ34X2lX9mFLQZHaHBzlN/uXRB+zJlWWVcH2hW+P5eZgJhnrYBijvfNjbe1aIP1R58uHVp7nd/F3di2ZRPPge9GrKYnBo2cAAN8xHe+965bwtvX4v79wkE23qME0vYrsNR5FQNCT9wwovD+escXn+PPPpYbDSsOrBVR8IffG7S/c59nA0qVyS+PHOriQcVSbkgenj2eS+qPVSrPLn0IYytn8UVfRJ/Nb/SRKGl5/lHYONdETshO0ShBef+zL9R1UWjVXL9J/0yf0NLStmCG0L7SWRrwWyQrgjibHVf2ePpip6zgBLSLhKUGzxNCWJR7CIMZHwQsbUPeefSRtJExKn0kTBHo00fTT6LMpt/mumAd4jb2OaE/C24QLodu5GeMyXk5fn3YsQfGF8FyGLOQ2FAqhO934wRXF4TSjOdoK+9f2uqU3twv/M07k2vNu4Vn2Smzwqoa/c8ywfgVaVEURy/94BzFzH8dv6Cs4Dln/BtLGVhEMV4k7xsTx46M1D+GWh0v8VFisrDn4iuuvJbyJr00/IXQOtCnD5s4/UPq+NbkiWM/spgYMdSRe4L3N4lnlXc373/GY4zn3HfmSoz3alvi3uR97hYkFLDvbqEC5TF2YDzLb5SBIpTnlncw9wfjB+5TrCewbHLjAvdcc07uD8ZbjCvYz/j+76DSgnpoEwEREAERyAACUlhkAFQVKQIiIAJGgAEuE18mfyeY0HMvK9bsOxO8GZaYGDGBQ4DBZPANSwinMNVnIMzgmcE3wiNcvTBpRtA52xLKCYR87OcYJosItJi8cj78x35siVWJnI/9rDRjUs+Ek9XmTPo4hn2sQGIwz8akwK0uRBlCPQOC3TABbzD7wR9MXh7rP3gUgqWeD7VtsW7VCueGwDN/pB+XLZw/D4UF7kj88hFHAmE+VgcuvoRfXreKNTxQq8vv3FcgVEMgdPOd99yHWxIvVxd5CxRiUpMD/+R+53MumpyQ7s62+1cq4+M9fJLofLxvtzgbXhPIqjVrX8xEE6HXjDdfnxR6zuoX1r2s96AXsSLIwWpbXLdEgc3kimvLGAChLwIIVstzTyGE4d5zZvNYCXG/4T4AYRECAO45JnwIihASI0xCoE95CB6Y/DMpZGLH/eaUBAhBKJ97jXuefTwjCBOcSwpWuCKsd64bUKpRDr+zwo1jEDggMORYBPOUR10KWOK+5m8mlAhVEKgy0cSPNoIJVj1zf39v9aXt1JdzcwwrQGkrKzkPEUKG+Eh2QuyDLFTsGLaACx+fzSs/WQOr6IPCIZ6/gKIkuNE+BHZOMUNfAEf4UWeYP2uJ5xs+1A1m9A11ggnFCgJs8qLo6BIse17wd/7knM6aAesIJvNO2cO52Vi1fDgb9UMwAHcEStxTMKFfRLhJ3+WEDu7aOp7OfQdt5n7lOO4DykGwQR0pxykZ2M937l82eDnBGdf3oC09rYuuuOb6JoVtZfmPZkGFRQKCdRQUFmt0d7enBo0IuE6a9PJorKVw84awybZ9JjPe99tvv/7KandXOSzU+M7Kd6y1ECyH1z38b/IisEeQTqydaPlD99PHOMXuulXLlgwaM+UdlMCmXAkEUw3dLEzCGS5OA5YDfsL9KjVrB1aL4wbJz/VI46Z38n7LMe3VcaPDrThCz4nPdrfi168fnzpxzIusICbvBRdf3pBYQbEwCBXOcQ1CY3WEH58nfwGeMVNYf8X79ZCtZJlyFVEuoMAhSDjfn+3d9SE/dy1FS5RGUJZjs8XuiFRXrBZ5r2Cx+EjbO5vgXz40P9YVTlkVKM/ei5H82TurQt7b5B/Sv3f3WPzfk/fqG265g89Xx744JHShAH7x+48Y/zpuYrZu2rCOMmPh7/L4+KLH5QvPMP0y7wCedfozxlmMe+i76T9oB/0YQk5+p79gDML7gvcb7rF4L/C+C7X08qoi7yW3IajkXUf/xDuQ9wjvmlmWCljC0gALMFZq0x/z/sRlDwJa+hvOh6ULfTd1ob+mP0JJiyKBRR20i++8Z50LGsp2QnWE/fTLvM+c0gUG9I30dyifaD99JjzcanDejWwwow/G+sq5U3KKWsqjL4UXdWcM4SWEpe3UgzZw7wUUEsFr5vrXSEpev32hio1gdQMfrkz3W6x/u3xwIbn3uVuswhiYd65bEMH7Y6UleNLH0vbwc4XWy/N7qXIVqzBmjGQhFrWQGDLwDnFKTrJjrReLCzfyMqYm1gR9SCTLZfKWLFuee9pc1e3+df2alcxXDtlqXnTpFTzzuIVbt2o5SqzARjychx/v/zzKCgJ6dzd3VZGa5vPcO4XWbrtWjIXcPcqYknEbzz9jSp5L7m36ZZ47ngMXx4ux0IeWeKZ4NjiOeQ/fsaRwCyXcfIrneqwlpwRl/sFzyxiJY2gj4wrqw7s67vskEgftEwEREAEROJiAFBa6I0RABEQgYwgweGbyyUTp2+DEyCkhnI9dXA28ZQnBm5tYMcHlbybnziSaSRam1AzMmUg5ITCDeY5j0onygcks+5msM5mcbYlVSNSBAb2buLGPSRnvAHwVs5LOrVQ7rMF341ub30PgUHzVvvvGawhX07y5yQ/CN79CLjfhIPsmjhr6XKQTseIzd558BcjDxCo8LytrCwbPg4KBOBNMtAY/3bubl5DJYtqiDMqxJUIQwqIl9wuhVi1b9ClKFyxPsBrxMtt3blj8ykPoRVkW22OyW9FLne++v1O321vd/xAT0Bf69nrUy91IaFuD15r7ifsToT7CEe41JutM9rg3uFeY3CGUqW2JSRr3IoJ1hBkIhLhPmMjhVoHfuAevsoQAb5sl3FxwP3J/M6nkGAQ+ztoHgUFAGGsbwhMUQEz+ELSECopYcYkSAWEUQhRWylE/JppuhStlUDfufawP2BAwUTc26sG14P5HMMHkk9+c0AaBEufGhQTl8rt7RoNFZPxHhKCRsHbKDie0o0JOsA3HbSGrYVHMsCFYGmiJfgKhLVx5zkdacisIEWbRT6EEQIAHF1auwonri7CZa4+AwK1OpVysFLBeoH/h/ChZuQ9QrnAO7jHKgC0CAYQdKFG5l6gH98QTlrhvuG7kp55uhax9PcjSxgnF+N1tAUVPlC2qgD9aAfHsR5j8+MARvi42XFkoQ0leZaPAMEOpX1Fy7P3zz4DCBgFVp179BhH0FCVwJJc95SpVq0H+tSuWLfZa/R+pPU45TJ+HSyOUEu+9OfmVjWtXha+MznGRrdJ1yoORz/f3tIqgX6p9yRVXcs457789zevcxLdwig/cQUWqn/XRgWcape4X2z7jeT1k22ZKZPpYFLm49ItdYbHfIo7t9QkvjYgUNwmFFPkQyHvVwbWHGCQX1Wt4TSR3hVjPwJlyIin47fV1bov79sdqGvrskz3CV3FzzVt37NortD5+QkaXp6j5jnLfidcxfcpEBHVRN97xtBFFxXvTJrMyP7Dhiqrns8PG8D7DWgN3kGm0rohUB/pD+gwSfSB9DP2Rs3ZjXMO7geTeJezjPUJ/gzBzsiWeLZQY9H8o3QtYog+j/6Rsxgnkpf9jTMXmxkf0nyh/6YN4n1DWS8Hv1In+ktXm9NckFqnwyeYs7FxZ/O3ccbr+b1m+qwAAIABJREFUj+OdEN/N1Z2w3ymQ+dtZmlAubeUYyqDObmEAdXXl0x7esXdZ4t7FhRB9dmAsGYxb8XlwnBCs7kEfnIP2Uj+4HdZ40esEmflbUFHtlNzu+qSpCsRSQwnNwplYrbrSdCI7yBbf5EfZ7Y4fN+L5Z2Itq1bderhSy0Fg7F3ffxuwHvXbKlSpXot9NoZd4OfW1ZU3851pKO0CruDu7dS9T/XaF9fjb5QpPTq2uSsWZXsMbeBaOeVTaN/rnhvaw/iFe57nhvxcV55PfmOfsxaiHBQZjGsYX7mxFWXRT3CP0x9wHBZIjIdRSDKeoY/guWFcktTPQAzMlUUEREAEspSAFBZZil8nFwERSGECDHgZCLsVQEf4DGyZSIYK1RhEH7RqMsjoQLwDH2ZbTGDJSrvQjRVBTqjjJfA7sOI7PQbdCExwfUEFxo94gVWGh7XhSokCUBywQjU8OC3CEXyj87uXu5LQk7PaE+EZv3kJhfBdzgpmBHz4QH962LjJWDO8PGLQIRNB3EQhsKEs3Dv5NdKtgNuweuWyJiG+vr3yOwXIJgt067WfVWz87iaFCMHadOz6OAHBmQgOfLz7w17Bbr3KCl5rJ4AJZAkqrBAaI+hwbpW4F1Ew8InAEkEMAkMEIawI5b5F0cDqfVabkQ+hN2Uw0UNBgQIBKxQEckwaOYbv5EXYg6Dc+R92VhFOmYIQBYUFyiEmiSjqEDCxH8VIqMICgRX1RsiOEJ66hrpYQ/DOOVldRz1QSFAOz4dTyLC6GQsnBPHOqsi+JscWovBwE+hQAUzo9wMu0ey6036XnxXAgWckuKFQ7W2JCTzXgjEj++EMH4RXfLqxpBMEOOsG9zt/hwrWKO8QQUkUhU1SXISt1nfgmgPh8okmvGLlugUtPQFlKa6V6F9w+XakdWj0aXzyjb7JxbvhJ/o8UmijsSZzfzepf2HltSuXBSybwjcXjHWZKY3jhRbqg/2WFm3aI6QaYkpbr3IaXnvTrfyOu6j1Fu/CK0/FqjUucPE3Zr775uteeeqYKzt+pwwvZXLoMa5tWKJFEoQPfabPYygssDbADV+0WCGcw7kERAg/YdSQiApwp9ixsB2eFhEu6Lm7hrim8nNXiJ94zo+Qc/3q5b4WicQ+YSUzSpIRz/V9PJwllj1cP87DCm/qGOn9xPHEmHDlTBg5eGCssaZ4H/G+x2oGKxPilLRo1/HRa2++vQX3L+/Yji1vabzz6y+d8jTeW/GQ/BH6hwA+68voY5zQkXeLO3dAmOmOD1lVT7/He4ON71icBcqy5JQKB+oR4fyhym0/RXcsitNQwWeoJYKfZV44o1CrwNDvKPgDm7WdMSHvSLdSnXr9GTr+c9/D22vHUj/e9wixeSfj798pO8Lrku3+ds/8yqUL52d048193QGrYxbYxOp2lXdMxWo1LqR+s96bzvvdd8Pazi0WiuRa0PXJKLmfGvzSpIvrX30dfQOWcvR70187NN5aWvhEef7ds+MWd3g9h/wW/nski1iq+VtwIQhjVBbhoCThvYyFRiRLorQ0UceIgAiIgAh4EJDCQreFCIiACGQMAVbkMGFG4Jspm8+APtNW/7CqEjccuJSYO/N9/Mof1maLjFH6BDZbTHZiuAuQKjX2uxrBt66fexB3fNVatS/mOwEBd3238xCXME5o9NmG9Wtq1Lnkclw0DbTA2JjChzfCCasQMPkJhJjsodhAePS9nQ9hEqt+vXwbI6x0E0OviacLjMr5/mvL6sZNn73QBVxEudKlXYtb43X9Et6m4IpKhByhgg7c9yCUYEOAQ0Ip5qxxEIQgGMIvMMe9YgkXAgi0ERwxcWeCh8CFslBIYAmE8gVBOa7L+BvrC1a6oehAMcJEGmUfCg8SVhWs6mSyyf080xKKDs7LCn+EMJyP76yide6omNSzappjR1taaAlFB8qMfawmtc/AZpNSJqFYsbBqkTodIrByeVPp0xiETrrdSlPXxGhCtkPcZoWx8fPrnGl9UmZfK1wevfhcP5Q8BzaE1pNmzA8oIns82Kb5Wz5BThHyIJC2zR7zE05EwUHq+NhTA+iPEOibvuPP78zlGwGu/dpWtmKVgJXRskXznQA2ZgxlK1YNHPs/W/LPOXEZgsVCeAH0V+48+Cb3O8ElDa5uzD4sNFjB75XPuYya+e50T4VG6DFVa9YJ9ONrli/hWfbdVi5ZON9ZWdzeun2naAoLLEUItE2BuLaK5l4Fl0/kXb18sWc9nIUFeXCXRX38KusU29vN8s/rfcNxCEMvaXBNgOWAPt06hSsWzIDw2La2qpn9WDY6xdOWjf73CSu0XSwm7lvclMV6ozghJYqRdp17PnVDsxatqQOLB8YMHdhv0JM9OocH4Y617LTmi1XhGbKqnlOF9kV+CoO0VilRj0NZzLPGGPXHOBer8H7kvUrfz7sDBbYEtwbB9YcrIjzr6XVDOAsvypv2auzPLX360UfnCsSu+nTebMZcvtulDRpd73auXPKpZ/9FDBtnudy+a2+swHMQh2j8iy8MYAGNX5yh9OKQieUwhmXMyhjVWVZl4ul1KhEQARHIvgSksMi+114tFwERyDgCTOBwX4PADyEq/vczfNVVxjUntpLdhG3j2tUr/HyVx1bS/lzHnXAC1imBzcu1iVvRtujjjxBgR9wuNF/mZPjIArJ6ZXTCqg1rVixr0rxVOxQgr4weOsgrb6Hg6jaEWn6rfIsFhV9fbt+25fKrr7+ZSeKwZ5/o4VUergTcJHK9WWOE5ylZpnxAOIZQrd/QsYHAt998uWP7UCuPyWqsq2KjMYqi8CK4YPhKT1anuVV6CPjZj9sfJsSsvncui7C2YB+/k1i9jLLAufBA+MGz4lb3O1c/KEZcvAZ3bo5x/qVRZDj3GOHNu9x+uN8SVhbvWBrDOSIIZ7CYIWGBgSuQWFe1RsOq/dmYAEqIHs8MGX3m2efk+dDcufkpK0CEchNlL4n+h6DK/N7wupubIWhCoD98wJM9I+HETVwp8ztOWfEGfqWuTtBdqlyFyihI/c5H4HDqQb/sZzmBIha3UeSbMX1qaCDeg5rgzrnokzkR+3EsNdw7hsDa0W4r+lusLHDFR//u5dbKlZH/3CLFELjzNy5MIpXNtURhQ7+7YvEC+ruDNqzvyMOPsQTDtfgVAQsLcxHvaTHDvrvueyjgCgol1JwZh7rWwi0g50RYiMJgwjtzA5YaFsPbV7FVKCQ21CyL8xGPcLFEUGFz9Y23BvzSc7+hKHmhX6+u0ZQ90a6b9mc4ARYPELsJiy2/wON+lXDWv9sswyGuNTO85gl8grIVqpzPc4DVUUZX09YGBfoM+hcUorGeD0ti8v5g8ZWcBbPfsfUb3dDU7fNbEJP/3MJYvAY2LK0mjRnxwmvjRg7FOjnWOiVJPudqDesi+mkUF9pEQAREQAQygYAUFpkAWacQARHIlgRwYYNrGVzlsBo8ZVcVu6uLWwi+swI4Pa746WechT/9HCg/EMSEl+kELusiuNHgGCw/3CrWWe96m8FbSIr9AThNaFfp/Fq1iV3hp4xw8SYimeEXKb5fCIWLmOtvbd6KFb5+AkRXHpNIr4DZ+QsVwed0YMPVxviRLwx4743JExNkBatbXek+w12cUe1oK/Ej3S7RVvkfsroz6PKDeBy4hkLAgpXHP1FWkvKc4tecZ/YQC5z0uJ9VRvYj0Lztg50vtBgOWHb17HTf3WkhYG7GA/2peZhC+R1xK1G2XEWsNLCKiBS82quQc4sUL+mCL6P4IHaFl3UFbkUaNLrxFspYPH/ebGJteJVXqVrNC4nPwL4Pg/7Nw/PxzkARgXIkmluTyxpeewNKW5QkH896HyVkxI3+FndVVWpceNG1TW5r0adzh9Z+B1h3HYhfgcBxzozIyhACW5MXVyxeFhFOkU6eNydPGIP7qkgVddZ9BDn3yodFn3MJONCsK8Lz4DP+jjYdHuZ3FEx2m2CxloPA4X5BwdnvFCV8f3dq7PGmUGw5QSXv5emTx48Z/+LgAV73SrRrpP2ZToB5P1ZKvOe45+N1G4cbRd6VBSxVsMQCimjv6ExvZGaf8Njjjjue5wmL13j73bTU1Y1nA9bFcSgH8lq8IM63Ye0qXHr6bli9uUU8KM792nT2OfmwgM2xecPa1TfVq1UhneJUpAVJRh/Dc0PMFqzwWIxDHDBtIiACIiACmUDAb2ViJpxapxABERCBlCbAKnB8/TPQxQ1Nym8uCKB5NMH1z2Fvzq2GxZllJf1BG0ITC18RmCzhliLSyRo2vrkZ+1EGIGDzyusmgAijUFRMjODDvHCxEgH/wZEmfS7gNsIoAqq+OOjpg9zEhNbBuZjyK48Ai+Rn5drNV9SqiE/gzFZWHPbFzKQCgv6GncsqzopQBtcX0Tae04ssNbCEX/fQMqIdq/0icAgB4szc80DnHqyCfbjNHTfFI1gKLQzf4Px9bEiQVT/cLg5DNJdJXsc76wW3b+Qg70DaF1xcrwGuqsg394N3pvvVpe4VV+JiLQdxKQgW7pXP5F0ITnN8bf6ivJTSoce4fnzuB+9OjzWQ86SXhj9PGfWuanwTsRX86orQn30I3rxcBoYed2nD/a5SsJjxKq+0uW/id5Qfo1945slIjwZ1Ig4Rebys6/i98a133hMIom4WGOG+5FEs9Xx26BiUSKyCHjPsuaddW3Zs37rFL24G5TpFCdxxnxWpnqH7TjEllLMIbFjzvMK9H2nfSsqKWOlleT7m/SjciBuDS8d4Y4wQ+wprYSwfD8RRyPJWZXEFzqtYtToWZWlxwxdv1VFI5y+437Jhlk9cIL8ynUJ6x+dbAvHh/LZmLe970O3zi0/E/v+dckpgbLX7l19+TmFlBU3k3YGrUe573I6itNAmAiIgAiKQCQSksMgEyDqFCIhAtiNA34o7HPzis5rtSkspLwD96Ydd33OlbdFsICD14W7OjZNXwD98vDNx4xyRBIH/PfbY4665qVlz8k1+edQwr0kVq4BRKpCHIN6Tx48aFmmVXGwWFvuDmVIeVhGfzp1FQGPP7YACZM1Kz1VvtmI2MCn8ySSXh8s0mxyPNROBpT+1xGpQVqiHBp0+CIMpOXheUVagGHLBwLMJKjUzIwiwOrXXgOFjETT3e6zT/ZGClkY7/49mekUe4vhEy1sgaI213lzbRcsbvr9shcrV3G8Lzb+5nwulBtftD7aNMNwv7gTtxrKEfF4ujNx5zBgg0O9GU+acV6lqdRe3Z+LoYZ6u+rzaO9vcJ6HwIY6IO94rnxnYBSws/AKZu2OITVTNXEyhhHp/+uuTvMpyLq6W2urnaEHEC5grKif89+KNQgLLEs7D+yv8fG07detN4GzciBHLiHo55fvOr77E7Y/vVrTE/pgdn8ye8W48Lhzd+4hj9U6K9ynL8vy4XUTwyoIaYsrgjz+eDUGts/jkneoXpyieMpM+b0WzJqMRmaGwKGTmwE75Sv8WDzwbNxODJOASyu+4qrXqXIwrPbd/dYR4QcfYAJt8Xi5b46lXEuSFG4pl4r8wpmR8qU0EREAERCATCEhhkQmQdQoREIFsRwCBKf0rE0KEpe7vlAZhluMEZA64YDot6M4prQ2mDBeM9Z2pkw7xKf5fs8GnbPyIR1qZ2/iW5vcgrEJR8dq4UUO96uNWmrryJowcPNCv3ig33OriTevWBALphm8oUohL4X4fN/y5/pE4OAsLvwDeByaFe/YejmultF6KZDzOKQe3W+VRnuGqLJLCkOcTc38EfDMscV1T3oVbMl7YZKgzyooh49+YgbIUq6h4BOxe7TOXUAEXZbnz5i8Qrf3OVc/m9WsPsUqLdmyohcWr40YO8cqfy6znnDAL4Zyfy6Hipc+r4OI4fGQWEX7nhhH7dv/ys6dbKXfcnW0eeITvWEAsnj93drS2uP0I8Fcu3R/wuljJ/VYUXptzf7J1k7cliDvmxtvuboNbqlnvTZ+68+svD1mdjqKmZNn9MYf8YnuEnt+9e4hJ5BVDguDWBLblPcc5Q4+94prrm9zSom0HfsPdFe5o+O7uAa/6ueOpp1NsxCv0dLE+cOMF31ivhfIlDAHehQhfL7UUry9+FuE4ywremXItbRBwO8fVXbJg3pyMvsrOlRt9Ff1GPOdzz+7ff//jGaMLS61OPfoSY+zAFikmh3VLgXL+tb4gnnokYV7cMaI4RmGHdUqgvT5x35KweaqyCIiACCQuASksEvfaqGYiIALJSwBhJzEsEDCvspQtVsazUhO/2ZjG33DbXb7+wqNdVoQpj/Tu/wL51q1aviTSCi/OxSpUrzJRVDjf3lMnjHnRKz4Ex7FC1R2P8ObrHV/gp9lzK1SsRCl2/GaO2/2EdYWKFitJvci3y6SN77/pvRKX/dSdgLp89wuQmo0mhdFujVj3I4SpYgnTfQKDY+0UzcIJU/8LLDW2hJ/naPljrYvyZSMCrK4fPumtWSg1EVj36eIfNyFWLK6fIcaE61f8jnV9SbSAquHHn2CdZUEz9eJ3FMBzP3zvLa9zVK15YV2UFuyLFOy1bjDYNq6bYgn+7ZSyXudk9XKtupfVZ9+IAX17xcrN5XOriU846STeyYdsZ5yV+xynhI5k6YF1xU23390Wy5JRPq6eYIj1Hyf5eNaMqHE2nPARRYxX3SpUrUGflGPT+jWrnGsw/sZdYrd+z7/I96kTx7z4xqRxo9zxeYJ+6p3Fo1e5ufPkK+BcOM6fHbs7KMrS+yjeOzCh8jM2JR4YSjyssHg/xrOhoMCVFBvKqmzvGsdZbxHrIdLYMR7IkfKaMjhgDbZ88YKP4y3Txdw58+zcebyOve2edh0LFC5aPFTZ6beQhuO/2/k11gY5UKrGW5cky/+r1Zf+3Fkues45kqxNqq4IiIAIJAUBKSyS4jKpkiIgAklIAGVFTUuVLCEwTfUVSDkQTk19ZWwgGN0drdp3chYS8V67ezo88pgT1Dzd45HACtLwDeGNc+8Uas0Qmq9Dtz79TWdxCsqFwf17d/OrR6HiJQ/4Yp5sK6Ij1dcUFoG85h58s295FiTV7Zv2yrhRkXz7Mjl05v1fbPvMs8xsNCmM91bxy4+ygdXPuLhBeYECKtLzR34moAg0cZehTQTiJtDo5tvuGj7p7VkIsBD4P9z6jptYGR93QWEHmPAo4NqH1bGhgZK9ynWWbdYVI2A5sFWufkGdpne1vt+vLvS3KIrZT0BrXAx55a110X7FAUL7D9+e5hnDgf0uSPRys8KI1P9ZWKFAfCeE7O78oefFXVKXPs8GrD1Y6UsgcK964TLqzrYPPOIVpyJ/0E3W9zu/CQQvD99cvCF+d8oYr3wPdHviGazn3ps2eaKf66hS5SpU5liUTNHcQZHPWTls/Wy/dUT4Zh6jSvLbxrWrV7h9WIMMGPnKNNigDCKGhNtH+3nn8Xckt4ZO6PnFti2bUap7ndvvt+92fhMQUnIup5yJ53jlzVICvA9RUmDRxHWP15KQ9+oISwSIZ7yS7RX7tSymD4rkSG4/0/OKFy1VJmAptmXT+rXxlutcBdaoc8nl4Qt9UAy3bP9wd8qcN/P9t/nEgurnn34kbonn5hTjeQsUKuzVd2KNVr/RDU2fe+m1t1C4x1vfBMrPc4Iimr4VqxZZliXQxVFVREAEUpuAFBapfX3VOhEQgawjwIQQ4Sd+8XEPFFhxn+rbwD5dOyEEYQL33OhJ03FbEU+bb2/dvtNd9z30KMewatTPxB4h2NoVyxaTr+4VVwWCu4Zu9a667qYrGze5jd+e7PrgvZF89joLC8zrF8ydhUsg3825b9ppS+n8MrnyEOq9bqtfI5e3XwFiOpWf3eq38PxuUmjzvQOWIKF5zDvW8Xfd27HLMy9OmIpJfzy8UzQvripwdxFwN2Pbxhja+aHlYQXd7GBKeQVjDEyUJQYCKAn6DR372qNPDhyGUuGdqa+Ob9/85mvSy683fRdKV6oSKQ4D+3PlyhVw8eKCq/K9Wq06l7zw8uvv3d+5V18/AXOl82vVdk2d8dbUV/2azcp+9hHg2SlSw/NybieIX2lKhkgI169evnTfvr17iSFUvkr1WuF5O/Z4aiBKXRQo3Tq0usOvrC5PDBjapmPXx5s2P1gpc+EllzesYOWiOFr4yZyZXse7QOXsczFAwvOx8hirEawW+j32cHu/erjrs2zhJ3NjuHUOBL7esW2rZxDck4Pxi1wcE3M3VclZ8LCiu8NdTRrBz53rmGOOCVi/sPkpndhX7DCEnj+YgsO5YTSXVp7vJFxZ9Rs2bvIlDa7BYk1b4hDgnYj7IiwQGSvEq1DFOoN7DKUHruqyvRzh2ia3t+Dy0tcxFkMR4KV8TY9bgHKLmcKSsiJZHvudC0U68WqIrdapV79BbrzIGHrg6Feno4RECeriDnG+SG3hPYBVCdZaNzT7f6tqFBXEMJr47rxlxHJCQXL8iScm82IQ5nFYQrOwhXmH3LOmxw2tMkRABEQgBgLyPRkDJGURAREQgTQQONOOwd8vK9AKZJeJHYKMu66vX2egKStYCfr4wBHjrrrhljvGDR/U/5M5H77n5/O6WKmy5dp36dXPWWUQpPaJLh3aROJObAv8rjdred+DCz+e/aELbHtRvYbXPNZ/cMBFBu4y3nx1/Et+5TAZK2BRDNk/Zfzo4fjljnROF3A7krsNt5Js0cdzZqK8OdzyPnhr6mv3PdLjycrmJ7lM+UpVVy1bTDDpHPh/hy3KCgR+uDPJeXTOoyOtaE7DfZyMh7ASLuBT2jZWhO6O0ghWzzEBZRUzk1LcG2yzFO/q02RkpTqngQCCcFt8+leN2pfUu7bJbS1Yec9z90LfXo/6uQtKw2kOHMJqfYTVJK/gyy7jD7u++xYFCn3gmKED+yE06jNo5HgEU9TLKT7C61K+yvlYAwYUp3NmvPOmV10p49yi+1fJRopLcfY5efMhsCLf1s2RY0KgpP3IzofArHOfZwa3vOmqS1CEcDwKCISBKH57PdyuZaSyFs6b8yHK5FYPdO6BxQD9M1YlTe5s1Y56THtt/Et+/t6Ll94fcJut/rU33jJm2MCnnWsXruvd7R7qimtB3g3dH2h1xy4zMfC7liXLVsCiMsea5UsXRbveWOK4OB+//77bs49ycS1QOjVp3qpdy/aPdEchRPta39Lo8nDrCHhSv1NPP/OsWhdf3mD65IljuabhdSlWar9bmdXLliyMVs/w/XCY+c60KbBCkdN+yc3XuPemxfGu0KJdp661L61/1X4O8Zcfb32UPy4C+yw3Fr8oNlE+kOLZUFSwsv87S7iVilfhEc+5Ej4vll3lK+/vO7v1HTSC5CrNWHefaRP3/3/v/k/7duC7/XbQfvbZhv0afS3KZeIEDezTrZMr85x8Bc7ld57ztDy7jBFfHTtyCH0JFoEX17/6un179+yhv+AcWC53adfiVnc+Fh7hMs8vHg5986vjXhxyb6fufdp17vkU70Usu4hhhFKEcjjn44/cf8/KJftjCSXphnLPBdqWO6gkvYiqtgiIQHISkMIiOa+bai0CIpD4BBASIADNZ4mVndlG+Mnk5vZGl9ZEcHHznffcR0BCEoKT9atXLEP45gQxp5sz3VImhGMVrbukuP3o8WCb5sTDiHSZcT/VtEXb9ufkzV9wxKS3Z8//aOb7x9pKL1bUchwrnXt2uu/uSGUg3GNVHOd67eXI7qAox8WwsPjivooI56JqrClpot2mhYPuqCKVRzBzlD0Eux32ylszF33y0Sybz+ZEeeFWUn+2cd2ah9vceXOkAOTR6pIi+1EQHhtsC88glhPRhCpOqYhlBpNSjss2z2uKXPdMawbudJ41lzyhJ0QYQ7wK+reMqAjKWJQVof2k13k+nTv7AwTJCI8QIrmYF++/OWXSoCcfCwSuDt9YEeyCP0+dOHak38p8lBXOjci8me8FXIZ4bSbjP7DK/+sd233jAbljhz77ZI8LTNCFonfyzIVrcK2C8oG2YhnxVLeH7pv+2oQxkbi+NGRAX6z5sEjo+czQgxTUsOvX/aGA4sJrKxb0Cb9u1YqlCNwnvDNv6SezP3iXvFVqXHARwjwE8j0fureFnzKHvLAuWqJUWb5j/RDtPgh1ZWiGMZ7BjwkwjmUHyn9cUlEmQsVWTa+5zAXZDj/Pyy8OHsC1533x9PCXp9x9Y8O64XmchcWnpuiPVk+v/QgprzBXLyjEXv1gwaotG9evxfWWsy5EODt68LNPcV3SUr6OSX8Cy774BSViAUsoKXDFhkVhvK5tyE9gaSyGiWWBAiTbbigPUEzw7OMSlQUwR+W0/2yAhrXCfhd1B7rDuDn9Hubaz1lXvGkK2LQuTBn01GOd859buChu+1CaukotNauwxx5ofaez6EVpe3aevPlxS+ensOBYFOMly5SriPLDuXLldywDJ9uYetzw55+J5J4ubihZd8AaOzVuQ7Fo0/gw666DziwCIpDNCEhhkc0uuJorAiKQKQQQgDKoRfC5wRI+T7PVxuTt2ccf7TjppeEvsJKrfqMbmxK0FNcjoe5HHBQEQotNEI+QA8VDLLBQMrS7/YYrEcog/HF+01l9OvTZJ3pMHDX0uWjlsEKM1WpP93i4fWhQU6/jWPV7pM1A2bfChGB+ZSPww52V8wMcqQ7OJN9Zh/jl7W7uUIZMeGMGQj0XgJa8+DEeO2xQfyawftYr0Rik4H5cD/D88YkCIqLVTPm8J/5jwhxc7iy3hO/+gI92bSLgRcA8avxJ30OfhWUXfVysfVZaib5msXWua3r73auD1lV+5Qzq26NLKQv8jWsjhGi4/5hg/eDAJ7oHLAS8jitftXot4iGgRB7tE0ya4yw0QiCwKgKtdauW48Pec/vC9tMX/WQdKsGio7WZoK6d772rKauTCf6N4Itjtm7asO6Jrg+2XTgvulCdmBEmxK9HGVjrueMnjx817JXRw5/3E+5xPos/fS75u7VveVtfc+2FMO/yqxvf7OpNex8zBTqT4NlOAAAgAElEQVTKg0htOc0UG86PeyQXhK4MrCPghFDTwpR4jhGmvDx6GEoALFD+sqXZuHQZ0r9Pdz8BYq9xi44Y0v22p1HiX3PjrXe6hQGh9SZALpYdBPomLki06+O1H7cxz/Ts/EC7Lr368k5yVoXcb+9ajI+Rg57uE0sMj7ScW8ccFgFWiqOkYhHNLkuMVeMVvm6xY3AtxbvygDuyw6pVkh6MYvP8omcd98+///wTPv5CuYvy9hgzhcVVoP07lr/pa+3fMfb9mJz2xR5/U3HkzIl2I0cwjhBjSGLF8JyFotm+9bNNWNgNerK7p/I5Foy8u9o2u64+inczLi5lhh57Nq5dtSL8eR3Sv3f38y+se+ni+fMi9nu0+8GWtzbGHR59L+1mAQ3WISk0JkVBR8wXXMFuTcMzE8ulUR4REAEREAEPAtk+WJbuChEQARFIbwIm/KRvxedpn+CEcIJ9vmWC0XhXs6V31bK0PFZrlSxTvqLJdXKfcOLJJx9hCoBff/npJ9wmITiJFNwvUsURzJWrVK2GyWDyffftzq9XLvl0fjTrjLSCQOmCqTv+itMjoC4WEgTS3WhCOy/XHaH1RLBVtWbti/PkK3guPgbwYYywL61tScXj7NmjWYUsPWjpAksPWHrP0t/2/Pk22Y7D1Q2rDQlWzEq6gFVGpGNSkZ/aFBsBFI1/mzQGhWdsRxx+LvyE+8W5CS0dxeqZuc/Ji2DM5PhfRIplwHEEvL717rYd3nn91fEImfxqyurhOpc1uBphVDRhNCttv7eI2gjYYm05lm4cx6pf3gn0b2nhy/EoZ6L1p9QLt1HDXpk+EzdKF1cocjb9cb2rG99kOozCvI/MpdGihR/P+TCaq0DXRlxx2WG7ln768UextJtYH0fbhcIXfLT8pow4KEuXpoH43oENRYV9kFxMgX/eHP3kMQ1ve8itBmbfP3bMPyhVOvd+ZjDWD1zLaOeNtD+3aXsqVKtxAYqfr77Yvg2ljp/bscM5j449fAL2jmOxBe6LnNXvn/Z++z7WkoPvVpcdAS4K0ED/p/dkrBSVL9kIBO97xofVLeEOEIUfyjrd98l2MVVfERCBpCQghUVSXjZVWgREIJEJBAe4p1gdCR6d2xKKi5Ws5E7keqtuIpDsBILPHj4YEMoQEBa3FwE/3VEUFriDwiIDH92sPNVkNNlvBtU/UwgEheUHncsE45mmyDmcRt7Som2H9o8+3g9XT+3uuOHKwykro4/1U1iEKCsQIiOURtlK4hqgwGBVPfv4jf4tR7Jcn4xmmp3Kt3cj9wAxmnBbhkXPRnsn4tZJmwiIgA+B4JgSKzyeG1wc4uo3MJeTok63jQiIgAhkPAG5hMp4xjqDCIhA9iTAgNYF5/xNyorseROo1VlCAL/aCGQQzgUEdNE2ez5328SUvNHiXUQrSvtFIFsQCArQ3cKnA65lkkkYXqJMuQpcrGQIDh1qUeFusKCygiCwJCw46b/4dIsjUFoErCssOYXGXxyXTNcpWzxQGd9IFFdFg/fHmfaJC0RtIiAC0Qng3hdrwR2ub5WyIjo05RABERCB9CAghUV6UFQZIiACInAoAQQIX1tab+k7ARIBEcg0Ak7pgM/hmFd6Z3eXbZl2dXSipCcQoqw46PlKNiF48VJly3Mx1qxYEtUlU4JeNCwoGGvwiaI23O0k14ffUVow53MWF3/bNcRFVMz9Y4K2X9WKnQDXf5slFFe/2vtuT+yHKqcIZGsCKCxY0KJnJlvfBmq8CIhAVhCQwiIrqOucIiAC2YEAbmnwc8qKHPziaxMBEcgcAk4Ix6piuWHLHOaHfZYQ10KeQlSvFeaHfVIVkCYCwWsRep2STvBNINz8FpwcALHEkEgTqAw8yJ4Xp3zIZaf5za5JpBhZ/1p+FLkIq48N9ot/2m9/2XGyKsvA65RARaO42maJz2wdLDuBromqkuAEgpYUf5kFrsaSCX6tVD0REIHUJOCCs6Vm69QqERABEcg6Arvt1Pg7/cwGvBIIxHAdLMDqEWEpRybGtI2hhsqSRAR45g4IZWS+nzRXLukE30lDVhU9iEDRkmXOI0D5js+3fkaA7WTCE1RWMIc7zhLWE1EF0ATctnwoNRBYo7hA0fEfrxgkycRCdY2ZANf9d3sXEmxbwteYsSmjCATiVfwTTIpdoRtCBERABDKRgCwsMhG2TiUCIpCtCKCw2GxJ1hXBy+6jfEDY4vygkxNBChuCSybVfEqIma0enbQ3NkQxoXsm7Rgz7MjwwMEhJ5JP/QyjroK9CJQoHYxfkZzuoHhnOgsLBNGxLoogH25NXDwLyjgQf0R3SuoSkJIida+tWiYCIiACIiACqUpAFhapemXVLhEQgawmgBABv6exChKyur5ZcX6nrHDCE/c3ny6QqLO6yIr66ZwiIAIiIAIpSKB46WD8iuVLkyp+RdAignckFhLHWGKsEdMWjFnhxiQsWuP4nEGLjZjKUCYREAEREAEREAEREAERyAwCsrDIDMo6hwiIQLYiEFzlLZP7yFfdWVWgrMgZFL7g1oK4H27VJ8IUvvO7GWj86ywuDir5iCNCDTSy1a2mxopAKhDQCu9UuIpJ1oaSZctXosqrly9ZmGRV53nhnUksCmJlxbX4DNdQpqDgncqiAN6xuImKFP8iyfCouiIgAiIgAiIgAiIgAqlAQAqLVLiKaoMIiIAIJBeBUEsK3kPHW3KrPRG+OIUFygz3HWUF352rqORqsWorAiKQwydwttx36d7IVAJH5zrmmEJFS5T6+6+//lq7avmSTD354Z/MPS8oGZxrqHiVfn8G36Ucx7tVWv/Dvy4qQQREQAREQAREQAREIB0JSGGRjjBVlAiIgAiIQNwEEJRgVYEQ5kRLrBplw23F6ZZ2WWI1KUIV56ubT8W2iBu1DhABEUgPAnuaHyjlgKA31wjF2kkPtplRRoky51U48qijjlq/esWyPX/+wfsn2TYXQPv3YMXjUvrhGipoZcEiAFmDJtvVV31FQAREQAREQAREIBsQkMIiG1xkNVEEREAEEpQAQhZcUyD0Q1lxqqUTLP1i6WtLuKw4ObiPJuy0hICGROBQtrgENQnKQdUSARFIPgL0W1iB0QcdYUoMhL9OmXpIa0yhoS1BCJQpX6kqVVm9bPGnCVKleKvBPYdSP/RdGFcZQddQHBOwajQFxr5gjItAOfZ34NPHKiqucymzCIiACIiACIiACIiACMRLIC6/p/EWrvwiIAIiIAIiEIGAE/idZHnOssQnCoszLSH4Q5mBuygUF/+zRJBREn/z6dxFCXKMBCwOiAtifuAzxkOVTQRE4FACKCzoj1C40n9hISb3Ogl+p5QpX7kaVUzC+BWOLMoKXELxjkxz/AmUFna8lP4Jfr+qeiIgAiIgAiIgAiKQHQlIYZEdr7raLAIiIAJZS8AJSBDsIeBD0IfQBaFfUUv5LaG4YEMYiFDwXEtlLeEm6hRLKDAC+4JC+KxtUQKc3TgQmZyEMsJ9/499h1EgWTWxrMTFFp8kftdYIAGuX3atgq3kPsKt5k5CBjw7Z1sqYqlA8JN+TFsCEyhXuVoNqrdy6aIFCVxNz6oFrSCcS8T0cGeF0gIFiDYREAEREAEREAEREAERSBgCElIkzKVQRURABEQgWxFwgbcJ/ulcQuH+iYQ7KH5HoO4sL4BT0BJKC37D8gLBe7Z/jzklRZCFC1qOcgI+WKIcE/wMtUhh/3HBPEdZGaRQRYdTeGSrm1KNzVwCKCsy94zpejaneEXpyjOWJ5hQYPB8aUtAAmfnyZv/jLNyn/PD9999u3XzhnUJWMVYquRcQh12LKcQBUgs51UeERABERABERABERABEcgUAophkSmYdRIREAEREIEwAggqWdmJSwviUZxjCUEfrqAQpDt3UeRhFSmKDH7/wRIxLhDUnGHpG0vOJUZKu7ZAMeGxOcUPu1wGFBMIUPkbK5T/BlnzN6zxe45AlTzs4/fdwWvBSluttvUird/SnUCoz/x0LzxzCqS/+tXST5Z47niWTgv2S66fSul+KXMwp99Zylc+vyalLf3044/Sr9TMLSkYNDs9+2ndo5l7CXU2ERABERABERABERCBKASksNAtIgIiIAIikBUEUEQgbEfIx/ctlnIHhX0oIlBQ4BoKX+MIBFFmkJ/A27iNYnNCdoSG+4IC/UMEL0cckcyLuCNeGtcwZ02BAAsWKCJgB1c2XG6h6EFZ4VxswZqV4fD/zRLHUp4LZp6ewrCIjdBOEUhiAihLsQbDuqJAyDOFAvZ9S/RdPEsSCCfIRa5QtcYFVGXJgnlzEqRKh1MN7q3DtjL0Uhwq2PbhXBYdKwIiIAIiIAIiIAIicLgEDnuQe7gV0PEiIAIiIALZlgDuilyQWgR7qyz9HBTA4PYJF1DsL2QJoTtCP+fmaLt9R1iD4t0J27MLSKfogQUWEighiOtBnA8UFfjTh1loQqkBv1MtIUwlL8dhbUE8EBRCxAfBioW8KavlyS43idqZaQTos+iHGFPnCz6TVe3z4uDzhgJRz1OmXY7IJ6pQpXotciyeP292glQpTdUIUTI4xXSaytFBIiACIiACIiACIiACIpCIBGRhkYhXRXUSAREQgdQn4ITugcDPlhCa84k7FVYtnxkU8qGMQOCHZcWPlrCq2GqpWDAvFgHfWcKygOOce6hUJQg3JxyFF8HJ+Q2FRV5LKH7g9IUllA9YqxAEGAUQ3+H0pSUUFXxHieGuAd9hjZsuuYZK1TtI7UpvAvRB6y3hFopnjmeIZ/MSSwiT3ws+o7KySG/yaShvwdxZM96fPmXS5g1rV6fh8IQ6JAVcqiUUT1VGBERABERABERABEQgcQhoxVfiXAvVRAREQARSmkBYDAbePwj22AigjYsitlKWEK6vsITyorwlLDFwu4KbKITpKC2wBuC3jy0tsYRbI3zG89tB7oyS3SVUkJtT8PDpgvzCAg4oK1A+wBFmCElXWkJoWs8Syh2UFCiF+FxqaVeQFUoMhKzfBrlyTeCI8JXYIf8kOz9rgzYRSFcCe5ofUhzPDQrD+sHnEIslrJ9QpqKwoI9yMS0OOjjXiHStmgoTAREQAREQAREQAREQAREQgaQnIJdQSX8J1QAREAERSFoCziLCCdtZ9b/A0veWvraEcH2zJfI5ywIE9AjqF1paawm3RrhhQeiOgBBrgVRTxvOuxv2TayMKHJQPKChQzuAuC4UN1hXsgwH7WNGNMoPkFB742mdFOEyxzqBcApcjTOU4eHIs5XDeVGNpTdImAulOgD6JfmyHpQ3B5xLFYWFLKAx5BnnWtImACIiACIiACIiACIiACIiACEQhIJdQukVEQAREQASyggDCdAR6vIewGEAYj3CPjdgLKCZYtcxKZQTs2yxhWYFFwKLgMcRhQKmBgB0BPgoPBO0I8ZPONZSHBUqo2yzaBSMYoJxAscDftJ24FAhDawS/o+zhWKwo4IOlBC6iYAJ3rFlKW0KwSiwQNudmivI5FusMfuMayZVNEJI+RAACWEWEWVnwjPCs8bygFMTdUBlLWC652DtOAXjQ8+TKkaWF7i0REAEREAEREAEREAEREAER2E9ACgvdCSIgAiIgAllFAMEdygXcOCFkZ8U/LqEICo0wntgLKCzWWcJNFC6hENDXtsSKZawCWNmMIBAB+w/Bv1FwUG4yCtpDLRqcFaQLKk4bsSJBmYNVBXxghSKCQNuVLDnXNCh9nPUE+8mHsgdrFPztf2aJIOcEB0bRQ9wLFB/kRSFCPeC4zxQpfP9XrqGMgjYRCBIIUzD8a4oHLCxwpUZfRV/0ZvA54rllH7/zrOEmKhn7Jl17ERABEfg/9t4DzK6rvPdeu5w6vWjUpZFkyd2yZdywDTamOjgEAhgCBIc4hHDDhXtzk5CEPMl3PyCElJt8IYCT0HINCSZgE8ChGGxs4ybbsmzLtmyVUR1piqafusv3/rbOGp85c84UaSSNRmvNs55zZte1/qvss///9b6vQcAgYBAwCBgEDAIGAYPASUHACBYnBWZzE4OAQcAgYBCoggCrkUmIDiQEiT2SOyVDqEPOYzkBib5F8o2lYwnADYnOfiwPtCsojoMchOgnT4hlcRq1AGXn+UzdIrFAMmIO9cRP/uoSVggLiBeQoNQdIQIsESX4H1GHAOUcp0ULHaSb63Mc14JkxdICSxfujWspxAruPyZChSFXT6POY4p6ShFgrOEWCgFxg2TGGeOSccZ4It0vGasnkwwCBgGDgEHAIGAQMAgYBAwCBgGDgEGgCgJGsDDdwiBgEDAIGARONQKQ7MRRgDCHHIdkJ3g0FgAQ9JDsJGJbsJ9A21eW9hHLAhdHiB2sYtZkP4S7JvtPdf1men8ttCBMYCmBlQmWFJCbCDdYVOBuBqsTVnBjbXKtZIQZsFkjGWuUTskIFI9LBgfOQwDCigKrFFxFgc0myfwOQCQaKl0XfCFcOZ9yOGJhEbmFMhYWgoJJJxSBT96Ot7coMRZwe6Zdu2kXcjXFs0+897ITWrYZXlyPRcbUeZIvlcz8pePL4HKNuDy7GFMzvKY5zCBgEDAIGAQMAgYBg4BBwCBgEDAInFEIGMHijGpuU1mDgEHAIHDqEKhBeAclQhwrATKkO2Q97oxwa8SqZAj6N5e2QZ7/smSIfAh1Vi7jUuocycRpeEoywgfb5lUci4oYFbohtAsoHTOC5zJCBfWHsEWsgLzFGgKxgk9tecL/4PNTyeDCim6EHhIYQp5eXzqe83ALhTUFwg7WF7ioQShCMNLxMbgv55E5jvLo2BelS5sPg8CJQQDRQUQLHetBWxkxDhgn9Ecd3Fr30eMuyN9tfSvX1uIm9+Q740lbgCEshB/f+ZXKe+k4Mhw/JhMSx/tDdzdTToRDxqYew4w1xiRCI3Mcc5W2LDvuOpgLzE8EwnuUZb3WCFMno3XKxM5yt4rjouA8ETRPBhTmHgYBg4BBwCBgEDAIGAQWBAJGsFgQzWgqYRAwCBgETmsEdGBnVh8jNCA4QLxD+EHyYSWgLQr4X7sugszHAgPLAbZD2GsLAq413+NYlIsVlF8Ts+BBPAlEGYjNiyVrN1AIM2wnIT4clKzdQEH0bpX8qOSNkhF8wJNEQOAnSjjxP9jpld8IRXznOhzPJ2Xg83R1q1Wq9qn7SH5nkPagD0OaQWJrK4Gqhcq9DSOhk5ekfDqoe7klUs0g6yerfEIsBkI+6hgqyaLodbGj2gHjHkGNfomIRt/UfXXW1goloYLfwVgqaYFTWzIRZ4Jt7GN8FD+z7jf8kmjBOGUMYtnFnKPHCgG29zXdOHhIRAssKrgG8xbioI5DwzjmeCzDdJ+IGl3I7amSnitq1lOIcZNOMQLShjqeEiWhb9myjXbW7cd3xGn6MW2pBeHy+aFqG5/p7VsmSFRrZY2vFh/BWMfI0gLkrOeIU9ydzO0NAgYBg4BBwCBgEDAInNEIGMHijG5+U3mDgEHAIDAvEIBIgIBEbICAxxIAwQJLAkg/SEm2L5YM6Q6Jf0OJkICIhzjEjRSBu7mGJtnLV1rOi4qWFUKTxRArEKCw1YgWbKeeZ0lGtCBGBSQnZC2rtPnkeCxJfiwZootjOR+3UOABXgTTJnEtSDQIMjACO0h0vXodV1CatH2pdA64s53zDMlTAmUmHyURQK/Sp63WlmFJu+COizgHs8ZVCPbyIpQTdPpa+rOqK7SPbbxz/HwpJ2WknekXkPT0Kdq7SzJiVmRVMJM6n4hjPplerxYFBctWYVC07PySIF+8odAXNoVFyq3JXe1CrbL+0xZJsORcxAiEB8S9ZyUzNhA6uT6iwgWSsVBCSmD+ib9t0Vcz3+9/96JCkGBccf7rJDPvIB5eJ/lFyT++5LonD2y5bxNuoR6QjOs1hA3EVdpfjz0de6ZaefW8oC09+J+kRdh5ZT1WrQILbdsUghLjjXFEWzGmsAiknRlT9CHiA9E/2E//OlcyzzcELqzk6Fucj0BG/+E43QcXGownoj5apNDPK8YK7aCFYu5ZEMEjUj1FED1l89qJqLy5pkHAIGAQMAgYBAwCBoGFioARLBZqy5p6GQQMAgaB0wcBTSxA5ELu4J4IErVTMiQO5A/fIXsgCjtKn9QQEgKCFaHiOcmQQNp9DPurkrfzABrKxTMYUhvSlPpqv/3UCfGBukK8aNEBAhRiCxKcldtdkrWrp5/Jd4SIsyUjYCB+/EQyBCfXhsQBX3BiHyIP12A/14RQA1/uTTlImiw1BE8JkKk+SmIFWENYgidk5Bsl05ZgSrB4MMcCRosWs8G23CKHovC/JrKdVCavAsd284lYfTJX8CWPSeCRwvrt+/zLHn1e/c6tSn1l1S3WDzvemHzAH1uas5PLfMvhGsRZgFSnfP8uuUsy4gp9pabFxQwgmfUhZVYp7b12fJ0IFhTw8IjjuIOJJYfeXOgZ6Qjy1FlbWMyqfCWrCs5nzDFWmDsYQ7TPayS/STJEM5ZMtOHlkveHyvqSH7qpzuRLfasTO0a6cuvTXhhrlO2vlv2IhYwhPp+U3LgrvfZHH73w75/7+2c+ypxEG3MvxhdxeUjEnnnYuUAdlqz7APMB92bMI4ZQBj4RD8nMFU9L5jj+1y6lZtOHSrc3H3OAgLamoL1w84XATB8gdgl9h9hBV0veJhkBgphCWAO+SjLPMNqPPoc1Ds8t+uJdpbbFpRjzBvOzcclXu7HKxQotYDKGtEtEfea4pSDChREt5qD3m0sYBAwCBgGDgEHAIGAQOMEIGMHiBANsLm8QMAgYBAwCM0YAYgayATIXsgbSYbtkyB1WKONahX1kVkNrl0bcoFMyhCvHIHpAAuk0n9walbus0KvbISXZjuCAOAPRdaFktrPiljgTF0lmJTfxKhAbEC2uK2EASc6qXaIOQ3xByGrCBqsK6o+lBteF9OQ71+A4yDQsK8CYDHaQa9qFDcG2DSEqgMwg0X60QafkLsk3Sb5Z8guSaQfwhhy/XfK9krGGgaSMVv5WWFDo22mRQgeT15YRy6wwXCQihe0EwdJCPLbI9f1s0VIHHD+olwZb4nj+vqahsVz9aLZrqKGhfkg19x2u6/CW5btXLc8e6BiMNS8+Em/d6FkupCmEKwki/R8kE3idMUa5PXEHdcL7QEmsoA9SFvrz4kBZiHSer6w13XayeHti+U//Z3YXfXy8PLMkHyGXsVSinXCZtkUyMXHeoAGv/BRRYoUfOn92pLiouDu34eARb9FYMYxDSuukA2rzP8IPOfODxTfuuGD4mfDmA3d0N3rDzGPc9+eSW2S0XywSR7e1aIIo1Cn7mNOY3/Q45Zr8z3bmAOZBxjFzAVZWzHmIF4xXHXOjVlXM9uNHoNwyjvmZuZQ2YdwwvpmLXykZgUqnG0tfeL7Veu9CoODZ9wvJ9EvEzkdK59HGiIfGqmZi++m20IsS6P/aMokj9dyqhQx9vHF1ePzjwFzBIGAQMAgYBAwCBgGDwAlHQL8In/AbmRsYBAwCBgGDgEFgKgQkKLUm7SGCIC1xoQJZB/nzCskQ6ZBzrFrmWMghSAqIf8hAVi9DZuLehU8IHsiJeUG6l+qnV8RTZuqJcAChgosQvlNf3IhA2BK7A5cy1BkXWNQHl1i/Uvr+PfkEJ0hwSC7EGgiv70v+Jcngw/UgwiCgWd2PexvEIAhRSFdW/CKSUB6OBbfIZ7/kyMKiRrB02XVmJiHWKyuuiTAsYT4qGQsXXHLh2ozECbQjIhIuhEifl/yvkumr4B3qGBEE6uWAv18UBYOmbzTGih66UX3Rca9L5QueFQTLPMe5xvGCzmLcXSEdvC9e8EZbBkZ2jTSk6tmezuTiy/f3/jCeL+7zfXfJAWtV7tHk1bFVg/taC2Fi+30t1137YNs1m8acOsbOhGSp8DYh6ulH90q56Bdzlmrgp8c+K9IZ97skf0oy/+sEAfkhyf8hGcurCQS9xm8K4Qf8mUuwXHiP5DfPpFKCg8r6dWpX7mw16LWpHx95a1gIkjP5/fzbySC3+RPbP9n9kd2fWy+Xeb3kHqGsm6y4rMZPqe3uK9RjVlNEeiN6MIZxD4RQRJ+4SjLWZswL60vlhrxmnsMShLF+h+Sdkhm/7KsZyPtMj4EwXVvPIIYIczfzpp63z5fviEj0Q+ZSLKsume4+NfYjOHH9+yUzz9O/aE8sNn4k+VuS6f9Y6bB/kji10Nu3SgwLbWEWxQopywh6GkOeoYwl7f5O/+/NUug8xmad+WlV+p9e3IA4q91d1RQlF3r7zxxJc6RBwCBgEDAIGAQMAgsFAWNhsVBa0tTDIGAQMAgsDAS0/25WlEKUQuRD5uAKhZWsEOmQc3xCzml3UJDFEK/a/Q7Pt3kRdFuEClqm0p2PdmUDiYp7GlaWIzxArkBYQqywqhqyEiKTuiJAEFoXEku7HMGdD/WE8NSrS1k9DsHJdVnJzz0QJSDYKAdua1jxzfUhctiHZQUF1Zhpd1CyyaQpENCWD7QJ5DJtiBshLVZwKvuwtsBSRqcPyxfaDFLywNtidwVfvyfCnzZM9LmNscszL8QP2m32gGpYL+6dmpKFfNjb2vJbnuuc5foqk0/E10Q2OUdTq2yXxg0hTC3fsVUu1YhS92GhNgsHFi0OY7tjA/XDQx3d6SXB88nz+3oSi1RzcbBeBItJ1YsFxRtsFbSl/Oy++q8/s/3Zey+MhL9SrgpH4l+OuZ/QJykE/RWx7vWScbUEOVye6Ktfk8w4QOwBv5msOqeNuD7zA4IFq9crxQqEO9oCMWNCQkcd9FrV3tw6daiwUs1QrOAat+XtxG23rfvQ7e/q+2ay3et3xBxmudWgVktOWcvUuVZd5B6I+YzxeItk+g1zG5YlCF/V0ltKGxn7eq5A5KF/YXXBnGjS3CFA/6HvkcGZMUo/fYdkbT1xvHfTQjb9oTIxl3dJ5vn3Q8lYPfGcmJU7tOMt4Dw9X7vlslzXjssMZXt+UGfb0eM2DIKQcc8sSdtpkZPnYZYFiioAACAASURBVFYEEP9kihY1BDEtSpRbi5QLMIhjOmg7QgwxvfhtwHxM+2vrknnaPKZYBgGDgEHAIGAQMAgYBI4dASNYHDt25kyDgEHAIGAQmFsEIEQhICFjsCpgtT+iBUSDXjnMSzuEI5YGWA7wHMOlEds4H2IC8p9zIDO0r/sT7tJmCig0qcIhlA8ilm2QXwgylBGhhRW61AXikRX6Ol4HggKuZDgHP+kIDRx7jWQIDCwtIHgRJCBkuSZkLoQG91td+g65AU569SkYIQxxP45nv3YHZdzLCBjTpPIVvqySxxqATBvphEsviEZSpSXDLSIwNDZbQ7ePhvXP3+9dk7089tiiAbc+3ms3rYn73oUxz/Pr3NyVgWutPlLXuK7guvQJJZ9VizaWTlr12awwqoEaSqXU2PKUEOyJuIgPKrvBXfJc/zr1w5FftUWQWJIICmGvu6iqpUDBjp8lbozcjUNP3/DOg3cUtzZuHNw4vJU+wticSxdr9Gn6MxZFEIm4Z7p+Gtz/Tvbjyok5YDpRUhOBiEaQwVgm/GqV6zOv6D4P4c+4UUFoq1G/Se0W64otI1epEZ/LzDyJdcZvj8br+u649F0/u/Xwlx6sa8q8xaqXsZ0Qy6WUWEQ5EZmKWzaspnSjImDUEisqb/5XsoE54P+VzLiH4HxIMqTmdNjMvCJn5pF6fGs3YvRP5mUs2X5bMuLkiUxYXyGMIFjfKZl5m7nln0rfeUYyJudyPJ7I+hzXtUVcmHC+triIxxw7lYz5QahSgRcmbMd3xBytQVzmqYIXZFQY8jtBtIuQZxtjjHbVViqn4ndBuUiBUMWznHmAeVA/u/k9QFlxL0c/0+7Etsp3Fm+Um/kx1qnbqajLcbWpOdkgYBAwCBgEDAIGAYPAVAgYwcL0D4OAQcAgYBCYTwjoVf6seEakgKCFcIe0gVDErRGkHOQRRAQMIi/0j0nmpZ7zIPB0QGte5iHmT3gqWVJU3kcTptr6AYsJVpJD1OJOhAQ5AQkGaYqIASlGgoyCLGPlN26wqO/FpWPAgBgIuO1BdIDcQoyA7ITQwKUOcTAQb8CNFduIIRAbxFSgXGCJWKGDumqxwhAfpQYo/6jhygjxiRXQ75T8+1VO02JFlV1qsRDav5NS2faElb/zsN2+77Db8op+u6FoBWpxWzD8qqLjtD2aXgppOeM0KkIFCVdGoRDuA1678obS6ulwk3pgBOMFWV4sva810Ws1FweE+cJgYXIadhs7n208/xO/uXfksnp/dKfEuviBG3pdciQEKa5pGFuBWFYca39hDIBfp2SsUoilgRukmaS/loN+VzJ9PRrfVVxB0ce5PiQgK+Eh9cvFpPL7IID8H8mIfghL/YLfBnGddb7kJ9piPZ0iVuhxOX5eys6opYl9o7kgtV+sMLozfj2sKmNzPGVV6ncfbrjy3Bta7hu9wNl2teUGayoqOJGJnUntJx6DWPb3knE7hksp+iPB03Vsi9lf8cw9Q5PJEMjMx8zL9AnIZBL9k37KXHssibHzt5J5rm0s5WrXYU6vtDDimfYHkiGtee4h5iNORXGHZAX/lBZQC9FlkAgVdiLuxusSbqro+e0qYdf5vh0vFPw2iX/T4IZBfxBYjgBTZ4fqiKgWuEZkIQTPSU9Ej/AkWlno3wL8dqH9mXi1m0DmQp7FV0reXPpO/CN+KyBe8uzHFRyxq5jg+W2EyMsznfgnA9L+iBjMyVXn44XY/tUGjtlmEDAIGAQMAgYBg8DCQcAIFgunLU1NDAIGAYPAQkBAv2yXuyaCkIQghdjHdQpxACD22QYRD7nDqmiIQAhJyCZe3tmuXdmcCmw0QQHZAImJaEFGQKAuJLbjxgVhgeNI1AtSAt/0HAcm7MN6ApGD60KkQUhSZwhLyA7IC3DgWpAYP5GMixncYjxcui7fEUIgNrgOGOnV2GZFdqkBZvABdvQz2g/yC3KRfkr78r9OO+QLK6KfEvngLUKC/7fKax8Ml74j5l9w/hXBo3du9LdcGbP9FtfxN+5JLHa6YzTz7BNiRZ2fV2PiEWVX9hy1yz9HbRtjse7LSYJIqxa3X12WeEDtHTtLxb2C2ueiDb6c+uLtLV9a9YF3fea5j4tJgL1KeiLBnhEFIc8Qxbrztx615plOuKgi+IATfZV+hyUKpHtlQlSrBgIkP4WlDNVIOtqHMcRxWGwQs6KWWME9Py4Z8YNMWxYEn9FfDL1uVWfyxYKIFayonyBYNLlH1Nnpp5UfxuoTdtYRsWJgf27tP/V5Hf9Djh23XMmpZNOecNXGZ+3z1y1yeoWp7FF2KOvBi2KtEo/G5lwk7qfdCSFUImZSFwSMUzkHzkXdTtY1wBACWVuxMa/Sh/gER9Q+BhFzsXZNWK1sCAk/LR3DNSGZ2cY4Ya7/jmTIZvr23ZIRNRFEEEGYP5jLtTVHtet/vbSRa+HC7AeSEbQRnrnPGWFxsaGz3RoZy1uu4zSLB6hG27ZbvCBcEwYqLQZobWJy0WjF3D3iIuqIZakGx7Z7CsXA93w/IcKFfv6dFJdKIiboZz8LFrDCQ6zg+U3CXSBtxvMdkex91RpdtnEu6TfL9rM4408ls2ABcYN+yu8GfgeY53kNIM1mg4BBwCBgEDAIGARODwSMYHF6tJMppUHAIGAQOJMQ0FYWkOmQwIgPrHpmFSIuaRAteHknFoMmPVlFrUUMiGTIOu0W6VRgV+4uiGctxCSfkIfUBWIJkgkCDDIDooFVs49Lhqx6o2QIB1Z+Q0SBBZYk1A2/9RBcEMes/oXQhaTQ/u8hY1iVD/EFKcb1IdZxLcU5iCDgRnkg3nSAbflq0gwQ0Cv3O+VYCMNXSiaeAO1GQiyCkPyq5Add5W29KXb3C0/6F+/vCRct9UN3U0HFOHc87QlWn7fTX9M2aDUv3p9oVHslvoQIHFMWJSEeTnB7srLYqzq8QRULPVUX5NSBWLvqtVtUrGCpR73z1bbspki0qJbGgnq1JLVPhcL4xe28uvDQVnV3Cq9ML6cGb1T1JBar5bmD74sH4zGdsezRAZ8RZcZEuNBuVrzpxIvS1SHYwI7xAKmLUDfBOkH+f0Qy4+R/VSn/+2Ubq6UflVxuRaVjVkAEQwKyahkLrVqJ8xkzlJ9x5O3NneXe1fdeq6ew7Oyd2XPrjxQ7WFU/IZ2dfka1xvpUm9ujVid3rBdLjFWHxtY8+LOBN+89GCyboPyIlcW67cF65Xqeep37U9VsDVpWPPKvP5NEvA76FuObvgdmUyXmBKxFcJ31oGTwq7nyeiYFWMjHlILcM0dCFtNnmGe7JCNMXCv5VsmRK7ZpEuI5czFCAs8fLCG4Bm1H3AnmXW31Qn9FYObZBnkNwcz9tbUd/Y0+y3OtVsLajswYoH05Fus5rAiY0xds2rJv2BoayUUigLh/agp8v7Xoq7a4qxblMl5bqPy0Zdtpy3IcV0wuikU/LbPpMtex0uLmzbNU0COCBu01IFYWxRNhZSH9SgcCR/TScareLd+Z43g2v0HydaX/j7WtENO+WHYyAhgCFlYa9Dn610zi/Bzr/c15BgGDgEHAIGAQMAgYBE4YAkawOGHQmgsbBAwCBgGDwHEigCUCpD3kOi/9kHWQMfh8h9yHCOIT8h4Snxd0iE9IIQgbCCCIoay4axJewzpW1zWzrYYWKyCrEBjKg/7yP9vxWw3hwmpuVoBDWFEPBAzOh+CgLhCfkFDURQcbZ1U6gg11p37gAEHO9SAnwIhjEXdYgQmhhVCBgMPx2qIicoshGYyDk4iP3O60TrQnbUCA67dLJggyZLtO35UvrLB+st4avf9PEn858LH4P6g/zH3qyAvB2VteCs7ydgednZUIfCX/G4uzsZha42yRxqa5qqcWf0S1e8NqXf6gKtgxlbESqt7PqrQsGk4HeZUMiqoh9NUjhStVwvVUtqi92Uy8XqM7qC5ruF+8qGTVpQ0PqpgIFv1J4WVxQFaWdtSfpX6w+Ea5x6i6ZGgL1gHsJWg1GXIWYhyCjH4YjVERL6hAcQrhgr4K2UZfpO8Sw6FSrADH/5TM2P+gZCxVytMvyT+4QYJ4JDO+teULQoUeD0f9YE1OiHlflcwYYLwxLkc/tvHO4tL/3OkMeG2Qz22HC8txJ6VXN0dXaY31Cma/UHXOsGoWSwvH8oh3kbDqgte82/vX/u+Pvs3f7m/QgZSVtLn6bP731Pti31AN1oh6rfszGaBVOWX6DfX9hWRc/TBGfyQZPCkfoiO4fUDyJ2rUi81YXmGx8m3JtM9WIVDHxC2MiU1TAq0kVJTPzQg9ZOZk+hLtfssUGJfv+n/kH2KqEEuIz/slM6fruEx6xbt2OQVhzb1J2hpHP88QshCqIaIhuKcS2zgfF1OMw/9PMqLFfZKxsFmQbY1Y0T+YSeTzXlysJppc11peVOFay1FtEmx7recGzeIFSmwpQj8IVKsTc+P5oi8aRlAn+i7xuPfIgOf9l98JLBzQLhFn2NTTH1YSK5g/eM6jFrMAgfmA78x3PM9PRKLPkrHiYe6kHzKPnBFWNycCUHNNg4BBwCBgEDAIGAROHQJGsDh12Js7GwQMAgaBCQiUYiBoQoN9msgo9009iXQXonkhIqnJR+qmrSpYYQxRDKUKCc/KVP6H4IHQ65IMCQQTCBHKflYYaiuCkyFYlLcfBKNeuQvJSFlhj8mQpRzLcxgyi+8QTAgU5atwcXlDHc6TDAHCSl+uCQHBCl3EGyxLiOGBWx0EEQQOtkGKIV5AynAPvdISjMaDkRuhQtCYeaKdIJHpW5gbaDWAdoJYpD3jYh3xnLhl6m9UIwNvd78TEZefSv7Zhp6w/c0v+htGHw0ve+Fvch87ZyScKCb8wnulWhk+EwV7dqyXOSZXBIg2f1gtzR9RLeGINL6jUuLCaWnUjeSmsh8LC0cYubzw2vslTMK+Yqd6Mb9edXsMm4lpRaJLrU9vU2elnlMtYiVQ56BlSUeTeBcX1T+mnh4lpMTR9Hz9OVFek9mtzhl5YUedL/6jXk6s8P6qZATDf5QMEYfFAgQqq8UZu5VJx3OhTyM6YClRLX1BNiIEcTwEfGViXEMuQwpiocT/mvRFSIJ8RlSplrjuv0lm/OBOhTllALGCg0WsoGGwmiEeBL7kJ6QVid25ttjhZFLEHsQKEu3V5A5YVl2m/bPhH6i3DN816b7PBuepK4NHI1ddTYWhAZUJt0mP2W8lZd6KRZY5rMon8R2rKvoTcxtCI/MDcxi4EqOCY3FfhHBRK6YCAcYRchFBaBeuecanklhBX2FOxaKCPv0KmrGEJfFopntHouGJpUL7QA4juN0umXmXOTyyahGRqPy5U/59AoksZWI+YSDSvlyD/czfWNTQn3VMiy753lnRiIzDL0uGoNb3jkTDiuNO+3+7e0dsy7ZifhjWhyqU56UIFl5wsbiDardV0JAt+MlC0c+I17XAdrAcc9an4rEwDIKDRT8YFXdQYnQRStuGiJCRO0mxsrDmysqi5P6JSZd4J3zSv7Dyor8wTitjk5yINnkb9ZKMcEU/ypZiXHgV/fFE3Ntc0yBgEDAIGAQMAgYBg8CcIDDdj/E5uYm5iEHAIGAQMAjMCAHIUMhkPTfzqYllvVpYEx4LcvVkBUraNZQWHNgNEc8LOKQOhBOMLaQAxCjHQ9gjDIAj+8BPr2SdUSPMwUHaLzbENgQuq7cpK/VAXIGwYB8krw4SDqFIeXHf0lk6D1GGmAEcz3mslIRg1TESWMmLBQXCCOdyDOQt/4MHxBUrsqk/mGmXPVEfEqHiTOhDVHUuE9jSVoxHiCj6GgliG3yfFxdQfW1W/wuyin7nZ5N/srjVOoIlzKsd5V3YYfVdIT5K1L5wiVoW26e2F+DsX04xq6gOFVaolDOmklZWGi5QZ+/fK6z0iMr7MdXSO6zaUqMH0vV5O1bwDrj1wW7HDhqtIBwWI6Jn805i/f5gee6LhQ8u6VGLLrvXe/UkVzarnL3q5tTX1YpYl8rHfeXJkmOMj4h70RE7qC6s2yzCRasSt0gTypYQd1AjbkMu7Wd2iiBTueqbcfkZyYhoiBWR5ZNYWuAuqlCytNACHWIPq4w/IhmXO9USbD99FvdvEL/Mhbg3uqYcLvmO/3csEPS8yThjfDAPVIoVjCfa6x7KJBmCGUKYezBeIgJZYm1wLcrPfh1rZkIZl9iH/t2VFdxplb8o7ziXafddiBdWPFBeOq8+7H1efT7z4QnnPeNfoPqctsH7u6762Wt7f/poor6QsepUa5hSL9hNQjYnIsKa8VkedyKAZBTCUSfEFlxXMR/Q58D8a5JriRa404Iw/aBcI7IEMpYWUR/plMyzA9EHLPn+G5JxCzVdwnXfJyUzv0IMIwrThxCXI3H4GIlh2p7z6ZeIFswzrJb/S8mIK8Rv+vUpCod7NepF/+HZoeManQyxfjrMjnu/CAt2T/9orL4ukZJR0iCLPFYVimGdxKlI5vK4gZI2CC2ZL8IGqXBcZN+4WFkk4zErH/g25hWHcl6QdJyg4MswlQIxn/N8RbSoGfNBxIwZlb0kVjDncgJuvZgXuc/EiX7qqyFE8jxHNaZf0Tf5nUA/1QLrH8t3RFXEyFoWOO+SffweYCED1/uKZIT1BdEXZtQg5iCDgEHAIGAQMAgYBE5rBIxgcVo3nym8QcAgsBAQKFlWQJJBTmi/x3xCjGr3PdFLtWS9KpPtOi3kF1DtFornFWQeL94QAri+AA9IHYh7CEoIelZKQ0JwHsdD3IDlyTZD0ZYWulz8z2pHyoS7GkhbCCgICeoCqUGGJYbMhZzAJRSrQCHCIE9pZwhg/kec4DqsrEW0QPzQwckhN+hL9BG2gZ3uRwgVC7m/SFVPWKINIcTBHiKbdiJWCImxuk3c/PzNUvuQLS6g4u+O3XFtozWMxQzE+VUiCOwK5Ap11qg6y9muNlpPqD5/kRoOmlUxPKpBZYUCf3b0FVH8igvcp9RrnnlC1Q1mRViIFepa8j9qSY1uj2W8Q44nDk+S1n43DCAlW6WHJ7JWaudP/evDH3uvvfSh4MrfORAsw6pnUrrA3qYu9F5Sl1hPqnDMV3c3vmxNIRYCUSyLZdl9kwSLB9quybQX+jKv6/1JX8rP1iLJEG6IbQE+d0omBsV9IlwcVHc355tuHKRfghnEai2xgtXkjGvIX/qyjuXyc/leLlhQN9xyHUnZmYQIPfaS+H7taopyVCbECoj+z5WuzRhDIBwTy4pyP+/a6gky8J2SJwglLdbgt52C80RbcSQ8x9td/0R63TibSbuFTqC2p5epi4ti0FAhWHgyFP+58JvBTfXfH75i5LEj8d7+TDigDoqFxRNhWg2Id6/iDMQExi/jmrmNPolF1V9IhszGtVa1BG6flkxA8JwQqz0zuE+NS52+m0uuesDsIslYVCBMISgzVgjeUnXMyHbmbZ7B9AWsW5jLIZZpB/aNxwg5RqGiHFRtUakDxkQr5CXTR5n/sQyi7LR3ZUJswUUUlgOMQ46tjPFS5bT5vwkrCCmlNZYtpGzXbq1PxJrlIR/LFQqtuZzXJAYVdY7lJP3AXyQHNtqWKL7K98XyIub5VlGsLWxxDNngWmqtb9sIvWJwEcWRYSFB7ngtLEpWO/QR5nzE7I2Sr5gBsohf/IZhcQOu4KgnfetVknEhtUdyl2QEV+ZFRChiVfD7gd8Rk025jt6UuRDRhIwoy/m3YclzJo79GbSDOcQgYBAwCBgEDAIGgXmGgBEs5lmDmOIYBAwCZyQCmkzXYoV2awLxDiEC+QCjSeZ/SHCIbgiNYknw0MCdti6jari2kuqJc/6jRDGrg6k3RABEJuQNmCFO8D8rZMGMFYUcD4msV06fTJKe9oQsoK0QUWgnygOZgfBA+0FyUVbKDRl1oWTIMgQZBAiOp8zUjeNZGQnhAInLdVlNDWHB9cEAbNjO9aizXs0O2RVlI1QICseX9Mp7VjhDSL2v/HISm+Dhd8W+dWidvevqm9y70yJWLBELicg1CNYLYhOxPGMn1d5Yh9obb853hLsSS/y9KptLqaJYT5C6CyulwW31Bu+76rLHXlC2RJJ1R7xRWYj/3+1G6+ex/mLSHg7GrBWq38pL1O3WqG2jeeP3c3/h/0fxrQhch8Tl0KhcZ5Jl0Rq76/kPxr587jrh7RcHfSpeKKrXjDylHk9vUMNOWrli4eGJeFII6ZoT0z0dN2QTYf6RSwefeHG5f+C6aaBEhPstybh8Io7CNyVvvWj46eTTjRe9V76/tsb5XbKdvsyYh5zTVkCaxGVsVJLK7xGXVv/c4AxRaIQK3PlcX+X6CBAQg4wjhE3Ei8MVYoU+jTHEuCU+yYS02Dq88aLw+ew7cz9Z0xNrvHqxWKMcduENjyZECzTBxviAekfyjty3cu9kLI+n/Wp5q3PEaxjprl/bMtK/Rw4/CraIFe7HZhV3QGNDXb4lmTmFFdhYrlTzkY+YgUXAfZL/U4jLyA/YHBDslRBV/V9iD5Rvj555l6xsPGnzcllwbcYulhQIZxD/07no+Zkc8ynJENE8f34omf4J/jrj+ulEJfohYgX9lzHxkGTiuXBH4lbwnCtPPHvokNSR4N88M3YtgBgmkQVqLu8lZTZdVMz7bSJCSJyKsL0YBo12GBYQLQqeH/e8QMUcR34bSYgfcdImXjNjEu8iIb8lcqFt1cvnubZsCEJ/nxxDm7oiiIBx1f5YaWFRZu2kcadsPKeZ9xjPYD4TC0bmo7+ifSQjTnCeji1FfB7GM23OvMd4JSOw8BsHsQWx9GHJ9GNteVneF/R3FjfQH4iRs53yG9GiGkxmm0HAIGAQMAgYBAwC8wkBI1jMp9YwZTEIGAQWNAIVwoKuq16JD8mAib92N8PKT4g7Mi+ivAizEhTygm2cB7mtLTO43gSXPwsITF78eUnXK9ypN6Ql5CwkfRQ0uoQRGGp/7+AGPvx/slJEqkiGtECc0O1DmyFMUE5NSFBuVkez2hzXERAnrEiHDIOI0O0OMQFpQSBW7ZII4pFVvpCuJOoIyapdY7FN9wdjVXEMrS+ugcrPoh1ZoQ8RroPzQiCyjTZJrrd3BCIIrL3BvTfZYff0iFhBm6wKlDWQt+MtQ05dYsiuU88lV6tetynR6veps9PPqCEhvDP+y/GmJciz2tlzvtpdv3fL8uyBry/dt502vTfYYh22nMAPhpQf+9PJQVST33m/Fq4eFdKcFbWvnliB4MhYmP7mnmBVuMnZ8sepsJBw5DIb8vsl4rqtdsaXqj3xxRKLQYJ2O+hgE5MT80Zb3L7Hf9F29a63HfzOa93Qe4cc8dulvjeBlC87kzH6kbyd6PjB4l/6l5ydvEDK9lah9JnfqiXG9hrJz0hGfNMEIuOHlcSsjGcl/HiS652zKrlzuYgt58t1N8r/1cSKr8oJrF7Ggok5FAIwI2LFhDgC0uaM3xZpu2sFm5uKJQ5QrunJtaPfzNe7Pz/rvbF/O6s+yCjPs9T6/AE16NSrvDWRL3wxuUz59bmMjMxJ2DyWumzd2sZd+ZtHvvmIBDOn3bKzFCvKIaAOzAc4jYrqJRmCvVr6TdlIu2G99a+SDwp5iVXHSRMOSoXifnNu9VaFSNYY8HxFmKBvvUEyljnEGJgq0V+w6vmBZAhl5mrt+om5lfLPGW7TCB6B1E0/BymDdhV1n3wnqDzCWmVweeal90tmvkJ0+blcY0DuM6HPT4PBfNoN3nUSP7vJKniLHdduSbpOnbh4SngFLy7mErGjbqKstKgYfK+TWBci1Mt86TiizfqNMtAssbjwpeWWupbVKzuPyO8y7UaOeQGMa7bpFP2LsvHbjXkKAfGWafoXwgOWFTzvib/Dc7yrBDa/E/i9QzloZ21pw27Kx7345HcCizY+KxlLS543/G4gfkW1xEKPTZL53YCVVe4UjPsaRTObDQIGAYOAQcAgYBAwCExGwAgWplcYBAwCBoFTi4BeCc98zAo9bVXByyjfyTpqrg5Ay4ssK2jZB3nBCzefZNKUL92ntrrHdHfqW+6yBTZVx4UAJ+2/Hvc4+gUfthl8OBfrgpmsdjymwlWcpK0iIBwgDiERNDlHOSFkaSd8S9PmtCnlZvkxbp3oA6zkpU1pd8pNfflkG/XGlQ0EJUQG5BPkh3YZou+ly4FYMRf1OtOvAYioCli1sDIbEnA8JVW+Z5Pz1Lnvif2702QNFiSOxVohuNOBZV2YVYkn+u3G5SNO6uy+oDHX5zamWYVPnIoN6WeVHzpqfx4e9eX0bfs94YC9ZPDXhr6xdWNx+/5Cndu96pX7x93AJW+c1ByUj75Bn9ko9/5glQa77UjY2vON4rt+Iu6qnpAyvkeOycRD7zfX5Q9K4G4cFvlqtxhmLE/sUWlndIKQMhC0rX6g86pLftL6+ueW5rp3Xtv/AOML1yWQZrinwbJhUkIMGXPrXn8k3tJ45cAjB/alVg5knVQ1wQL3NawAflIyLqXKxyzf8eX+Y8kTBAup61sk/0Lif+B+ZUK7lBUGIh83VowxXKyMilhRjZi066yxZrne6zJh+tdFuBgWSxUxA7BccfflfzTxOUesZ1SbdSSKL9IoosWa/CGVlPge9zTABb6chCtVcSfb2ugMFof95glqhliZnHP2yPZt5w0/13/VwMP0qWnTDAhtiNL7JRNEnPkE908IE5WJZ8efSkYAZW4ZEfLSPwXkZShWF1qwx9riuOboGmQycy7YM98iniFUYJ0GeTtVIg4LzxD6HPM116APMa+XW/1M224n4AAt0NN2lA2LCwLEV0v4eyPjRvExyi84DZ+Ctp4TGFzXthwJT++6jiMiRKMfqnYJrr1ExmdDKLEqxMWT67qWH3cdTxrelv0J2ZYNA9+SaS0VEzsLeR6OiHcoOwiCDjGEIlaItkQ7nsDb2rqL/sEcfMsUFf6E7KPfY6nD74FoDErWQlL5vFQtaLq2NuP3RZdk6oD4wZyKuyjEi2rjniJ9TfI/S8YyZ2/J6uZ0FbDm7my+rwAAIABJREFUpE+ZixgEDAIGAYOAQcAgMH8RMILF/G0bUzKDgEHgzEKAl1DmZF6eIUZZrceKUIgnSHhtTQCJghWBJqYhrnnZZZv2da1X4B0XATRf4C8R7oGshNQWA2DSJRkCv1wUgMDX5BIYaIsGS86Vy5yU2A2RQFJqM/CHREBgIFFWVuTrwNuIE5o4w4UHbUj7ImJwLvWBjCCzAhPSjL4AwYHIwTEcD6lRLujM2arfUrnNx1HswRVLGMgg2iQKcpyyssPXOA8Nvs79qSXBtmXNfZgSMjtRUO7+nBXP51X8oucSq5xdqaUSiVf8LpUSokW9M6wa3AmucqK9QpJbT6UvsS53N/cO2Q/vXf3Xh/JJQu9WT/R1rgtjThDqG8oOw6VIROLLNZ+R/Pyj/mVd4r5KB3yPSzn21gW5Pzo7vz/Z7g2rc6wDqs9dps5OPaO2jE5chD7kt76zsWngxT+46lM7Hv7+qxAX6LeMs82SIe0+WllEXFwNu40tI27jm3an1ygRK6rVAjwRZCDeIInL+zPHa9GSmBPcr/wiMcH7TYUwkYhbuQt1AOyymyB+IKzgRgWrjeFqYgUug57xr0k+E5yvPpX/+PJd4RowG3ettMQ+7LzD/Y4EQ8/JIPSiIOWuLNZu9keV4CeMv7394fR5K3J2nPEtlip+JPysSHZ5z41dPEGwSPq53KHkkoRnu8wPWtSs3roz38p8oF1ZfV2+0/aISG+qcgmeNbjpukUy1iy4DCoP9D3plNm4PCoJETN1+UT/jck5zJveHLqJ0uMCoQqhAiEMsfFDU0BKPwE3BiW4sAK+SzJ9U6/An3mLnLgj9XOGO1C+L0j+nmTcXf2Z5EoR7FdlG3XD0uL5kqXFvHxOiGumaqhFqruoDZ48x70wCDL5omd7ftgqEkQhHnOG5RmfkWUJybqE68iBgQSvEC028rXnxmN2xlI242NABI8u+aV1MF8Qoc6y+iWcPW17PNYyWnTDCpZA17hnqkwICTzfEVxx9cTvFOY5nt+RK6rpxlcNQU7/TsBKA0ENAYRYNSjgWFNhvVmZcNXH7w7m6i657uHTVcCqUjezySBgEDAIGAQMAgaBBYSAESwWUGOaqhgEDAKnJQKaNODFGgIeQpqXWMhsiC8Ibl5KiXHAd150Ibh42eWTVdUQEbws65X3kC0QV9on87wkJo6htbQAg0ADDuCDuANm1BlykRd2iC9IfO1n/BhuddyngDltSptArkJMUibKS7n5nzaGREOggGCivAgTnENdOJ5V0BCtJAhhiAkIEup/qut43CDN1wtUuIOif2H1coMA32Gp4GkhyFNijxAJFoutnh3iDiorsStYdf86IcyTXujsljAFbYdjLX39TmPipfSKS6VDTDJ1gVw/a2xH7zlqm/2COl8LWxEsffH26z6z/uMrP73hj19U/1jLg1J0KCInZBiJeYCy6qTHA77SqUeXZFbTe0JUwQwyf+SkHMNCvl/X6g+/haOuCp5Qvel2tTN7rhLrgPGL5cPE8jp75KpcOvVTCaC9Y+juZuJBcF0SRClk3DckjwfB8C1H9SQ61DMNF6gH2ibH2ZZ7Dzih/6+e5dLXKR/ju1JsZTwxpyHUYdHBfBgliV/RPei1bjpSbI9L0O1KlJlLkXqwPoCA1jFdxuvEF8HCyYSpxa3WwEUXO0+vEKECkntCutZ5MBIrOqxelZZ4vloYsaUNJQ+JHPqkuNnK5VQcgUhi+0ocC2dQ3H49rXZkzs2IoDIuVg3Gmpvvbb/+xssGNj986eCTmx0hYT95+72V/WPCvF3pR7+yfGX/a6ur50t1Z3X9RPOPowczLyFafFLybZJxO1cpFE1xmyl3zZQA1qvFOT7qMyJcHK9ooXHkecpYwMKA+uPWaSqxAizov1gisBCAPggJjEAGoTwfn6O0NQI2FiGMQ1b317LY+d+yD/EKV2DfkT7fO0/rVKtjhbZteZ4vZk3i2Uk6SyzmWhkJRXFYrCyaRMhod0SqKPh+WMz5IcG2LWXFRaDwsbLw/CKCR724iWogxoXEvtCuI8v74Gz7O32NZzXPAn6fTYhrVHYxArV3SWaM7ZbMvKTja83onjOwsOL3A/Mj8WwY8wRbx1UYwkVlYkwgrtxZKsdk1XxGpTIHGQQMAgYBg4BBwCBgEDhxCBjB4sRha65sEDAIGARmggAvvDrmASs4IR4hsnn5hGzkZRhCglWfvOSyUpRtWFxAwHC+DjDNdoQMXoghtiHCCcq9kAIuQyJBqiEGjLvIke9shzzlxRsiDjIiWjl5kiwrKtsaEkS7hWIfZBzPXMrOanJECAhM2otVkBANHMPKSMpO20Fu0Ob0D+pC3ainFmQi11+nqH6V9V2o/+tV2vQpcSsTxsRl0EtCUV88GrriJD1z5PXuPYOvce9bvdbaDYkdE2Oe4kChfuU2d3VTd6LtnOF0emU1saLj8EDWLfrFIB+7s9npxxvTBypBFHdKuPd4SASUWqvwte905gPIyl+jz5ddB1cxEJma6B/LvU08HnHQayP3MBCz9Cvmmm43DLob/cyHltq9ap29W7XGeicIFsTXOD+95VLHDy65pf1zBxP/EglnEcmdvzXqs6wgph7vlExfvlDcYmFZotZmmK4mp5sOfe8r4o7qqcebX7El5WezW3/9iqqWYYIB94HkYy4cFyyKYbxVcE/kAhlOk72fsfKcoLScV6yMWSH1Z2wxDpf4yrl2e7BhWZM1NOArG0uaCelSZ4sMaFeJdYoAOu5F5Sdy0FYRqnY2BNmhlYWeHw4nUx8QkebVnByz82plYmfqrPRz6rkxpu6Xkwg06Rcazl/xk8VvumeFn+OCzGnaOq58BT0nzYYs19YoiDQQklybuA03V22Ao8F47yjdgzm0ZvDhGudP2KzdPM3CxRPtzVzJ/BhZMmFtcRyWFsyjPAsR7xCezpVM7BJioFRLkP3cm1XwiGXgp2OBnA7uFXVfwfqIeYC2ZPxVS5hMQWbz++C/SrjPpFlP2jE1hLlQLC/EoiKQsBW2WFTYOVEhchLHYkxiVzSKlUROrCyyRd+3xDWULR6fLMcK7ZhtZfgaBKpBBroE4FaiXYSLRKx4SXJBBhvYHav1DH0GkZm4EZD/uNirlpgXEcJw1YaFF/ebzXieDfZcV7uI5D4E8kaoHZ8vyy52q3yPYqLJPLgVEXs2NzLHGgQMAgYBg4BBwCBgEDjRCBjB4kQjbK5vEDAIGASmR0CT25B/rNKDdIBgQ3jgO6SlDkAL8QgBBeHAClqINVZU8p05nWDU5Iigk8y1cae0kAIvU39N0rD6lXpH9ZSs3XbwfaarfKdvodkfwf0pG2KTXvHMUnXaBcECkYky094Qu5AFkKfaLzXEnQ6wDvEACTHenqVzKdWJIj5mX+MFckaFdQV9CCuEZiHFIT2vS6nsYyJa+KPiMuhS58lusayIn22/mI9bhd7Asw54nrP0YKxt0+H6lqZMLLEkVvAdESby2VQCITJKsaJXXL9931dkW8eh9JKHuuuWu7GweEXRilXGYIB0rubHXF+KPoNQQVwH+lclZQ8Zj4/7r0rGDdQEf+WlFdYFIaywWuiTOjYnw/ztS7z+mxv9XKy7MIm3l3nEP//KugfecIF67qEv3CMk4Msrz+nzzGE/kgz5i2/5Pxxym1/5QNur1NdWvn9SD7lscLN658Fv/Xo8KHT+yYufHluSPzRUf6s6IkJINdGCvg6GE+pQCBKJlJPBfZPyJNZuzC5o6wfIeuZG4hdAxI8n3D/JP5rYhtReU1TxywfDxlZXFd+5L5hc7wvsbaLwxIcEI8YlVlK/I5k5uiijcDQRFg5K0PL20LIhKCPBQrv9urB+8yTBggJIPI/m7658T9PlQY7r6fhFtKmeC6irFjFm6+IPvHhuICIx5yBOfXhSIxztP7gTwq89fvVRlo6XVLVFdAjLRQv5XuXW45u8kkso6q1d7Mx2buM8ngW4KVtfqiv/4yaJFeXVEn2Evqr7LTgh3jF3z6s0zQr7kHgEpbZmnJPfLPnsKpXApd31kgnCHQV4Pl0sLcQywhMrCZXNea7tWG48dAYTElDbD8M2yUXpABLdwha3UWFSYlSESr6La6is7BOLJ1UQa4x9thX228rekQv93XKIdqE27diqcMlEP6VDb5CMIKwt3Kr1GcYW/YrFB8c7rmbSJ/XvSX4jItJ9XzK/I++pOBlLDJ4N/KZMEMdGPieMuencVM2kMOYYg4BBwCBgEDAIGAQMAseKgBEsjhU5c55BwCBgEJgbBDTxDsnFKmoIShIvj7xk6pgMV8p3CKc9kjmWF2BWGuv9kEyQMrxAQ0JA7PHJdXi5Fs0ilMXOJyWOw9wgM/VVyle+gqEOnFlO8M2W8JqrcmvxhDJqVwsQkqzahdyAgKZ9EDN0EFf+18fTbhAb2q0XdauMU0FZT1X95gqneXkdsUAYL1dJvGirt0ZXyAr8xRIg215j71naE7Y3yyr7fBDae8+zn9+7zOpebGWDweGxVOtQvi430pRaOdyaXpWPx2MtAyM533GGsqloZbNqGM680N439GI2nahLZfIvLT/c//Tw+tZ2OQZXNOWCBWNaC1oICvSH8qQJWvpORDrVABQSGlKW/la1zwgxFeDXXvbfIRf9xQvhhs+nfP9v1ri7rnqhcN6Eyz4yfIO6rvWBKy70dq17KbFchIADEPhKRAauTe4TawvIucb+eFu+L972se8u+eU34haqPF00/LT60+2fVE3eUPuK7P63yefOWADnqJ6X8yFcvdI1o9OkXYLmu7p7vTC22Qvd8dXMCTsrg9+X4OWuGvDaVVvssPhjihYLf00ycyLWTNslR6RkyaqC37+0B8Q2hP07RIh6vaOC+BeLuHifmC52tqp94Qq1ztr1fFHFHkuoPIKitujqkfMGlxaP5PJWrBgoi7HK6vUodkRSytfkDKil8X0KAegoG48bKZkQkos3LM/krjyYWpIRxpNYG2ymHSkf5aXNo++ywlwLlpPKd3QDC70nJa6BpRaJa0Ni4gKqMq2WDcQ+0S6+XpDvUwllNcowfh/muWlJ4IqL6HkzEt2w1KhlZVHFn7+2NET87ZRMrArc9EAkI2DUSuDB2GDs0U/KrfamquN83KcFQywtvltq67+pUdCPyXYsSx6UjJXfsbb1ycQhWgRQKMpMbFuHbdvht9ByPxDzJLFqk983RctWOfmZo0TYkCUaeGoLAlEqhiQId6Lo+Y78CmL1xrB4jULPyEpmnuJ3Fwkrjkn1qWLxQV9j/GMZqRchIBhXS8wDWDgwtx6X5dIxAM39EFQZi3xeLfnPJb9OMv3iS6V6YInEsczjp0M/OAYozCkGAYOAQcAgYBAwCJyOCBjB4nRsNVNmg4BBYKEhoElE5mTECF6CeSFGsNAugCCUWPYLmQ05qYO4QuzxwklsBFb18skLOBmynJX5rOZH2MiW3EPNlkiar3iDm7ai0BYVlPVkEwPV8NFlQ0DRbnNoO72ym5XvkGPs00HTISdpV7L2rz3u/mkBiU3ztT9VK1fSVd5aIbOvHVX1a8SKIrMzWLt4NKxPiGCx7ZXOw49fHG49EssXUgXPbezxmzt6nGbLz9jbRazAIkMNtDQw/sgqkS+MSQ84nKlLbkuP5R4RS4sdCS/fNWbXDYr7J2I/4J5HJ1ZCsyL+ackHGL+SKwUHVuXTlyCaL6pSAchprhu5CdHuoKpVlFXWQgQjahSW+v2dh8LlX+y09mx6QZ03QQgZ8+vVbr/z/COxJ/64Q+V+7wePXf78L13+2ASrBxEaPBF7hteN7dx5Q9/Pvr6j7qxr5LrMTePp5gPfVBvGXsyLFUaiUYJ9u4EHkQZpjFUEK3/3i3BRLLe2OK/uydye3Pqdw17zAbF2QGgQAtJRuKo6mF+lmtwj2sTk87KLlfUEBoeFzBBom1gV8h3xkHGIYPFBySukDK/0ZNeATL3SvpPgSQoPKiLFgaXWod0ijkBwQ/YSbyZy8aJXqP/d1jjjGbywangTwoQr+kWz26+WSQDuo4KFLPzmIAnYPZTouLo79A61yjXrZeW3MKoNrASXRqad24RQxRWZthqjzFMGxp5U8KMbaBuEcNoWMhvxm9X35Yl9N0rmvuDGHATReiwEpn5mVVr71CjehM1a9JrtuRwP7vjd4hq0A32uVkL8R8Qi/tN9knmmHgu2M6nTyT6GeYL4BQhVYEJ7VyPUvyrbPyH5S6V4FhPG8Mku9HT3E+EAQSGKQSO2EwUxtOgVYaLzqGmidUS8zsmcLMG1ZYdlh8tjjiWBti0/VKEXc9muinL8qJx8qOiFBRlbejxFVg9cf7oylPZzHkOY4xEB/rDsPOZZxhJWOsQMQTBDWGEcnQp8gYfxyDxCuZgXEan02GacoyQzjyHs8XksY36G0JnDDAIGAYOAQcAgYBAwCMwcASNYzBwrc6RBwCBgEDguBHiRrpKwfNDkNrs5CLKaldasFtUWGLil4cUTgpIXS8gWXoa1i4Gb5DvWFbwU6+DNkDe8OGsf9dG7fbQS0bJOO9GiFn4ljDAh0fjxOVPy4bjatPzkKuWLyiDlggjTZIX2VQ9RoMlm9tM2WmjSMSt0HU4HP+pzhuN8uZAQ7rTDoqSVvyavklcVwjiWFt0SbDudtLJ7r3A2/+CN9o+77cPenrGxeCHXlFh0JGxYvHvF0gtziYi4Hk+uRHz1XCdWN5rbE9hWzvb9B72Y87O+Rc3Fmz70mJ/8ThySCP/yCBMREV9KiJba5VklNJrcpX9ggRGt6C9LEFQE2I2sFbBQmA7bkqVF5nDQcfhR74rhwbDl53LO6yvP2xOuVA+mL3j9a3Ob3yrxKfb83da3jiII6OMEO+ax1M66dRu70p1XSkyHCWIFxz3ZtEltGH0pccnQFiVBtyHycX33z5K7JBN7giDIhxAt5DP4wkfeau3IPlS3NrU9JvEgBiVHOIlwoYa8FvXQ0A1qfXobA5+5EREHUppg41qsAEfKgfjL6vtOyZDzV+JOSlxCKREkxPcXsE1MEqPi2Qucbd+V+BaPx5T3pOyF2IMYDsrd6QgGgWDBqu27S/f5mC1TbaM7oFYkdqutI1ermKwAd6WUdVLnpEzpllu30lWZc5ywEBMW1BW2tVt87udsS8UlwHuXEKzMDeCJ0KLnhkltOY37FoKs0yeZfz4tmZXf/1hWS54vpF+SjBhDzAsEVPrVbH3ba0KX6832XF2k6JlYaWVRxbKi/HjqQJ8gbkutGA76eKyO7pf8A8n0E9wiTTs+yvCaz1/BTsdKwiXQ45L5HXBLlUIjaGJNc69gS7+ticF8cg9ELIqiBM6WjjYorqH6LbFgC7zQc+IqIQOkXrZbxSIGpfzosjzf9/e5LuNKrCu8YGcQBliVIOJF1mGSZiomRPOaZBaPMEbeXoEpkwe/yxhbxKzQVpNDJ7p/TdE+keWNtC/tjHiCtQXurJhLWByj3aixWEa7nqzSVcwmg4BBwCBgEDAIGAQMAicXASNYnFy8zd0MAgYBg0A1BLRgwYsl5BwCA2QRGZcVuAqBgMNFDNYUCBEQ3hCckFBsQ8TgZZQgkLyQQn5DxjHPQ0Sw0pIX7egFWkj0UxWM+oT1gJJgcNKFihlWCNxpC1ZmksqtLrR1iF6FCZEwThwZy4oZIjyHh5UId2eN3bU4E6YvS4m/JyGPD621d48usvoOdgWr999g37v77NyL6UK3taqnYdGre2MtwyOplHuktREyaNxhv4VZk+M4yWzhUQlW/TMrtLYGjvO4CBjFm3513DJBB1SP3EZVJMa+tqgq3wV5BtHGOVhmvEpyufhJoFfGvLZCmhFCEPD/8V9tA93BkscyKk18h0mCxd78OvVKcYne4Gdu9Sz7W3VBbqcQYl4ZeU8fhkBeJ2LFRF9QpVKMug19aX+svd4fFRV1Ak+Kq5U/k4zQQsBssEEgcFvd3uX5ILVxU8ND8fIg1tkALh91Y8Xwolj30+ISipg+ELWRkCJl02MPAQhhl7nzf2hAxMmMGgnr1YvBenW/N3lh/piq/9aD3tV3nOu80HO183DUVrX8/sv9PBEtmIu/LRnLmg/RACvie8VW5Xl1ILde7haqlAgZdTLM221pv9C9wrHDoiwRb5IV4atFe2V1fCYI7LxEDN4nbmxysjocchWRsyirwWdNrpcsaBCzeY4w//xM8muqdIo/KeHOcwQyH+wn+bevcp7eRHXJ2k3fFIe+vKtKjIuZzOX6XowR+hl9p5ZYQT0YE1gj/btkxCwI2pptOaOCz8+D6B/8BsAKCGHtryS/Q/LRgTIxIQxiyYW4QXvPd4Ec64hDEkz7qMAfSkBtS/UEtoqJn6cGcQ81JG6jjkjnyYmFxSKZflsk7kVMWeGIjKtu+b9fonIfCpSvA2AHs7Cu4PmNKIY1ErHCmB/LE0Ioid9jV0hG8EUsmqkgUqV55maTjH9f5kF+UyJc8FxAvEW0YZsOPK4FnLm5qbmKQcAgYBAwCBgEDAIGgeNAwAgWxwGeOdUgYBAwCMwRAnqltF5pzwsk8SlYxcc2Xiz1SlVefCEC8TcOSYPvbU0OQr7gzwS/7bxUk1lJyDVweaFjIkBaFEor/1EuZkIMzVFVz7zLlPDFkEYH1tb+orX1DKBokaJ825kH1hQ1LlnQVB6hzZbKP8uxJNj8rMnd0k0ccRW0JK8STdkw2SCxC4TxamhsUKN9g37zvsxAMh47kmvMFpKLeppbOmWEdsmdDjcOjfXnk/F0Ie4mZHDZDLBEvvijpqHRfxDB4vnBlvqR5oHRwZ1nLS8vF+QbMU4QFxEgyxMkGeOe32zl7jroKwgZnZLfWjqBMa5FCsa8dgkyqzH+9jfd5a+769MDEoB6f8LKD+TDxIQ4AC9lLlAH8mvULmfnqk2F7Z/KWbHfl3sdhhArEfm0B/MUc8+5kxst9NsLvY8uzh++QOJWrMZNUlmK3GdJwpUVgWG/kEknnxX3WYHEg1gj1hR1Dc7Q+mWJvZEbqPIkMSz2isXFLrHY2FyvModeM7JFffSeSKylLIhIb5N8s2RiHIwnLCwGwha11Z/sVavN6t/eG7TH/rbwUXW9+/PRa97w8EzIR9oJ11FiMSO0qfwlcA1lD6teEWeSMuU2CC/cJM2TttVqx3GtRMIeSqsgIcvBZV53ugSTHvluFT0rVSh4tCvushAsfHGNkzlG0YJYJRD2PCu+VvqE5IdcLU8IOgQLhpQl0S9n6iqGfk2/c6aKQ1Fxv2n/rRG3gv7PKvFOyTz3xkWoKhfEMgbLEhYBIGix6n1W42LaQs6vA7SlBaQ0OP2K5J9UKSLzy22SmX8QCBE4EOXmHTZlbqEk/kTgi2ghUbVlWFmBuH5SA45YcsVcq1mcrqVF1KgP/TAT2lZWBIshiVsxJKLFS2Jz0S3nDch5kPSTxIoaVjzMZ8wjLAhBwH215Mm+446C+yPJzL24XQLHciH3lPaQkpUH9c5LPSkb9TrW5+MprYu5uUHAIGAQMAgYBAwCCx8BI1gs/DY2NTQIGARODwS0aMEnhCukAWID5Bim+qx8JLFCGMGB4yCv8FWNsMHKPl5EeQFlpSmuCSJyq/Q/hAUr/SAe2cbqZT69hWhtMU+bvHzlqg4Orou6kAKinwz49cpqTbgwZsiQbzqweTSm6N+l8TJbca7hQLD8XHEHZDdbg30iWKztDpcmloUHB35l5LuLLh94NO32FPMjra25gdYGd7ipbpPc57G60ew2iVGxQm62UnjpnOt533aL3l+P1qdeGqtPRe6NPnjVf1WSRNqFSzVSGBcj1EXXS+NLfREzmSt0KrewgHyEmNZizqza5UCwDLHhybiVZyX+r1aeTGyGbcnValXQfeOKYi9xNlhN/IhkxBfKAVFKLAfEjAlJ4lU8u6jQt7nJG35QxIXrZCfuVaol3FzdJaRjbuXenj6v07UvqHv8+j25s6JYEOWp3hnJ7cieO1TnjHR1xA9u/8P8bYUVxT5ECgJrY1UBMY9gMUGsEFFKOs7R5rjbe4Oqs8aKY2HduEWLBNS+qz9sHZDb5b9ceL+M249Oi2OZa6jNKrS+LFY1H2hwRtS65IuqmF+ssv4i1Wr54irKUq22o2KWWFbY1tpULNYo9ji+rARPyv06cgWiifurA8cSkt0e9fyAVeEQp56IFoVjFC2wOKHP3CuZiiNWVAoW1JH4HpCvCE775JzItVityle4pNHPs2mxOsYD6NO8wyyV/IrS91+b4lq4Rvu/khEqeJ7qQMvHePvT5jRtaUF7IFQh2jBPVUvgp59LzB1Yds47MrtMtMDSQoS8MOYHkbWF6MJFW8QK6irjNeyQmZ/5dJ8fBPwe2iGfBxzbHskXvGkC2E+Ch8UhLADhtxWCMGnCPFLaRj/DnR1u6fg9lpuvotiJdlF12owQU1CDgEHAIGAQMAgYBOYtAkawmLdNYwpmEDAInCkIaFdGZTEYICZ5Ad8imZdvVgd3SoasYpUtK5B5cdarXnn5ZhtBfhE2IHNY3UvwWl6010hG5IB84KWblX9R3NfS9c2q/pPQ2aq4rJp3K1hPAgzHcwstUnAN+i+CHNsYKzpYOdvp95Dt2mc/OEdBzGWMIQzNhITjOqIuuK4E144CHweh7aRUJrM8e/DQWUde6l7ae7C7OOYsD1qt1GBLw+J8Iha3g6BFiLKkuHtaK66ghkSweNpz3c3FmIuLn0hcgcyuAoK2CoHogoQtT6+UfyCOIVrLkxYiCFCtE6KkdvuCCFC+r8pta2+SmBcSW2PwkB+63xRC/01ihcBc8vKNvEVqcXy/GrAbk2vCQ58Qj/Ln2yosCrH9+JqRw86hcDEr3z8kGZF1QpIA47c90nLF3b/SfWdvR76HWAK4roEYv77swMgiSWJ+/KVgml655/DnDy9pTXnp0Usb3UHVHjskVh6rxw8f9RuSmSB9ccwqfqElU8yucPsQZ5knET2YA5kfcac3IYlgIYutbbcnXBSKlQWYTnCUxvb7AAAgAElEQVS/1Re25aTurJimP81mzBZDP7FZVnXT994dU0FqqXtYeentaudYu2qXX+DJhKuEbZUSCCKWGovF7OZUMi5eoWSzF6z3wsD3/LA37Uit5Gs2p/aJaIG7KbDB0mI2wYLH611yD4WlAf2KQNy0EWJOeeqUf1iR/2XJ9EsCmGsRvRLG8f/FtVMolhUnWrDg/YVnGSYxjHfKjlVIZYKkRzRDdKOekPCseJ/JHFCzjvNxB4JRDesA2gLynPb+nGR8nn2gSh3AkkDRHIe495+SER3nHVZlogVCRLbo+TGxmsBiwJE5nt9FMqwtTywrsjKgh0UBzDiWPSJS4LDEs/Dl/JlaC2lhjLmDZwLPFQRk5uTKxPzwGcn7S8ctyH42H/u+KZNBwCBgEDAIGAQMAgsTASNYLMx2NbUyCBgETl8EtDsNXrohurTFBN95WT5bMi/mrISE5ITgg5SDpOyUzHkEe9SuoxAlIHaY77dK5gWfVdm4neEFGwKHVeh5IXJn4urk9EXWlHxeIzCFy6dyCwFII/o9Ah0EOmOCzP+462CfFuro3xD4rCaHtIOkwhXaTOK3cE9W5y+R+AbpI2HLSFwVugLfSu33lufflPn+noElqbyqb/deOnvFpmwqIQRfOFw3mh8qJGKRX3PbD/6vxKp4Rlb54raNsuRriBUcTvlY/YzF1HUVDfVu+R+f+6xwL09gAWNfHnQBaysSAgljHfL9eAjHvNS/SwQLCPsJ/tqxcpB4EeqhlASVDsfc83Jd74iF/iPbgw27CirGfHSeZO2qqrzcWySuxegjLVcO/bDjjblLhp6Kgv5K/oXkcyRrwcb1HdstxGNpL+aqbDrxibG6pDSwr1pjvSKWEJ98YgpDOzycW9lxdfJzZ4lFzCtiqgiWzJkbJx1c2pBX8e/tCtZ+83OF3xHKV91aeZyIFdSbdsmLiDNjwaJkZTHkZJPPh7b6p9AOPuoFaZUXj09iUaGaLE8VxfF+PG4rqWa6KRn6cdcZS8Wdegm0vaJoqYa0CBpCtIpHrFhqLFtoi8X8ncMj2byIFlGbzsL3/qTql3zaM/8zPj5Swun8igMZS/9L8nck06Z3Sgb4KZ8VIlr4iBaIF7VwP47t9HsIdfo9QhQr3d9Y43oIFYguCPgIfgTXPhFlOo7qzN2pUwRexqqGxQzfl8xchJhXPjbpB8yhWCIxVhAP+S2BoMU8Mu8wK4kWkcUa7SrWFrovRwKzFHkQKdCyFS6hinmidJeEvmqIVxF7eJYgioMLgh5z7X8vYVN5CSzZfl0yzyC+417reObduesU5koGAYOAQcAgYBAwCBgETlMEjGBxmjacKbZBwCCwoBHgRReikRdlXsj5vkMyL9CsIoVgwgUL/+O3G3IS39ysJIa8ZVUk2yGVeHHG/znEE6uYETPYz4s4ogUrdSOXMsS0ECa3psuPBY24qdx8Q0BbU2iBQrvwYCxAtrHKFTHuaODVoyIcfZzvrIblf0h2SCz6OoQTYyEiWomDXcvSQgfclsPwUQ6BO2AF4TMSa6FYsOIJWQ2/L50eXj64uG7poTXNa3o6Ws4Ta4qs5JFcMt4eOLYv3++WzydErGC1MuMzJwT2BJJX7lOOOWMeYhBxgwQpDEGMlYJe5VtOGrINDHB39LvlFyp9Z+4g6PTxBnylXMTyKHc7Fd1i8/Cr1Jrk9kg82Jpao5YX+1SrP3xJQuUf6LT3tkicj0Yh+3UQ2vIi/lD+2S05/5n1Hw//6KXPUO97JNN+vyWZoM9XSaByNVaXULlUQkn8CnVgxdFwCriCklgWanVyh1qT2q52Z9EjjiYpZ/1oWP/ZvcHKz0mw9KEma4iV5TXFCtxBZcPUZ187drcr5zF/lieE4T+STKBm5tBJGFQcP+lfb+hcteTIM1Y+Ed/V35YaSDuZljViYUEXdvxlqtkNVT2iRMKxi8rbEIs58YBCSbFsW+Vijpt306GbiDtidhHzEwnXzeWKy8Ow2C+iRr9YWLBa/JiJ0ZKlRSSmSSZYNbGTqiUsGBAJ6J+MK/rilPcVseKYy1WjDHpOwOIQYYvn3/skMwaqpf8jG/+51G6Q9aPVxArBsFwQLXepxjXHx5zgPF1zz+v9pbZmPkAgZF4iPgyBuEl6AYOuQ6d8YV5hHsKNFufNS9FCyoV7NPoagpTEtgh1zB8przhXe7kXMlZmuiiDPkH/YtKhf62SjKg3KR5PCTAsK8CM5w+WsIWFLIzN645uCmcQMAgYBAwCBgGDwIJBwAgWC6YpTUUMAgaBBYYAL9aQtJCyJFbtQZjhWxqm8wnJrDCHEISIhXCCYIPI0XEq2AZZC0EB4cD/EG+sSuW6EJ5cVxO+Y7NwmXNawi2rKCEz1guZACa40FgsHwRfzZVWWEL0Qogh6pDA8yVWI5+WFT59Cw1hpONRaHdJ1Ib2YR/kKSvx6c8QrrDWV0qGtGIlLL9vEN9Y5c85kG0Idl2l7TksOmqIFtyXa3OtuyQX4kHBcwJ/Q8rO7K2LDe9uzA6vGnSTzUfaGjsk9sCYuIIaFZHiaXH91Cyl2yk2HAiK9CEEwt5KsaJGszAeIcgQOLCK0gm3NpS9XEwEA8Yw9cTCqjJhsYD7nlmT7BUXAjfK86DkST7bJQB2ZPEw4DSoISetmvzMe4X4H5aYD8w1BPmtlnBJBzYcEzbdOMjYGhy6u5l2hOz7quD3w1wq/hvSQJ1iYaEeu/K8ccGCCzoChcSpUMvcfZnd6uwJrqqkVd3hsKllZ7D2wY3O09eIS68axVAHcirxH18u3FIvwdTPEkuScsw5Bwsb+gLzLX1hVnNA/lZlHb7zTjsfj3t7Vy17zvITPz7SlL3RceMNi9PdKllYqtpTjkqLhUVCBUHKdpviMccLxEFVPO44ntw6q7wm8WJ2zsiYOLUJw4TnBR0SnPsZy44Nj2UKcyIIlIhs+hZ9DMEI8hVMta9+jR9ucAg4TN9GGGdczrnAPUXQY55lzM2vkvwaybgwqiVWfFP2fUkyz1Cei2OfOrRZffL2CfFctFBBPRhH4KljOETu20p53hH1tTr0dNtLVjU8+26XjPgLnrQpSbuS05fBggUXUrh12yrtomPTVL3NFNYd0xXruPeXRLtAhAvdH7W4Ne6abBbWSPQF+j8iN3MYzxaEb54l1RLij3a5BbZZI1Ycd5OaCxgEDAIGAYOAQcAgYBCIfqCbZBAwCBgEDALzCwFesnnx1sFBIQz1CkII9s5ShpBkue6rJWNRAYmkE0IE5CeZVdqsaOYFHJcxEA+4l4GogaSA0OFcCAxc5tQicucXSlOURsgV6gKGiDdgBtmKUBOtspf9YAHpBTHdLP9rYQjiAYKSVcS4E0EQukr2gyMYagsViFVXiImZ+sI+bbA72QUti92ib02/1ISTDqwLcYw4waeOSUEbgj9tAXkJ4Uxf5xhIfs7V1km0I9elffmMXCXVcA/F+az6p62JF9CWdVPLEkFucZM1eO4V9gMdQ53xNYeXNJ2TT8abA9sWoSHsCi27T4h27tslGf/vjLHRWm6gxL1QOdShWFxQF+pI30OQ0QlB4lLJ+EanrtSfOlB/rAIQZMrTHfIPpDNucBjXsyJcKyw/ohXnMiP0i2VDn3yyEns8PZfZpM6v26JEyFGPps9RKe9ZtStcc63EhOgR6wrGW2XC6oP5BgF1Qkr8iyru/+Pm0dYjI7ihee9gc/0+yenuZW0d+1ZN1GQsKRFCSYfP1Dg5PeFf8oZfiX33ZnELlawhWHxPzvrfPcHitvv9azqkbuBaLSGC4aqLvjAjHBEq5NjIbdnikedXenb88paxbuuCneri/YvObfj59VereqtPhYFMw1ZcJUJfJcWaxI25WVc8X3nKbnQcR4Jvh75ERfGKnpVy3WC1TMtNrmMftm17h2Nb2T6JxTIyRnc+/lQSLbgYrsd4PtxW46p/Ltt55mAlQ0JkOpFz4DiWch/6HuOcuZx5/eoaZSQmCn0M4fKx7uK5I1/u/9fKttOCKNsZ74iFbAMDPvUcQ91oy2ktSo6/FU7OFaStC/I8wz0kz0VcfeEy6y9L9awsBNZJYM5vDdpaW2TOiVg21zUuEyVmNFYr7k87a6ECIQyBjPYnFpB2U1dZ5KdkA3Msx7GYhN8Xx3LvuYbCXM8gYBAwCBgEDAIGAYPAaY+AESxO+yY0FTAIGAQWKAK89LLaE2KAl2DEC8QFSEv+v1AycziBRBErdBBu9rPKD3IBQgJih6CjEKG4k2KlIG4e2K5XorMPwo7rQ+RmhCzLzjA48byAXwgYSCbEGFhg6lAuUkAca8sTCGWIXkhItkFyQ1RsLlUEYlgT31xzk2RWUIIvRBlEBveJxAu5LyvFISsQOfaZlZXH1B3An1QpVDAGaE8wZyUwRD7kECvfIZZoG4QFxCRWv+IKCqKfFfy4gGH8QK7ixoO2Y7xwDRJtRvtiaUEg7nKSifMYb8QuaBcye5MIEa+SQNr+cld0iUQxsbd98aVe0l5mB+FD4vapXsQKgjkjbhDrYJdkxlhNsaJUhsoPxiFEItfAl7xe8UwfY9xSfk2mIrBBJL7sD+nlq+G+hLFNOcatAiSmQLSifJZxBcAF8pcx8IjkN5cXel9urRr02sS1Ub/qFeOS/W6HGs7XX7jCOti1P9L6JiUsVhAruOYEYu/vtr7V+g9Z1d8yMDKyuuvQHftXdIwNtDb8icSxqArXpmefV+fkDqQluPbIPzR/DMJ5PL0YrF80HDb6klXcKkjHGudXIeSZD0Oxqhj6YuHWwuP+pavFumKS9UjpYhC1zI2ZmcSvKIkVEJ3MF7TBZU7o3ZwqDK/PWulWCWyi2oaHlds6Ksx4n6qLJ1RL3BXxwnft0EsGQTwXt23nqFwX5sT3vqgVToPlWOLpJtwnbqJ6i8XQLXpeY3NDcmCuBIsy6Hhu4F4Q9ze4U6oG/r/J9l+WzBhBMcJd4YkSLRATGN+MRdr4Wsk8495VtVMo9VHZ3iW5yQsTT/d6a4ceHns/jc/Yob/pMcTpzCFcn0R7UVfam23MN/RT2pLzirJ6X8dLqHrr08xlFKIUOH6jVFfmib+tgSniFeL9JyUzrzKH8rxDvFhI5DzPFZ4huKbjNwL1vElyLbGC+nMMzxss2hgLBNpeSJjU6BJms0HAIGAQMAgYBAwCBoETj4ARLE48xuYOBgGDgEHgWBHQL764ddGr+CAhIRsgDCBweMmGSIQ8gkz4qWTOg8hk5TVkD7748T3Od86BSeSlnNWkZF7IIRAhZyDrefEuCpFbrCByj7UeJ+M83JdQjw9Lhu6DjAITMECY4BORplM58azyC1hXRBYlkiEkLy4Vku+QVZCNkBaQV+DFsexDrIBA5n4IRZDM4P15yZDK/G9SFQSqBNXW5LsmRfVKZ/ok7cV28ESUgJzHYoA+St+l/7MPtyW4qNGCEm0B2U+bcw5txG8dyH/aB+ITsh8ykn6uV1JHY60UvwKRBAGEIMwyvsKuhJXLptxM07Km3QeteG60GHdekF7m+U7k+gmyG0IfoYGV58ciVnB7iFXGIWO63D0L9UVoAy/qol3FQZhVI5SpC6IF9Rx++DJbu76JPkW4mFK0wPKjzMqCa2GttVmsK7rkE7dAlGc8jfiNKh8mJdCFp7YlV6tsIaW8vNtZfkzpO+Iqbofwie+VCwCIFbKNMXvZQEvDFWJZ0eMW/RERKyZYdOhrth4ZVg25jGo5nFONbWMTxAqO6Q3bna8W3+estvdKcOshASKyRNgiGesTcMnvDVf63yjenBwMmySShMW8UZloU/oc9Z/WHZSIFdpyh3njRsnXS+4TV2FX2NJkiWJO1Y8NqPqRjMo3u+IKalQ1JTIqEWuS6SgUs69ik5i2+aGKFwJfwrXbdjqViEunEDVDPET5XtASis4i/TE/lvWaZTxBOM91or0ZGwTXRoh4r2TcRFUmLIh+TzKuCZlne0S8JaD1Ma+8r3AFpS0r6GvMzYiW9IW3S65muUP5sMyBWI8sAQ55G/p/NPwH6lDxHOYM+hbX5Lt2dUWcG8YTzwDGPHMO+2h39jHn0+7MPxyn+8Ax13ESinO4gXFNHWciSJZIdeaPEcGd3xe0J/V7neQJomSpiDwvyQiOWBKAM0T93Jj4zCEOs71UabEDzx7annmTxQ78ZkKo0XNn5WX5zcWih/skY2XBWPSNWDFb9M3xBgGDgEHAIGAQMAgYBGojYAQL0zsMAgYBg8A8QUDEgWolwXe5Jkh0gGHmbl6QIchYEQiBCcmC2AB5xz5IM0hX/SLO/xD6kG+8aEM0vCgZUkb7zYfQ5TgIUwhhu8rq83mC1tFiCNlAfSGW3ygZskG7AgIbbR1BnUZU3blJZafrVcu1y5RTV1BxWYxfEDc8sYYNavCBHjX0uDCJezpLdacxIK24vvZtDlZa6OGaEHqaQP5z+b5XygNhfY8QF+Bs0mQEdCfXK50hySARtasn+jOEKfghFCHQaddlEItsg1TDioi2RqjQJKQm7xGVSIwHRCZcxDA+IKo7S9fHEoPrQbYShFuGX2RlwTUYD7Qvxzc7lj+0JL7vqQZ36ML2xKF6O+4NCY1Fv+AY+h7jkntAbmNlMVvLilJxx93OVLp4ot/9tWSCUUMSItRQb7AkKHhl+ktbhdmE+Bz6vewu1d27LMJl6aIGvcI8FHJTk6/hDAhOiE3mCtoE0QGRaDx9r+896iMr/lzFxJJht3iMssIm9bjP0Hs5iZVKzlHBVyQuA4LFhLgaJbGCNoSQZgX9KmmNl4pxF2uISem8Z3dHFW8cGVWLhL+/qflutTm4XP3Yplu8nO4q/rJ6u3unWmYdlEHqfVHakTrQplsOhx37Xz/2fftI2Eq/Y7teaV9+CUjZKAaJ5KokdcmiQhPh9KlOyYhNzLUQv3I/omgL9OLTqSEzpDr37FJ9a1aKG6g+CR7ermK26BRiReKGdtKxwya5WL9j2XlXLCtc2/ZzBY8g7jkvCOrFJVRDPGYfFCEj31jn+Le87uwTQZ7TTyDpaWtI25uBu0pT/I1sQwAiUDfCxVMy/zEm52KVuRawECe0IIgQWU2sYGxjDcK4QGh+bEvmbYN3D/8RRaa9ybSJFvqYw/nejAGLjH36NXVmTENW0xf5zrjGQot9nM//2qpg3q6ix5JqBmN6vDnlWeVJu4EhQgTz17cl/4Nknn+ViZgORB/XcZ6wXtTCc5XD5++mklCh3UAhVjCnaqERwaJWor//XDJjQ8e3mYs+P3/BMiUzCBgEDAIGAYOAQcAgcAoQMILFKQDd3NIgYBAwCMwSAcgRiClEBshcvTJU+4KHbIDUxKc37m/YjosjiEFIHkgFiCTOLV9RDjmsLTYg7CBjIGUgbBEvIsuO+SRaCMkAmQspRYasRZSBdAAfVrvDlGrXPwOq7pxlquU1oYp1LFXxdlfZwl1ld+RVan1a2SkvEjGKvYFKn2WpuvPq1fDjMdX/X+JQXvgpbwziSruuObp62m3tV0FukQoyEOFgBTEJbohAEGGQlDdKOSH7IDYggPYQ1Fs+z8hUsqwod/tEW9HfwFeTvayAhhSF9KX96M+4PYPERniAJOc7ZBluu0iQjhz3jimAxeoIcg0CElEBwYPV1IwH2guykuswthgbZAhqab/wAimcK0T3q3JhqmGRfchP26N1juV1lsqEMIjl0ncl75YMyTsiMSuOlczUYxOStDLRrxn3EGsch7VQVTdG4mBoecpWj15s5Z1VS5tT2bxn5fPFICZsd0tjkvNtWb5PfaN6C8EZTENw6vg53HfSqv5ckFLbxjap9elt6lB+hQqcSr0louwlloSXlngSsbyK29q6oiRWUC/aHcKQ+eotkiHJJ1mPSHDzQujaT67fu+/KVm9ExRb5kg+pW7zbVU+hQ5aLNygJtj2O3V9kfz/f6e7uXjJ2+OnmuqGH65KiGNjqQOfIi9QdDFmNr92EMU9qsYtr3CcZa5Cpxq4mt+ljN/z/7L0HuGXXWaa5djrx5ls53lKpJJUlWU4ykqMcHidswNBgwICJxszQAzPNTHcDPYanaRoGZmAaTzPNAGMz0ID9YGygDQLbONvYyLYky1YslSqHe+vGE3ea7z33/OVTpVv5VqlUtZe0au+7zw5r/Svsvb7vD8r0R9zsMIdaXByROJqCso4bbpyYac+f2DO6mA5lY253rDp0RVgEfkkDoecRLYpCvxp4AVG2u1mexUGQ63d/uJy7BbVbouOdkaGKrC58X23nq+0uB2nBPZnjKNT/rHymmBbf0+9HBLlmLOPSrKP5DyC3R/ReoNY590CG9AfeT3QmLCz+t5ON+vQdxh79GcD9699ovxaywqxdbF5hC6HBvSU5b0j6AWvVLIwHEY9ep09aak7IJeOeRQZ9hP7OuOZdyDxv6yYIv4sd52epysX/pH7AxRdbJvo47ywIXMbFzyv/pzOUhvn4XyszH/+WMvMl78nL5Rbs4oWywpV9ooJ+Rt+a7NeXuqDwwDg+G1nxG/3febfzPYW8zml9taoVKG5WSKCQQCGBQgKFBAoJFBK4TiRQEBbXSUMX1SwkUEjg2SuBvuUFlhZUAq1wwCAW2yyUzW0F4Bja14A7BIoFoOUcFuCvVEZbGGIDIG1K2UgQiAmAT84DvDPAg4W8ERwXHLh3taUtkAEACnKCuuHuB9c+gM1oxFJWiBfIAeTQdJUbtrjJ15Rd/XaRD+OjIisy13zEd95I6EZfKpRzve+S6a60nrtu6M5JV9m5XkRE5ta/veRu+OWqaz+WuNnPJwqKK/kmNedVM1fZtuiSmWHXPTrtajdIlby01aXNrpv7RFvhmytu4QuTLpkD9AAkpxyvUEaj/GGVHxcSX78UlymrLdPVvt8ZXD7xGNqOTN8C4AXYMo1m+ijay2z5je8SSCBiQmDBAClF/wQk4zwjK7gvff9c6Qd1AoDj55QB1gBC6TeAsaZxzX3MPz1lALBDkzuU1UB7Ijxe31g6UNpeeXx2JJybk7Y8roX2KjNe0MDHBRTXty+BrKAeRljQV9D6B7y3BICKRQ/ALLKkDrgmOyUFLj9Ycfktu4PuA68vtcbLpaDd6sTxcK3sBYE3tNTsZmHoi4R0fqUcBgK9kXci4Ls1SFqcFhCcZ6RyE8VcgQXR0+IH7O/sVByLE66RDbv98dPxPhEVmdwzPdB2lQPbvX3xty67gKIejBPGzHf2ZchYpq4rplq7877RcuOR0YnGF7T/E+GuvB5IFDf6j7s3h3/r/nP3nadc95B7Tvldnfds/vX5n//eA/Obn3h54zNHN39jv//6F91bvXfd60F4KceLlGnDQfc2uHmx+e8UDfK+6yfkBtHC/ANJDDhv8VYA2okBMZDyp9S6zTCN4yAc+VDFm5hq+tnNXtDx01xYr1d2IaRFHvmZS2RvEaiJRPN4LlIA7kROvZZkcTGrQBaL+uHJKFRUC99byR3YmUR3Mcd5v9DmaNzzLEDqqRVuxPjBdRSZvstY+0D/WlxFMU6MVDkboA6JabGVMJeh//Pe+v6zFJ6y0ScZL18UWZF8aumdRobafMK8QVvJakWvgNxL9U9dBVkruSr7eSZRZ1kmeXuxjms3r0r87EOQYs0FmUWC4KCf9CyzrpXUD7oOoUM9kR+ELsGmcbO1UuIcBtsbld+t/HG1M8QfbsEuljS57OLskxX0V/oEcw/fERDjjNl7lHEjeKaE20eIOcY5RCb9uiArLnurFQ8oJFBIoJBAIYFCAoUErlcJFITF9dryRb0LCRQSeLZKAODHgE0W3uaDGw1BSAe0yO9QNo1QgGDABTKEBiAdxAUgHIt2QAauBdQFaJ/q3wdwl3NY1KPti8+cKwZECFhA+52yUEZALMqNBjPAE3WibBA3AMvmQoh6tNzkW8Zcebzshu6outLkmEuaj7poZL0beX7NlbdUXVBTPcKmvH0L0MqF8XbbrrRN900FOuPvP5UFxo6DbuhbJuQuvuwW7jviyhvHXKbz8s0LUsDd1iNAkkXPpbOe2/D9VRfPP8+N3e25+c+nOn9ExMajiqRLHYglgjUI1i8fU73QRAUsB+zYK3CHsl9LiXaxNAhKsw/QByAN+En/pE3R7DULGcBAXHuhyYyLGQgoYiYgK9oacOlCk8Vpgaigf5iPesB+nmtawVKCz73qX84zpoAw68P5wldeWb53acvYE897tHvr9o2l/U/IugLixFymcQ9zXQOwuxrgFfIADKO+p6df1AG0nqkTQCF5nzKAf1eV+afI5YdH/GzupZV4emOUj3ieXxcO25ldaLk4VvHyPFKtS/VqyUuzzJfVxaK0zVuVUtgddBO1kpDv/lJGmT6i/Ev9fPK0ZlqXe6OWzLHKrup/M4xLpKaMNUW9MbzX/+ny79YVTyLYHuzd8JHkRUsnwuGNmfOxaKAvsIXpYIw/LSlo9v2C8OeiUvqVHUNH54dLnRtDRZ4glcThTvlPudv8h9z3Rh8QafGTp1z/teC26MPdt7w0TOIfv+HIEw+WSu2Pru0en9/a2r+5Eda92Wj8XcKr6RsnLSK0z1wJUB3PfwR8UvPnj/fmWrOooD/Rl3Fh9SplKs3cRH9dKW0RGv7RPCj9ZTK5+/7xYPcaP0tjLwze4bx2LcjrmtcjX+VQMyVtz4sIBC9yKQgVz2JRvezxwPf2qc4LIizaartWkmSDY+0Mj73kw7xvaHcCcTMuIb8hJs6UIJQhGRm/EI2fUIYMWiaSl8cIDUfZuTdjELmSIaruVrZYNj+ifWJWnCn9s36ArOiRkSfSrU6EhZtOdnA9z+MZ3Jf3x4TIH5n/uHE/EuCc+bXM5dsV1Fy0nadg564igR+URcsBERq7VMCqrtY8nevd1yOkiKFBzBvekb33p4JsX/D7sB9nYqX6XJAbp7PI5FJ+oj7Mtbi2M9Idl3eMefr9Solxi/XLnyr/rnKmdxzfDqb8cMUIjNNioJxeVusL1ANCnLmGgQ0pjmLBW88iuM/qN/IfKaMYQeHtLS8AACAASURBVN8qLCsupacV1xYSKCRQSKCQQCGBQgKFBM5DAgVhcR5CKk4pJFBIoJDAVSYBgAUDftiyeAZUwnqCfbS+AdQAhABgITLQyOY3APMegKPMfQALzVWGgTxssdAwNw+ASsIL8/RykxYCHXgvvVoZsAswwSxJKC/gLAQFxwDPcO+zVxlC4HYXDj/mNr1zQpYQdbl4Cl3nkIiG7SVXG55UzArhpmtU16jrogpapFPK1Ev1LAFiCJyMeDaykhyroYvW4GLqCbmRGpH7qO2uvT91fjipOBhSfk46zh8quXRUBEjFc+H8FldqjriwsuRGXnzEzX52t2t8te1icJ+TMUbQWIWgAFADmD6k+tJWH8ePOCc+yxOg0GBGrsgYmbKlzgBFyBkygv5JPwMEBRDEJQnn0qc5B3/pWFQADF9sog0BknkWICrjgT7EeIEMO4W06D/Er+atA+u8I8/ZGu/PO4u18XrSrnSc4p5EXkNXQFhQJkgKSAsIqOQSrSusftSdPoJbKAKGDybAW4IhIxuInXvsR3WoUuDlL5fA37cpSJ7a6rqj5VIosiJfXwr9dbGCRyw0OnEU+UvlctRRXIR2u50cTrN8aaheGkprpa5IDIgQnr8i8SKrC6wsmEeMtDhZtidau3txGgi+vb/9TQsLyArSWDDrRkvTP5aX4hc/JU88mec/qQA5WwS5A1JjzYBbrx4zcHoK8mzfhuTEoW3dY8c3xzPDI17ztUEpY8yfDEw+pGa5MXjcneiseAv3aHVX8NKZz3131y9992xprPWymc8+P8pi/8Mbv+N5Igmw2DqZRFYdHE3m7/vhfe9bfMf+99ncSXsDXPM3ZaZizJ3MpRbT42zk4595efbrWVDuDi/sq9f82kIrGn6gkx/f08lO3C4/V0E1HxOGHjbkO8vJGkaiEaeU5y3ta572Sr6v5+W9aBjYViTlyF8NgmwlkZ9+jOcA0n9MmbkXt08EiDgl+PrARYxprCKY/BhnzAO8jxhr5kbH4kbYPA6RyHX0+b3KkHAkjmHhdzpgzn0h5z+pDIicf631RhEWrzFyftD6SryE2yLbihvVSaMszXdiviL3WuOyVFGHyRVCxGvGaRrq+BrJuxJ4riU5z4nIYN4gzgXvQuYRiP3eM37lj7+UXyhp0XfbNCCqk7sXTH6sdJNVOEY5mAewsECGtDskHNY1Z3K9B9mHRdG3KeMakffrPylDVN2vd9yi3m9Xqq+uJALeSfQf2g/Sm28LxjzKBPQzrFLPlCBh/oMyY565nr5INsWRs1xa/FRIoJBAIYFCAoUECgkUEigkcCkSKAiLS5FecW0hgUIChQSeOQkYaTHoagNQgMU02o2AKizQAR4gKtAktyDEAAm4lwFoY9EO4Mp1pjmIJinvB4AI9s1dzmWtrYAN/NYDkuBq4q+VARb4m/KiyYmLEIAuygRYRplJTZEVj7sbfvU1bun+vSIshl391roLyidc9aaOC0b2uCD6ln6dAMa4L7IxOVE/AHMASIANngdACQG0w1V3AsDkrrzpyy5Ld7n0xGHX2hu5eHZM0QBEYIzVnTcz6soT8y5Z67mhuze5+q6ua+5L3JH3fd01H8U3P0AJ96fdaAeeCQCC1vw61R1NVNxNPOsSlgkqtGXaq0dwKQPsI09kSd8CrOQYv+OGg7agHbEIQisbMJi/ATchKnDTcanJQH8siehD9HuAZ+6Phjb9gDIaoEY5N9fTpc5k/djw8XzNS0biha0b3YH6huRQudZqf7pdjyBbANkhLOZEVKym73b6B2Oa2Bi4sxpMyAtQkOfSp3oJwYNpizYTKps0X1du+SMl92KRiwJ785v8QEYPmQvl52YxSRQHwYvnu85f6MSJDBdyuT1z6cJiRyQGJhgu33d4PjsLEEv5mC8gl3DRdjI93jrlz5PHJ4IZFwttf6C061WV8vyrRtMGQPbBKE+qqedvEGHw351Wz5N/Cp7P72jvefjGzsHy2mT+DSIT3qaA4rQR5TBN/R5ZMuU95UqHOsf/Knvr2l+a/F/dN6LdruUvx9P4xOQ97qsjz3PtoOx2Lz78G18ZfZ776FqZN0XwDaemmxuPTvt5uv32xQdv3tQ+RD82khfXUcgdN0UwIz+jzLxi6SSBctot6XOQZcc8mYjIouWYm5haWwtbQTeO75OxxGg3X1DcikqEb6LI85LIq3UU06JB8HSdjzPAbpKkzFczYRB0Qs9vlmQVs5rxKzT/nC3FmqMgjJmXGc/MicQa+b4zXPSt/eM/1N8C9EN0YKkBIM44x50WfR3SApaL/n3PCvc7naz4jM6BqMBdEeO6Bx5/euknmFcYDga6Q3ZATjLfrtNJE6Hv1cgigoZlATeUZUGVuCC+nHBFeb6B+CAaN/IZpTgWYivEdHTFIs3ojsd1U7NCZJxcbndcZ2uLK/GbEZfIE4sLgnAj6//hLA+HRCRjYUH/4NuCtn4cy0L1L3tfX4ny96bFfn+gregD/I2SA+8eXH1h9XimxLuZOf6jynwHQZANBly/WgimKyHL4hmFBAoJFBIoJFBIoJBAIYFnRAIFYfGMiL14aCGBQgKFBC5cAv1YFqdf2PPW1F9Mm8sNgAHAIdC6HlijDDhkmv2A/oAKADCAOgBh/A1IYQtz9gHguNdl1f4XmIGG47KVxDJoDRiA1j3gAsAH4CCgAy5aeG+hHQl4AnDZcJOvr7nxN9zlRu6uu+EXbJYrKJ0fPOVGttwpQoF6AE4AnOxVRlPSfE9TN0AyADHAOGRlLkQ4HwsPzkFGxKIo634HnL9W1hVjEy45+kXXOQYgfosrbxXwHU240Q2ytqiqPbK2G72nJrJjjVu871F39M+edJ393I+6cE/Ac+pIXQE95yUHLBAI0A1QclWnfrwKc0mDzNinPehzEDPUE3KCPkk7kiwGA78DWHKceBAQarg34hrA/5WR70uTCH2e5wGW05+RP8A/fYH2b/7FwdhIl4VK3gmHkqXxZjYyRVCBLcG+J8Na64TsjEYEHx+VfzRILcbMapIV1BDwFfkQCwDN8W+aKyzX/4eVGdsQPL1EZ1MFvnhDKfv4c6Nkdr2XTIZ+sE7WFZvEY0x6vt8UHhuKMwhldZHrAdVWqzsi30OESZg40l48ok7YQY1/tF7ubFw7THucCVykvxqRec52UgwQt3voyy4tt9yh2rAj0rFA+MkTgayezpJEQCSywHA3dg/Or49nt46nSzvDPB0Erp/mDqmWtQ4osPZX72g9kL35+N+84Mtbnm/9rvekuWjM/d72d7q3Hv6Qu3fd69zRMlPictrcPugOVja7m5YeO/aD+//ojvF4Nnn18Y8vRXnM/IObIuYQXMlQ7p9WJujuyTbo32bQpRSHIIv/UPnzPF65nQxtbO7/vvczyZTr+ZDmuuRLM8nD9W6erutknY2RTEe6WScp5/G87/tHhZi3JfBIE3c794Mk9/IjQeCmgyBkfjKy+myiXM3fmEsPKNt74x/7fYF4E+dKzOu43oHQRJ4k5gaIHOb9lU1jTr0rc/4HlbGs4DpAZe5h4DFbe1dBREJW3KUu19W7U0SPv0HWE+tE+ETqPOUkwT0aw8EplntW1jl1dbmmbhLrmo5eOKOKFLJZb8XNMncRn5FTX/qgvW+Rx6q9G+UuysiWFWV5FuuMc8n+Un5HpsyRyJv5CJm/QxnlgTMliH7OYTwwXrj2Pr3fsBpDZnyHIDf2bc7NzkGYnU8d7F60Ef2M7x6+G8j0UeZq+gsWI6dbr51+fwhZSGPeyYxj3hsWe+lpZVmFsp9P/YpzCgkUEigkUEigkEAhgUIC15UECsLiumruorKFBAoJXIsS6LtpgrgY1PoDEGBxDhAPwMSiG6CRRTegPQASvxsRwCIfwB5SAHAXAAlgwQLgApCdFVC5ENkKvADMINAugAaZsgGGoW1PuQCSAAsoB8AGWvckqw/a+sOKNbHPTf3bu11tl3yOVxS1dlhumXqunbCY4HrKT90oP89giwyoC6AG90OTHzCSxLNRu0arGvAdUJvrATg4n+fOymKj4oItipWxJXXxwl7hL8+Vu/PYdQ52nDcUuKFbhxWoO3RpY9pteNuUG/2WG9yh92Vu9h+eEpfBsykbdeR5U8poDaPjPC3ZYPkCQPJBASGDgYD7RbwqNqbBatYUbJEX5A59D3maizKIGhJyRK6A4fj+xxc+1g70BdqXDCi5mon+DOhPOxKYl/6EuxKAaLIRBPl3bY5yFQhwrjVTnlgj/19HlrrDe9px/cgW/8DnK669VWTFfKXVfaRVk/WO+tEquYE6vb7IB3IH3/C/oYxMBxNj5GRSQywobsVnJ7xkZtyltTxJdraybG25HFYF0kayohjzAy+NgnCp0eyUdX6cpHkkt1CQGgtxku1R4xGQOGlHAfFqwt/+4P1zCtAdr2BpQdsyTtG0t1gaZ2yvu0c/7l459t+EKCtwhtdxsqiQacW5PXzd0Dk8PdU9umEsbUyuS2Yno/ycHmUOe0E+MzEx+0/7prc+OjY7d0wxKt6+v7oVQtKVs44Q6LJbDIfdH2093XBFE4zHVCfTq8UH12Gt8fKZz7xQbqFeuIxn9zTMmU8G0+lkBb8B5hoL8pvaJxYJ4xxyg/m3ueedn7S4DUu+Fy1Ww/X3B+n+euz5r21mebuWB41AzvdSGb3I0oJrm8SsEHCehV7ezDLviPhp+nJzNa0rztiAT/+BhmAM4/qHscq75UvKWCwxfy0L8szJyArOYG6GrDVXWszLg66c7C48A5dEED/M7cgSsvBMpBrjhXboxTpSWqu+vVdExT617TYZ7dSc72eBZucky/0kzSRqLxNBlMoaKVH/j6NSlMrgKJfFy5BIyhNplgxr3OzQCxYihPIiA19uoS4qlsU5ZHS1/UybQ6KyxR0ccz9Wim9RPpNVEb+TGDeQdpAVjEXkB5HINwaWarQh79t2n7BnfNgYsUHP8watZ5iD7JhZWtHvaG/61DetI/uuF3UMF3pm9XM2+UIs/okypJiNW/pftyAlzia24rdCAoUECgkUEigkUEigkMDqS6AgLFZfpsUdCwkUEigk8ExJwFyk2JZFPYt+wG/AReZ8s7ZgYQ5YzgIfwIAMUGDaiaY9ClBgbmpWxQ2CgAlAY+I5vEkZIASgCm1YwA+08skcN3chyBOwGcCDOgF+DLl13/WI2/HuN7nK9jGRA4+JRACoAPACQENrFzAEYAs/1YB/1AmghPsAVqNJ/lxu3n82W+RBPQG92AK8m2yQF5YBkD2AI7i8+JoCeuPuqeGyJHJefcjFT+5z4UaVMxlx6966xglndJUdZVfbueTin7vZ7fvNg272412RGRYEGvCLe5mfd4gjykgA03sFlNBWV0USmAcwRLsYYESf4hhyoT7WfgYgUW6OAWCxpe0fVIYkgqwgk2gLwCwjjlarvhafgOfS9wEbcSkGGNUDHZWNPKK9adcXN/PaxP3uzvqa6Nhjd+Rf6WyrPb5udGG2XO50ljqV6FERFu3LRFZQb+QLcfLflLFiOKMblmXWLU8n/LRdzZLtN0Rpo+IH6wXAVirlsC0riuEs98pCXmMFcA7yOJE/ftcphd5wmvqj7Tiblv9+ntcNQkWLyPKG2AwCPvP8TIBsOkhaKI5FpjgW+LX//5RxqUXfPJNbIHdT7UFXDZouzUMhxytPH8NZyy36PV6hl2RN4WpZZ4NcQLkx7UNW9CI3rJyIpcBcAYhZC6rZx7Y1nnpsqrH3i995+IMPvm/rD/+PraCyTmSFEa8r3uVIeYN72YnPujXdaSfLGjcaz/eV73unn05WnKks9Ku/UmZ+YB/SCRKDuSYp/77a9fcZAi6VNj1zyVPy0HXC99y6SjC8cTGVY6/sRLkchPPNrDZX8quHFKxCbqE8ANNc+8cUDb4tF0YGHp+pHJf7OP2F8Ur9nlQmtgUk6+8rM//+e2XmxPNJFt+Cc1ciKzjOWCUxp0CW8WxzzzP4DCOhzWUYrsuY/zWveCURFb5sEeNMsUEisUXyvsUboaNtRZOA+n4mssiPZXbkp4nOzZzGTV4Xx7a/b92ITgCyZ77g+atq4SICalXer+cj9JXOOQcgn+tdxPsUywP6NPMqW0iAc7nu+1Gd82rlP1OGmMcVE+/7/0sZSzXefRBetC1tbQG7mVtoS97bvI/J9JG9yrQ173vaGLmZNSTjnPJwX9oJK0aItHOVUae4/6hMTCn6GRZuEHI8e1XbmQcVqZBAIYFCAoUECgkUEigkUEjg3BIoCItzy6g4o5BAIYFCAs8mCRjo0fPrPZAhBQC+AAAAAnDvAEAOkMsiHwCNc/jbAFwW7ubC4ZJlIMADtA5XPMSqgETgWRARr1KGUAHEAAgClFAMivq8q+4acuX1mRtVPOHK5o5LFrGqGHa13cOuvO1mkRRcB/AMYAGgAQCNNQRbngcJslcZgAOwiTrxG1qe7IOUsh2U1aCWMMeRmQFkFpeBc8i4iuFduqCA3MeVN7jo1rXS3a3ojp7LllrOG1eMC8GSlR01lz3Sdjt+Yasbf0XD7f/ttmsfNPCLurMPgI/rEeqAm6RbJTdiW+wXoEQ9n5EkoM4sKYzUQi7I1mIp0JcAkCxmChrO1IXjnEeb0ga0N8dxD2OJen1SGS3YM4GWl1JvCCwD2szSxiyIALx66Ve+0bN8obxCDv1sUd2pXlpQSPbmrJ+mi16WzQt1//rhTWsWLiNZYcWxGCeAv8jkp1YSAAWuePmHb42Sr06F6Zp64NYFftBM0yxQXquozXUhsZ6AWPVHeStzXiTn/NIal3+oIEhLisySB15UKUebpU3ebXWToyI5UhEXEHs2h/Q0nUVUWBE4zh+0JX2TvkHb36N88rvyZWN/72r+EjixBgqhMlbGY42seGHzMTeZahiJUVmbzB0TkdGQG6gdZyErAMwZl2hE2zhdCG5xjS827mx8YfwuET75BgXaPmOMDKtQNW25X3743T1LDLIcM11of8PqAXdFn1DuuXZThhxLe0TFyilrp9OSbRJ2s+mwnW2dWchrFQXgfnwyCmbFnO0Z9r2SwHKsEDRGFBval4+tZQKkJNKDftGLLySw+5wmKBdaoXOcb/MldaOeH1VmDmZOfLsyhPQvX+IzAcQhN/9AGUs4xir90oIer3R7I1Mgmemjj+EOSuTDZC4jChWv4ft5rC42rFbBDZSE6iri6AK5geLvRRF8y8Pfk8sozxvTRVt0/LjiXmCu0dVcCKDek/uFBt2+RHk805fT5sgeMo52oJ9jiUBsF4jDs6Up/fhvTjvhe/X3x5UZN7iFfIEyZD39G0IE8gCFAsYWSgrMzRAQzDmQplwDmUibY7lDWfiu4BzS6e70zlQ+LKj+i/IfK9u7fjBmxZmuK44XEigkUEigkEAhgUIChQQKCVxGCRSExWUUbnHrQgKFBAoJPIMSGATgDawHsAf0gaAA6GPRb26e+Nu05c01B8dMmzXtu566qCoJdAfAxg0QQDzAgwGMaJDzvIYrbdrsyusOurVvnXbJ/BpXWjvkfLkbr+2ecL5c8GTRN9zETRtceQMAmcXkABhEe5Jyoq1rrqSoI4AXhITFwOB3tPghNqg35wC2AvwNAnCnExbIjXMgKzivZ/3Ql6EB7Kb9CeARuSDkvgJUx9a7uL0o/d3IJXOZCJhRuYRK3NDz227nr4UKEn7EHfp/ZXkxA9CCJQzXIRPuQxmnlN+h/EXJ8NMiLajTFUt9ooLnUS6LVQEYyL4FtYVwoKxolqPZCogEKQE5AKjFlnIDaEJwAGaaBjYAGHJ9vjJardwTIGq10vt1oweUAcEA2ehr1v5mRdQDlP/dc6pYDwBUoek7K6uAjW1Xma/W5/c/0bqpeUvt/vnqic6syIorpXHL+GO8QlpsV8b6BDdD9L+7lPdI6H8xEuTHR0p+NhXIJVmapiIn2vJvI7xbMbXTdKHZjstR6A9Lc3wizbOqSIy420rULrmMKvyS6AnFr8hndHwkSTLackzg7Xq50Yn1dyIri5WA2Z5VhjJzyO/2ZfY/adsjByajo7+3Ljq8S8YbUZCnCk6fm4uYp7XrSNp0O7pH3HPaDGUGTyrSoLtOZEVzBbICkmSvMn0Gd1+Ul36HnAA2CV6vMfpreeWD/+YpEQ9/IFX5g3L59PP6zVyTnSzDy058pivXUcdvW3hojYiK8ob2ETckq45SflbCgmfybIBOthDBjAkCSkME25yZiaw4k9Z8b75pZUeDTnakHefN6UU57ZpPJkbTqBGtL4892cj8xZHIn1IbGwHL2AK4ZSzhbg2SiLI8JPICEJ2xxt+Mt6c99zLGQOBZEN5YW9A3mcf+Rpk+wrzGeAOAPp9xzfjjHr+gzHxAok6MX5tLzmaJYBaBbG9QP8Z115KseyYUQ3uX+uFEFufDiZepTJ7mMAXXFpvcfwtiakSIc8WwkP8wl8/Kxs0pfoU8qslnlFOg7mVChnoxd1w2iwi1J/VmTiX1nnMZ26//mPPeUB76ODEekMdnlbFkgXAmtsXUed9p2fKCbAk3kZa4v8WaMItLyG9cCa6UUHy4kIS1B4lxBWlC/+L9gPAva/teSCGLcwsJFBIoJFBIoJBAIYFCAterBArC4npt+aLehQQKCVxzEjhTUG5VFFcWFhyYhbhp4wIC4PYAIB+AnL8BvkiApWSuW8n9xnnLT0A74NrPKJt/dwv0DeC234Vjt7jJN4254Tu6rnN0Sn+LrFg/IysEPXkmcNH2I668aaPUW28WtsS9BuMmcA/eZWY5AiGxbPGwTIwAUgNyUC+sGEAiORfABeAFbVHuae6muLclA4y4JyCckRKmeW7EBkCHAWWmmW6AR+aiSkuEhfymb+oIAOu4YKjihu9UzI1gwtVljVG9Ydod/C/3u8X7KQP1ATAH+MFagbLTBlhbvECy/C0BsoBDVzINfisgC0gH+oS58DJLFQukTXlxD8U5TyhzHLAd1x9Y2CB7ZEZbfFoZ8B2LF/K5EuASWrhnSxBaPJOA3rgYgbCgrQG0AbZ5Dm1oroS4l4GPAKbIvZSpSWeS9Yc/1Hj7E8PhfPyTE3s6sxPD+W/f/9ZTni0C41xlPq/f5W5p0IrBymQa7D+nA1jz0A8B+JDvx0pe/jeB50YWMlfqJHE7jBRa21fw4CSrtTvdRCr5wzpSirOsEkhlXDxamGaC7zWqPLFqIilKsqzY3u2mLXX2Q9LgX8jS/IDGWltWFswLPdc3kBa/cipAi7wYY2hBQ9rRlv+H8iMiGVBRRx/968PB3HG5MRoVdfI6XcAYUQxz/80l4cQjacPt6hzysKoQQdGzwMD9kwJOO5EV/D3oxokxgaY94ChjBOKCY6ZR39N4XyYrlpPkmbgPzu3V7h8qf0n3+1WRF9xzpyRArIp2I6jf94Zj9z70mYmX7Sln7dabjv7tdCnu/gudN9jI3OO9yswHEHFYdNAP6cs8D6aFPs1cihxw/3RWMBv3PwKlk/3tj2hqzirySrSvm1WaJxQvPXCHvFYa7Z2O142tL7lJtS9jDlnTn5m7mMcgbCABIAlwzYUmOnPGPykjZ8rCGLM5HTdU6aXEvTiXyyDqrfkJOTDXUl4jMJgf6Es/oszYpU+hBW+utoiHgbUM12FpRf0Yq8iQephlhc27OrScBsv0K+jHf9MqiLovx7BgrOT5BrmCWpunIiokcb0rY/V18XiKWuFlLblHU7/MEgWEz7zQzxWcW7FeFAHdyw4kSRrgJkr3mVCBzK0cfZ56XJYEOdEnLZDBKcTFZXngxd3UviVoK1zEMREyvoixg7UEc9alpMHA2N/0GXcpd1y+FpL1V5UhgZEvlhmMZ/vOuWxE1KUXvbhDIYHzk8ALX/YDzBvMvWzJpmhh37iDSjr5fZ/546Lfn59oi7MKCRQSKCRQSOAKSqAgLK6gsItHFRIoJFBI4JmSgFlHgI6pDGjgsmgBcABgAgzoAX79Y4BLBnbZouaCi94PrP0SXQjwAJAHeAbgRgb4abuNPyhHHNtHFLxaVgjt0I3eNe1qN0bOr6k84awbeRnAJC5RAK7QkKbMXA8YBcBg2sRYUeA2BE1nW5AB7rJQA9wzcMnceZiWPUC6ac1ynYFiZnlCvZGBWWmgSWzkhgFJgDTsUy6SuZPgmRyriWhRoG5/Rk8CsJMFieqfN5fk5kquor57RO6i7nBP/doDbvZTaL4DngBGAtyhvW1thgx/VHJF8/Rzlzsgd9+6ogcy9+qwLEfkTqaP0B6ApAZaQxIArqIZzW8QEZQdEgcAE5CP62gnjt2jfK5AqLiEIR6JpbORFWif71UG2AXQh3igLZAnz6bt0U6nz9AXT2qiMz76Lo/o99yDfnRIMXkPTccbYvIVcAM1UM2Tu/Q9+hHgL2OAOjAm/o6/1wbZoZdGrcN3lPKhcuydkPuncRlOdMqlIFlqxpATFV9ubDqdblMgfcVLPUVK8Lw09+T+KQ7VaSNZWchv//L4UJtvkOuboyIylkRY2DciclrJqsRIH2RG/we4/4CIiqHFZKwpK4t2ye/Ude+yjv2TSInmzR04Bvfh9cnsmDTZd26Lj/+4yAmBynlA0IBlZCWnjQCpIRPNlzxjDmAbcJ7yWDB6m5/y6sKcCJ+nidACBn9VZfgxyaAu8uTOWtps1NNGWsnaw5vah46+Y//7ZF6y4DZ0jpRkEfJh3QUXR8gZedOXITXpux9SZvwxt9DvScjBsjsXWWElhDx4zwNv1zyXL8joJepkc14jOVSajf2FZtZa2LYM0WJtRR1xaQYkT782KzHmA8qE/3+OM0axYqDfQ+oYAIV1Qk8rXiD4U3ruBfu7sjKfa9snjHhWR/OUaatbMOQP9MvFO4dYH7wDaGdIFhKWcpT9c8rMF5xHO/fI3/MIesxzzfKN+zCvb1Z/vlk/QK7OBCK8dbOOSKB55XImDk9XiKPLCTYvPjkvefIJ5Qd+GoZO1kd+i5guGgvT6qQzOgWymDn5lNgu55LL+fzeWJ2VagAAIABJREFUJygGT7X2GyQtzudWF3WOSMnB6+zdZsckf/jSFRPtM632Zkwgc+Z32pex8p+VLU7URZVrlS5i3mDOpF8xlnlHYGHBu43yJupfV8pybpWqVNymkMCyBERO0I95FxgxwZb3BEo7vJ/NhSnzLfOuuYDFOpH37aLu0SPblVckLkRoFOIuJFBIoJBAIYFCAldcAgVhccVFXjywkEAhgUICz5wE+sRFsqxkKshw2fLCQD+LM2DkxUmN1gt1ByXwAvDsNcqvU2Yf+I3FEiAUQN8ut/FHd7mR21/gok1VV97syy3SnEtPtFww/DVXkmuocAQwG1cygFYW24L3Fgszysw+Cy5z7WOkAoCSaSUDlrE4Y8EG4MsCzvxUs+U+gOeA8dTXLCVopNM1W/ndXDXZ7wYoUxYDlswqAnTWfse6AEB/2cIjjOS+p9Z1WVUyb0du5M5xd/Pvvdjt+4/T7thf7pZLLM7r+WBXNqAfcgCgHQuBIcn4YwJZqNvlTMiatqNOU8r8DRiKfKkbf9O+yBAtabSmaQfAa0BUtFgHLVuQIa5DALfOJ52MMTFwMjLAcoO+gXYsf/M8QErKQpsD8AJ4I0f6D1uzMuK4aQefvjinfLQbWsP0Gbv2fMp6yedgZbFC6pVVhIqB9NSd+uY/tLAnWTtRL5U7QlejICyVZE4RRVsUSFuK4fm+ZrO7oNAVbQGwE+UwnJSmuJekaSj3NotpmkeywJCSud/sxKniXqRdHWuKrIgEzJoV00kQ7wxlo7gnNTVVRmTrxXL/f2P16xzH2kUDy/Na8rKzs3PIV2yKwwrvHc6EI9XEBX8iX2lrRVpw7puUcal0vzLPp/8bsYQMaF+zYHoauHiW8lGErsoGcB/JwqPRDGrtKIvbj9dvTD625jXpu/b+36XxeNZcynH+IIkLoEP/gbwwkrfXb4yc6Px4b/+CU5I3FwKv8mWVSc9euHNT+UtrjnXXl/7hxO07tlbyhVeMedMC1nk21hzIwsD9f9S+EQH0eQhY5iYIPc4jMachL3MhxbzBuOu1yeVOBgBrnmKOAjSjPZExiXmNOd3iB7EPYs4YRcYXDB4TT0KgO+1C3+G9UFM/3iuiYevyy048ncs78vk0JoMJWVR47SDPK7KdyPxcceGdn8pGpyWrijzu5PKtJkulLN8moguLo6b2j/RJC+qz6tYV53D5dCW0n+19d/qW9jLZ9vZX6jsiNOxdt6Q2pw14z2N1hUUYfRR3dsS6uBJrT94bkM6kP1WGoGC8UK69yvyOpUXPyq4gK1Zq0eLYlZaASAO+9ciZCALmzJOpbzHB3zY+Oc+ICCOs6d82h0JM8F7gW4i+z7hjXuUjg7gzKIKgGAM5D3lnLh7tm4fn9+ZhrC94fmGFcaV7RPG8QgKFBAoJFBK4Eh+NhZQLCRQSKCRQSOAqk4AREH3SAvCFRZBp3p7U7LxQooJq9sEKiArcp7BgQqMRLXcWP7e60oY1buTFJQXTDtzYK4ZcPCul59aSiyYed2vePCprhBt03kuVTWMMkgOwn8UZ+2xZgHE/gGWzuKDc1IGFHKQFv3EvzgPAAsAw8A4AngUZ57IPSGYxGqgGyQgIs0YZJDDsN47ZQpBy8XyeDahM/fkNGXB/zgX0pCzCaqMTqknN5QrUnbRbrrP/mKs/r+I2lCru4HuFKXchVwAgAfqwHqDu/I2WL2B9IFn/1WUGW5APBIX5x0cL2ha/gD0sjgl4yiL3PmVc9mBZwflf7dcZcgO5UG7qgtUNcjiXeycIplcon54Aky0mAucAjCErykNbAmxjmcFCfZuyAef8DthobdG77wp9nP7CedauKxThyh8SID+ocd0bq7+o/Lt/81AaRX47COV4P4oORyVZ8ujMUhjc3/K9W2rlYHOShWX5aep24riapVkiH/1xtRS05KJ/SArk8o6DqyavmeWKOC3kXMDsMYG9PfEoD7pJO2vF+2XsXfmzp55pxzL12YUv1Hd7uzoHF0t5vCSywmLLQFTQL2gnMvIfBGCMGFmxDKdpqD9NQ7zvDqkj4gJCyp+PRjOVN/0l/aHcFukwaFVl9eaZPXINcoJzzteC4myCGnArFqZ5W67y2qXIq05kebXqe3FVqPmO+xfzfU+23EM31dyU2geygbHHmKFM5gqLOWEwYYWCPJEdwJSRu4w7yKRecIQrmfpWF6nanXFnpCHjy+ZQinM+FhTnU2zuuRwTaTkfUT9Wn/ZeIddoWNPdr3GwU3Ep6rLoKceZWyv3T73zRWakYvIj/e7kMk3Jaysid9PPklmRenOJy5i/VO4c6wpzq3g+ZbrqzxHRY25jzIWMzTV+pQynSTCaIJtfavfqfR7Bxrke+X9EmfcC5BnvY96LEBi8x/5cmfH9ZmX6M8d5V5wrUQbIx6kznPgeHf9PyrynflLZ3gdsKQPv556V1qALuXM9tPi9kMDlkkCfjOD71Kx9Mx1jLECsGXnLdy7fwfRd5ncIB76t2YfQ5jueeZ6xh/IIY473xiuV36oPnUSDXEZkOUoljA1Lr9IOtokcx7UbcZm4D8/hXdlQWTjX19asKW3+O0leFhYYAxItdgsJFBIoJFBIYNUkUBAWqybK4kaFBAoJFBJ4dkqgD9hibXEKyHcxZEVfAt+rLYAyGl6ARCyOAC8qzotqbu1bWiItGm707u0u7Rxxpc3bFGD7hIsmAfJZIAEgAbaxOAJwAzAEOEeLjEUbGsK2UOMZnA/wwQINQI5FncUnYLHHPQArKIsFjDbwjDo/qQyxYQDaIDBsICYghwVdpZqDlhhmmWGWHoP+5bm3+W0HPAf0ooxTyixI94ugiVxUG3Gjr9zhqpvmXXz3JufVcnfgPQ8qJizPJPYH72tkaDE6WJzyG5qr/5UCrWYaCLZtdUPO5pfetPrQUKWNKBPlYQsghBwgJUi0HZrTtB/xKmyhi1sd0k/36wCAyUKZ9qe90PybGqgTdQfQxlIFsB5XQWiPc09z7cE96B9cz4Kba5A/dTDXWtzSgG/MjE4uuFfQ0F91LeqB+qza7l13bE0f2zvTrlbC2XI5VETt5IAsJsZEPgyHkbfQjfNNsUwnhMbKnEIdVyGEBc6WtOkmivasoNuYWsl9VBbS7tIkRygQP4wh+jl9rxd8uy+7k2UXcHne9RBgbSm/q/ENIxcNwLaYBRw312ynyP9cLoG+AoS5nAx8HZzPiBmREzsCkkLnPA1wPo2IoBznOufkAy/GuqJ/sWm8bhfnNHe4u2VB7rR21/2l6kKaHIvzgDEOGAUxAXk3OIZOkX1fQ5/7mWbu6WTGebfV5TjxtPYbnGNX7XF9Kwv6DXU3om1BI16xbOT+yXkzGvQn5H9Mc6y3VcdFGDuFeJFfKDEbCljfEXXS9XI/1cX7FI17T+4HB+RJ8SHNIkc1VphzrM+uWrmvghsxVsySLwlDvyw3WEOy1FoMgyCQi7lIf2dDtRJzQldzQXw20qJPBBDThHHN+5p3BnMzswCkGn0aKzF+4x3Bb8SGoe0g1ujr9yjzviYGEUQH71XIcOZ+s6LBeu+Tyrxjvk8Z4hpXVNyb99EfKTP38/43gr0HABdkBVIo0lUiAb7xjIjmfct4oY+jLEK/5W9cE0I+MB7o93yzmkUr39h8n/F9qWnLu1XfNq/W9nbP06XEhAoiRa2SPWO3rUg9vVf5w9ryncX3Et/spFuV/1YZsoJnQjbyDcWcx99mKbdX+4xtvsUu2Bqu/6xiU0igkEAhgUIChQTOKYGCsDiniIoTCgkUEigkcH1I4BIIipMCEkDxev2B5hfkA4CBgSAE4bxPrp6arrxhvQvXV1x154jrHj/kqrvmnN8D5lg4EeyWrS2GuA+LOfPJDigNmEoygsG00gAYAfAN3GdxBWjNIg6ywLTVDHjlPEB3fuMe5u7FLCK4FoCKMphbE/Y5l3pZGdgascHzKRd1YPGHhhvgPGCLWXRAxrAIZYFpgcjlCisccqVdmQtmNrtNP1FxpTUVt/jVeXfiY4sumeV8fNVzX8ppVgu3I3OBL/f2y7OaG3NzxeKVBbHFO+m5LOjXGYsVLCkstgREFW597lFGVtTVYkcgQzTEcWuDZcTLlJGXae3t0z5gFfWcOq0itMN7+78jC9qURTTWFshkrzLglsURAfjieZxr5e21+2r089PK9oz+CQj//s88mbRayZKCZ5fiNDsmIKKtGNxjedKJkzyUZmXJL0lKvhe05OymItf9C4kAceelVcW5ILJNM8nYyZejXyv+tSoFYAIgYQTAJdXzDITDSsD1xQIgg1riRiiapUTPIkWkRW+cIrNLqszqXcxYpi/vDL3kQDur1hX3o6XtUOhaR/5upvToDVWZAwS9ccO856vsJ4kU1cdA+bNan6xeca/+Ow2QFj33KurTkcg45q9F8ZOxeIl9iqrdLoV+PRUjLF9QowreQnRueU6ToZHGgOi91Mu8EzJFOiySYkFDY06cn7knu9j+edUJr29ZQblsnIicCMuyulonq4oRzZXznW4iK6y0VC1Hi0mSzeAea2yk0ta1PbDyPIiLHkHYj2liwemJD0NClry7aB/eu/RnyAVA0r9XRubM/RAbfAOIeOq9L7iO41PK3IsxhJY45ATXMh4sUD3npuciPPvlKTaFBK6oBGS1YG7xGCf0W74VIfTM1SbfeowNgtm/VOOPb6obmLCkaXA7BmFSQsDdnd4U3h0KwHODL7MxhnSgl35U1mtD5wZRpGA9qWvNTWvLp5MnBkMPzJIegbFsUZkzDvkGtwRB+Clls9RjTkWp5L398vFNbTHbrpZ36hVtv+JhhQQKCRQSKCRweSVQEBaXV77F3QsJFBIoJHBdSEBgBMDxzyuzoEHrC5N0SAesIizQdd3d9JsbXO2WQCukOVlZdFztJgBmFmws0gCrARtYuAE+A9CZhQKABH/zHEByi6Fg2tKmlYa8AasBy1nkAX5QJlwVcU+AcrTTAEK4F0A7Cy2LV2DgNvcF8AYoMc1M7gmww/3RCkXjjWRgYc+RyMAxA31xmUQ50IzjXpQfSwGsRNALZ8sKUm6iwm+4YP3tzh864dZ9j2pwp+/GX73GHf2vm93cZyxQIo8ApEF2xLXwJH/A/18VKGP+6weKckm75g6LLc+jrMgNUoI2m1IGQMICw7T9WNDSVsiLLTIGSKINKR+gEySRWWGwSEaeWMBsV6ZtAZkgQiy+CPJDa/bz/edwHs9F9hAqBlazgDaNXnMnxL2uSbJC9bKUKThwK0m9pVKYPtBNWt00Tl4e+Z0dgWtNpMFQIpcu8u3izXa7QmPzdFGxKg52Oimyl2ecXKCDByh+QgAvcqWPI3u2vf59Hm5gBopzeXZXCExsD6KtTUscoMfc3Nm8YPE/erFMdJ9ef7gKiAsr95Z6sHh8JJg7Ug0a4eHyts7XGi+o/vXxfKLiu8fetcV7SeT1XK89pLJ/jnJrSz2/Qxlg9gv6mzF0Cmh0jrgIl6eRroK74rKpD8b3rKwg4tQ5qgLueiCgCAiB8IL4ZF2BuyOZHbV1TiBgXjEuFLxe/vi6qVsSIDgnw4IDEipzCmB7cjWMg1UWsZHtJcliTRQGfhjIaZznz+if8U43HhciOq7RFcsqqyI5JbLCOlGKwulunLSwvDpPmQySkzZnc4x3H3MN3wtGwJmygVk6MW75PviHfh+nXUnEpuBdze+8d6jLRcdBWWW5FrcrJHA+EuAdTP/lewkXlXxfvViWtxu1/3lpE9ypWZ3f9H7Ox70gfGFYqjymbSuNu7dpnD4vLFdkvSzG1Q8W/SBkPIRJt+NK9WEXVZb1ezTn6Snd3rEw0ulBsFPXuzTuiMBIXCrLC/7undf3B6nLIE7eqIz16yeU+e7iWw+XrcyHlJvYNAdFvPD+MdLlafUuXEadT1cozikkUEigkEAhgdMlUBAWRZ8oJFBIoJBAIYFLkoDAcjS+/qUygDPAAyADwDYLGoBqSItDbuoXtrh4qaqYFZ4bedmnpfIFAM7i7HnKABWYp/NeAqz4Z2VWWrh4QIMLMgAtLwBvFm8AFlwPKWB+t80FjLmUoV4AkxAEgOUsDAEy9yoDfr9WGbCPMnMfc71kGsyUjWfzO9r/EB0syiAbID+4J6QIAIlZfRjgYkAkADogGSA8gQ4BVXBpwb25B2A+ZbTg2RAQgQvrTeffUHKtJyacF3pu7VsnXLKw4JYeQJYAO8jcSBvkwPGfU1v8jkgLynxJSQtlfB0bSYG8sRRB/mbhQjkB8ThmpA4EDsQCZBXH0YhFbpAptBd1ZcFL2bE+oX8gO8qLP3Nz88UCmPoAav2NMnLfqwx5RRua8x/anf5gIBXtRDIfz/0/pV074PrJDl5L2+952Y7sD+59uOfDOvQzhbeeOxT43Scir7tOroaOttJGUvayTbnCCzfSqgDbcpp71VR+/WeTJI8Uy2JB7T2jjOwYs0bSWcyPq1l7ctAFFPtVacXL0CRvKRD5sFzZCF/NU/0QzCaucrSTtyfCPNlYCzsC+dNnmLRgvmPeGVIgnzvXlQ799f1L33Iw9GKNE29LnLvwsWYvnohi+/TmyZ9SxmKLccO1jBOs2ghY/hv9cXKyrSB4rlfSQrKweZU+MSuhPCIgbpvmgnWSpwgKzU2eNySQ/pBIigPtThKJqKhIXxnZym9K/pRk/qisCpjnGRO4QbpmrCsG5r8eYS/3TzUFqxgqlYJ4fHiIcV+bW2zemKb+rVHodzQ3DAsc3Sl3UYf19+FapdSWVZbcaeWQQ8T1OOscsYKFwynn691l5ARFQ85m3cXfdi5tYfu065kI+qt5vrqWXj1FXS5SAgL4+b7i2xDljY7mops830mpINB+8IYgLG2TtcQakQivl+lX1Q+iPxeZEPlhdHOpMtTIku7dUbl6o/4W9xBputKQ8bxh/Y0lpSsPaXj4wbImh170EBGhLC58f6T3d1CqSm9INmbKEBbtxVnnR7FLOi2i+fStLnq6CrhYRbmEb1/KyjcvLtv4TuObg7kRl2xYSj3WmztPI84vUkTFZYUECgkUEigkUEigt9gpUiGBQgKFBAoJFBK4KAn0yQp8R9viC5DBrCbQzgLYfsj5tW1u6Laqq9+63w3dDhjyfGU0uiE5WLQBaLPwYWv+cyEOWG+xBeDnPAPNTXveTNUpv1k68Jv5AAb4ANQAEH9OvzwQGK/qPw9CxIJIcy6AO4A6oNVeZUgBi38BuQGpQjl5f5pbJBZwLNLMHRHlMK1VtNE4l3JSJhZ/kBuA9ZQLWZhLAJ7FvZfdY/jBMTf5hq6LZza4xje2uoUvtV3WOeCaj1AG6kh5eCYZ2XDs+9Qmf7oapIXuRVtSRggSiw/Cs2gPZETZ8UeOrDiHyIz8hr9xFrbUEWIIX8uAsgCrWLiQIRewlmCfcyErkA3tgWXFXmWIklcqI0/6Cr9xHvvIiWfRX6wPUB4jjChTrz9c62SF6thLP/b6W1KRFtKerM9XsyeOCbN/WLY35Zo3vavk5kf8PO4sxEN+nqybHQ/3j7TziTjNy92y3wnFWSxlmZd1XbWZ5lHPfZISMmTfrCzsUVfjlvFGP5DXiyyT9vxQq91VDOWS143TYLoVJ/N+aXhPy23Y3/GOTVVda3en29hYytsC9Xv1ewaJC0BYCNrnBl4y+XjrOcc3l59arPqNtlxDbVAlFpPcG1HlmDe+UxlLNohAxhdj4If6DYK1BUAS1k8ngfXrlbSAXBCQznxA+9KPIX6Yi5HZIWJWyIJiU5K5SJYEB/GDpkPVPM3GtCvrAndAGKAR1syDAPMr9v0LieVytQyevgWKkdIQXxDoGxrN7vPlIma2Uon0XvO2icS4WRNpR6xfLN53jQgL9S2c4ru1JZlidJO0sXHtMPPw02K+XEhdzzPGySARUZASFyLg4txnXAJ9koIxxzce31A3yzDiprDszWn7Os0/d/pBPhJWo60u80UauPVBVBsSWeHSJP5BXy80katOZMVtsqQQrxGKhCiLaChpOOIFSv9q4up9+mi/R2JoWhPx4YncWK6/bdkPlo2CIS16H6wqAPtxp+M6jdme1QXxffoWF9+qUywWGA/Zq8w3KIopzB+8n/g+ZK69pLngGW+oogCFBAoJFBIoJHDVSKAgLK6apigKUkigkEAhgWelBHBTAnCAFj0LFcB7FmKsjlgNPSWyouM2vKPrxl69yZXXmU9qzmGRg8a9+ajmfABsACYWPADZ3Bvgmr85j4UeGYCexHFzxWQABsfMwoFnoPX1I8q887BwgETASgJAFpLAXExxH3sWAZ6pyyP9++OCid8oH8Ao5aa+APVYDrBQY81nQKERFgD95vvcCBUsEdBWI1g098G8nntTZiwyKB/34drPKBh505U2DrutP73OHXl/3eXxEdfag/won5EkXEsb/IUybULgxNVItAVkDHWAMKANzGqE+gOcUi/IKeqEvCmLBd/mb4v7QZtBcFBv6mztxe88ByKCjOYepJUFSKddLIaIfbcYaUQZOJc2NzdAJufrDtCCtPjaJ35W1gXuhHQn40423Kz5x9uz8bo1Ve9EKU42ho0sP7zGPbi2HDRHjkY3PJykbqadDR8bj/Z50sEsSxfTj7xmpGAq8UwyFe/rvuCc2tOr0dEu8h5mXRHESVbqdhNpqPo1ufZZL6JiXTdtl7I0C+JOulmDvVbP/YmaHyrAuDs8HefDI4E7ni22l0aHK2k/vsUZNegvk6UC/RbQB2LvOUPBws13jfzj+PF4wxMikXoB6B9puqWvLuV/95JRD9/izKuvU1n/sD9+PjUgN8hf5jqIww8oG/F0kaK9Ji5jDjCXQ+wPC5SrC8uT5Q3zRs8V2rCAwE2ajXAb1RBmd1DbJ/X3QVkPQFg0REhcq7I0Yr8ugHNUru9DAaLbukl2a9aM5fXJbyljbhfpeKb425DKt4oFnhBRMZKn+ZejKNi/sNTpXIBrqGuiYxWVKCRwugRESKwkFLP85buR702+6/gGLGkeeo6+Gr81LHm3V0e9TS191XgKP7F2ey4LiCxpzgW1xWlNW5qUZHFR8koV6bEsh08Lqxqy2kJQ+P5yuDERE73fNMehqMFv9n48a2NxXVRjapQ7yCxVFJtaIFbEpSJCuq2GXEX19D8I5t2L99N/97xG2yeVmSP5JuebjgLw7cz3It9jRSokUEigkEAhgUIClySBgrC4JPEVFxcSKCRQSOD6lYA0+TETR2se9z6sogDMAK3RtBp3td2pG737C652w61u4luPunCCdw4LGSwdSCzcAOAgAQDuWBUB/kMOYEUAYA2YbRYLAPTsmxY9izFzB8X97Dz7nWOA2SwOOcbzWTCSKC9lAYy3QNmAUpyHtij3fa8yWswQGlgIQASYNQVltbgaPIPruCfHjUQwAsN86huRgny4D66U0KxGDlbfG7XP4g9giLI9V3nOlbdlWizuceu+a8pFI19wR//0Ntd8gvpQZkBWtNwgCb5L+SG1zbw0Vj+n/YtOfbdQPV///edQR9rLZEj9IFcgJZAxmt1fV8bCAkKIOuAeivpwDtcR5BxwFjKKe/E37c0x5MM1kCIsgiGLkB3XIgvOpTwshGkjymNEBQv0a9Fdi6p4fkltvuw2LfntIPWHwwV/qnOsu3muki3ODfvBuCCPmXI4HQ57h1zdm1msegvNoWi/W/JHg4q3uGMiPKCxlity5/zHy34j9+RJq+w1s4q/UP6Fj55CChmheAohdLrLF5XHUg+w0e+Xi0CiH5RUdNz7yK1PVpdxRXl+qRNVSoJTQzeRxun4SCXshC4LTqTphtk0mBMA2w5b2YO3DvuHdX6zouAfug/j90r2I561XH71e+nUDpX9dnk+mZjE6kXHHmymrvThY+7Ru0fdIxLk7Tr2BuU/EYHSEnFBPBjmiE8r93ygK/2xMnPDn/THCsHGr3nXUGewfqDPWTwWcx/UEuYmF3c58/BR4Xp75BKNdxdJc3J+RH8fVm81l3XXsrYwY1MxK3zFF/c0l3vDsqCYVZCbDQIvS+CdYitq+ncEJpDYvfptUfLLIvmbky+aUR1rVCtRp6GwOdbfbOAX20IC17kEmNuZl/kmtO9djvG9NxVE/i/W9GYe35QrtkRwXN6gJqJy1ioP5UmnWR1LOl7PRVMYyZJCYSpCuXHC5ROkAVssKGT51NuKnGCe6+E6spJYlPUFz7uQxDeUfEWFsQro+eWyr/g9PYJE1h19e9Wem1BLKNswb/KNR8YC4y3KH1bGepZvwQXFrrhc7/0LqVtxbiGBQgKFBAoJPEslUBAWz9KGK4pdSKCQQCGBZ1ICAiO/Xc/HrdIOZUgKFijEhOi6cOxhV71hlytvbLmR54VyA3VQgbYntBACnCOOg8UtAOAns7ACtOadxAKIc0gcR5MecN+C53IPA+rNPRFAFGC4WTWwQEIj3ywQWDACrKO9z/OmlAnCDeFi7pgA2wHHOceIhpdrHy3nu5QtXgOWC3cqA2ZZ/AkWiraQo2w829xi2b14DoAOvxvgS/1w8WKxGwy8NPc2nLccIyKINrtowzGXtfaLtNjpqlorPvmrB13rSRaKWD6gpQ1EDKlCm3yP2mitQGIWj5eSKAP1gVCgLMiIDNiHLM2aAZKCRGBUfqO+ZMgKiIe9/eOQP8gNwsECq9P2WFXQ9siH/sFvyJT2wCUXxy0ItBEVBi5bGfpFuDY3AwSAVdC0J5EN5I/1r0qQLUbD+aN5yw+azXT0SwIV9wWuc1c5PzG6mI09Wg+PLZbdUrPqy/ogCwPBH404L7mR4Nj6mjc7XvEXm75LbxUHBIEGIWcakxBJ9AlIRkikk0nlS9XfToL9EBg6Rtl6Piq0z29GgEFgXHA63cphIAi3wFSv3OkmI0utWFZIbqTZjtfJyqIsrzWVTjetxbk/Np84f6mrbVRpiG1ciIMkW+t78WQ13K8bRIp5QUyLK0lYIBvkyBhpqw2iLy++ZOhAZ8cOQUWMM36b/MpivtjNvN+X+cvmuLyWAAAgAElEQVSP9eXJmH+SskoGX9M+LvYgL/p+P3pkK/Pf7/b7xQXL+hq6gPnBiE7mEPZPWuGhVqy/OW7uorAgQ+49d2gE8L6GZLFSVRRi22uRA99tKEdhOQ2yNYoBMxHHoidcHklCJWJ8iL9QDw0bsmBaF4byki88VR7YHlDw7UQxLXCZtXQdyOsa7w5F9S5WAgSWlpXF4HuZ7xgsEToaX7GmGr5TsfZ9rbw0uZENJbf+xtSNrI9zGTSMixwI6uOtoU6z7UrVRB6bQr04fdfUWzduJ8pNVxke61lSyPehyATFqDD74j5ZQdkVo4J39oUmcw+nN7Z4Cz9SyKuuV6oN9QiRRO6hBoJxL9/b81AUwO0rCjOsA1BGwi3hx5WxAuT7k2/lIhUSKCRQSKCQQCGBi5JAQVhclNiKiwoJFBIoJHD9SkDA4xtVe8gKM21nyQRIPuzqz227ydfc4oZuTV35xkU3fMu4lDMPSD0MwgAQCECNxdSu/pZjANz3KANcm4slwHFz2TTo9sjM6zlmQBSgOMmAawApFoaArJTR4l5wzZQy5QUuBQjnHI5DGgC6s+U42mGcx997lVmI8RzAK8pvABfvUYBBA2K5xiw2AHdN65nyUQ4jVZADMgP0hxAABMbNE/XH+oDnUB8WgpAQj7iwtsV5Ny649p69Lpwcd1v++wm399dudfE0ZcAyARlzP65l8fgqtVVXwPBFu4fqW1lQNuqH+T/lhkTAooJnQlBwjEUrcmDfXLBgEYH8Ab2/ogwphKwp54PKkC2DZBVlpv5GDkHC8DfJwETT1jtJUuD64DpMVBpZWt9lSz8ygqAbep32Wv/h9Fi2q3MovrURum4n9Nob93RedDByi7jCmR4JjuxaEz6542B8+xdb2Vi6Nnzy1bKuGBYuecT30g3ylo1o6ev0SdwNMVYBy2ln9iGeSLTHkvob7WVBN7mY8UCZbLwydih7onONuOvd4GIIDHu2tLtzxa0ot7vpplY7HilHviuF/lRTBEbVhXmkGKRpN66Vcq+8URqpGmjRCRcJEvJ2LeT+oeE4nZX+eEJ8bhEAvb51hYgLZIEsezIJvHhha3nP+FwyuauRDjGeekTeYur2zCXuw+tLvbkFi4p3q5zvUhnbxN7Q/l4dwyUHLtcs/Y52LBDqwOFrc/cccSSIZ9Hro/3+yVhhrmROp4/Sjy1WC++Enh/26wB8p86KTeFyEXvzof6RadUG/T0p91BlkRZdKVfX4iSNFfCjKzxVnvVdRYGBb4jTpKtoFmXNv93A9xcVrpf5Grle6wTPtTmAilpdsgT6ZAXzCt9GvPM2C9S/UcZJm8QivNDLsxdpHOlw5sY2ZG7tFIGwiRuReWEpC7M0cLUx3EG5xsJR1+g03bqK3sZRacnNH5NZU7bskaln+bRsUTpo8bBc/jx/QG/jid4b5SIThhal+nCsOBleEncCWWv4sVxDxS2mz2VDZgJ1ax7AmiMUEYMVLN+qlviuw+KiIZn8vbatwtLiIhujuKyQQCGBQgLXuQQKwuI67wBF9QsJFBIoJHAhEhDI+GKd/8PKgM6AE8sxGipbn3TrvuNFbu3bhlzrMcXu3eW7cPzLLlqP6TuLGcB7SAoANxY2rHoAicgAn4CcANuA3cRFQNuexZhpw3IPlmCA2gD7AEoQALzHcM0E6MR9AGDYZwsYZVYKbImzAJjCPbkX5wOOY8Vh5vp7tc+qDFAW6wqey+KT53Ac4gIyA3N4ABqIESNOtHvKApJyAvaSWMRaWSg3iTpwnHuY5QjPpUwG8HI9ANodyve5oFx29d1lV5qoCh8K3fDtnjvxj2b98HD/POqFCysIkY1qsxmBwV/sP/NSNpTDApRTd8Bn2g3Z8Tyei1yRJ21g7rQoH0Aqx6kfQCxtzDkQH2xpd3P5ZKviQcsJficV7gWWZQzIjSyNKGMMGHGHnHrHI6+dTwZ7ISxaX269dX5L9MA+YZOVRjbphoPj07KkqI8Fh3ZOhvtekOZBp+w1FkOvW/JdQnv2QHRlxiFtbwQU4wgizwKy0xdoU8pDhsQyiwyzgrIyT+k3+jvkl92TPuQNWGD0Gvp8CIw+WO8Sxa8QiKNQBHlHcSzyMIy216shc9S6JEEWeafsC4pNknUVmY50/XBkbZBns12vs9AORkeSXn3nqnLhL/dQTu6huhAXVyAQN/2ZtsRCYnPgpZ1dtYcmD3anqkvpcNbNKrEsLSjb0idm84fett5Dnlh8Mbbfr/wRZNWXA8Hqke+/UX5XT4jOvVP5XytfSauR/qOvro3Ih1ykhc3/BvbxDjMru56jduXeOdc6WYE8qKtk0sGCQpYSXskLltIkLSWZIr8oVK+w1ZrcwpSkcC2XUYIv5SxfTmikG+6lWZq3ktxtDyNvVuTGoXIUHJSV0gmCeffvfXV1gCtcmn5Q88Gn9izNyIV8rnBjXIHH9QNq853IN+M9yj2rU42bdYoJcXcQlZ8rYkIHlp7y/XT75ts6bnxLUy6fxKbXc1efaMuKIexGVS+WS6hFz0sXDj5UbdTGW1vHt7TDqJq72cMyHsxlWiHbC41OsxKDpPikHoRSwQ5tn9tX4lhmFi4yabg39Ln5z7lLRhTWaqdXKVU9r1pP9H6ErDh5axRG8nx5DhV5qX3e589TxlKaMn1BuSv5ZCItrvv30EU2R3FZIYFCAoUErlsJFITFddv0RcULCRQSKCRwYRIQoAgY+VPKmLlb8Ok9rrpzyk2+5flu5MWx6+wbdiUF1h7aPaeYFYBqANJoXbMPEG2WAyymzMUQ4CXg905lADmAfhb3ZuxuoCzX8GzuAfFhmpwATRAZ3I9zWSRBhAAEsrIatNCwYOCApVwPMfKPyoCwLDAhJ7CK4Pp7lI1UYBF2g7KRGFgHTPV/p+ymSc49zZKEOlBOygSoy7NNs1e7vbqwoOR3ysM72baQFtwXsBKgGJAXQPo25b0igg67td+5wY28aJN79Gcn3YmPPqDjyJhnYsnAfSAIWDz/lNpunwBggOQLTn0rC66z2BGU2WJ2AFRDuuzv3xj5mCUKbm4gXGhPay/6ArK1uB5Ys9CuyMUWs6do3ut4T0bXiyXFCq6fEK0BD2zpJxAG9FOICvoHMqP9kT1jwVxrLYmUiP9+4V8hY/9IfEtS8+dKCrK9oKDayYtqH3hwyJ9pKabFZMlvzAQuOS5sErDBYscwdiAbGQdGrDFeaUNc5zB+jPyjH9CulAHXXxbPhTFhYxOyEpdglJdxQn/mfpzLefRR7p1KDoPWNCsSGP1A2QTczpvtbqwgyRV88SdJfkuc5ds7SVYTSCRXN8FSKQwqIjZGmlmednOv7kt3vNvJphZdsDUdilIZVwQCbmfkBmdehMWVBFaYS2m724T4iLRIWlW/oXHhLYjGOSEpMC8t/P7BPBFhgasN5pofUP4O1f/vRVYgSxLyggh8t/KPK9MHfk4ZDVeuu+413/tAMcQF/Y1+S78eBPV67X69AMp9UF1zeS5uwg/lAEqO8V1Z42lMWuFtSUaeazwhpLn+l9eaLC/3Yls4GTRlnjxI6ezQnxDZsU2B7B/VdcxFRvz0u+X1tenL1PpUUKtEuNzKR4bEAytVypH78Bf3JfVqKZ+Z47Xnsre9/IYrOd9cXw2yyrU9Q2Bt2pbvOb63diu/SW3+NVkmvFzbN0WVmgvLVQWvlqunSrB9jWb78lAgT5+JXD9lnfp45g2vTcI8i2XNkIfiACrVkWSyNp4sLh13jbCch/WJJAmi/MnF6dKmuBOtyVJ3QuPwmEgCWW8oXhlWDhbHK8/FJea4edM7gAynkD+lv3kPT51DJEbm7g/CcCEI651gLBMXGeR+2Lxj/kitnHQi11lawDJEE4D+Y4bIMxmQZNzfFHJ4zB0q0+t7hMryu/0UN5Kr3DTF7QoJFBIoJFBI4BqUQEFYXIONWlSpkEAhgUICl0kCBHsFkAbkAahc4yZe47uh2ybc+KvnFQS67MZfteD8ioCOOkC1uX8CjGMBD1g5+N4BAAWwxrLCQGzAVgveCfCB9j4kAtcDyAHEm592jgGMQh4AehKQFpCfawD12LfnsTVLCMpv7nQAfAFoWUwB0pr2OASDESoA/xAIEAGQIVgScL4BgAC6EAuUF9CW8pk2pQHMpv1O2QzMMJc5nLtsqfJNqxKOUX7KvKV/HI017o+8prUOfcB1j0+6rT8zpMDmd7gDv4eGNeXgWiOKkAsypu3eq3xRqe9+QB5zcnOpQvtSZotHgmxMU5n6IR+ei6wtQDbAKnUyKxiuNTcsJktr55OWFIA9F1XoZ9lFZ4lRQf2RLfLGasDcjNGH6a/I3oghkyd99qR7ll/YcCeAP9rUWVOun5R7/fPvFv6X9otq779vW+kr/u4KIVB6fRrQmz5MX6cf2ThkDEFIcF/GBmQV7UsySwwDLBkvADjW77kXfZc+Tz3o0xBajG3uCZHFMX6n7zylbLFLGF9nBDrkAsqXD/2yOk5FLm1GS6WsHgW+/GV47UgMRhiELYAVdd6KWIlQSOtwtx2XS5EXjoeSq++9bs7z91Wcf7/Yjs8LX6TMPM9k2a/iZdnQ3yGfCFKvEKv5g77LjkzH6xVL1X8sywOIwB6BuiTvIXHu9kder02Q73cr/5YybqMs0VeYQ/+t8m/0D0JY3E6A7itgMXJZhLTaNzXiYrXv+yy9n3gyvyWziZLeTMIoPfEOXlNkmca9bCvkkUYu7DXO84qsKoRNiqrwPYHwilnj+7EvuyY5jNqkd8NWXcP3QQf3W9cL6TPY5n2yohe/SbE+ZJDiSpJTTbFxfMkwFKkT+RWXyoUd78RWqRSk3W6WicCIt20cO+t8c3r8nmdpX3tWF3sFssKUN3gX8+31QuWt+mZ5ux+W5HSwvuw6SYGrZWUhcqImoiJ01bFpt3h8Mg/CRmN0Q3O+MpyOyj5QVoLfFA/hr6sjWRyV3RMiLJLKvCfXS2lan5g7PvOUf6IxV+c7lLle7yvv2zVOccu5fAeIiSyX5VQ2q4DZvGdlHhVpTAe4aTpX6umG+EG6W9Fs1mpMHxmazFIN92ZlKL63Nhq9YmZ/eSwIJ117cb4X24ILchkwrpD0utK7aDl+x4ckP8aGKSCdPJ3YH0UqJFBIoJBAIYFCAitJoCAsin5RSKCQQCGBQgLnlIDA1J/RSa9UBoRcjlGw4W0Nt/7tY1rHRC4Yit3oXeu0aPqMq0xtkusiyAniFuA6yfzqcx1gG2AgZAXgNSAmiyxAOUBXs6zgOYDjHLdFDtcDJhoRYVYSAH4WCwMrCK4DBAUUMJcrALEArCQDTg0stGeZhjjnWMwNnsfCkOsBD83NlGm3cxzQGFCV662uLMoMfGdLHVjU2pK0p/GubJqV1Ml+p/zcB1JokBjg/iTOe6WWs3Nu5K5jrrt/Vm0w5Vr7Mjfzd8gIawusYZABZBEL2VvVhqMCrf/P/j0uajMQ04LrzfXToAUM5QbERvueLb9ZcGyrL8dPJyHyATcGF1W2a+SiQesVI9nYAuYzpujzgPzIHrCCvs+YQt6Qd2zNWuVpRM+AG5hBTfKehv5phAlthIuxvcr0I8plLs3oy/RL+j77tCtjA+1S/qZsFmiTtud3ttyHODWQGow5SEH6KuQIBAhji/tAaOB6jXtxHvXaT1BvygDxou3JpH7joa0sP/sVuXOqyF1NJFICLVWVwxtRIO4NspoYlopoJ46T4VIQ1MNQ/VIIijxxdxeTbHh/M/MU0FrusGJd6SejUoruP/9yaz7TRswv1HujkOPDQ8FC9c6RT01+Yf7VT8wma2zOQrb7hP5wHgTFj/UF8IsiIn5YYKa5TOMw8nmf8r9SZh4gQWx8u3JPpbtIhQQGJCCvT5li0gdt7CUErMsUwGvItEJchKcI9PIsJwBU4wddahzXM1UrbIXcQuV5FMfyva87yMqipGsZ4+aS8boS8gBZEYWBrzktL5WjaJ3kyNhNw8hvuSQbWmzGdVl7zXh50hAo3alWwsVqOWJeXzp8fDF90ws2X/eWUM+SjjP4rsaK9BXK36d3ziuWCQpFTyqVZYWguNT98GpeUBZ2P+a6jWghTUoz1bG4MjTZJGZFolNaesvyPmAMkVoagNPqP3+uUBE3VkezqDrvjjXnwq3V0c50p1l+vVxI8V2wRsQEY5frNTh93icE3q6ncfe4mIpdCs6tbwbvvAJxa2zLmCJr+5oJpCvSCktpWBtVSCyXHa1P+l8RbVIq1xe+ZfZQOD7zVKUXkFsGWi7vtpwfqa4oB/RcRvUSFlk3647v8cMIYuMjKtNCEc/iWdLDi2IWEigkUEjgKpBAQVhcBY1QFKGQQCGBQgJXswQEFL5W5SPwMwA6wPw+t/bbt7v137/NVaQ4ncyccMHkiIvGYlfe3JEWF2CmadGjWW3unwywHgzWCwgP2cCCnYUamsO4QGGf30yD2xaHgCHsWyYQMOSBWUOYc12ARq7FwoDfTJN7QIftFJczlBNw0MrIfQBUjUgh0DRlxJrDgFTOwY0V2uDE5zC3N9R30KLDyAqOW7by29+m1c3WAhqbOysICrufnc/fQy6odF1lZ+Y6R2bd2u/Z7Vp7vuaaj5rMACctiDdtd7fa8iEBvj1V+otNfdKCZ5hWPbcyixL2zZLFAHNTvRt0B3by8deLqyer8FlcPiEnc6lk2rYW0B1AhD4M2A8hAHlh1gi0BUA2Y8fa/qzNu5L282kxI2g77kVmHEBoWDsamE9ZjYziPEgKc+PGJbS3xTmBvKRfG6ECIcjYwcKJY1g5cS/OZwzgNorEMcYVBCfPI7A3MiAuS6//CTgNpfFdabVTTwCqsEKv1Owk49IGn5CLm1I3TerCUKr1erQgP/sVObeQTmgQT7eSqJu6UjfI157I8xeELe/JkpcdCgL50ErShlBH4liklzn4NnKmjpAQuwX7bDnU3f7Vf154+bqDnal/ob8Pi8RAJsgoVllSlen/0f53Kr9EGY1eSOHH0cDWb32x9cY92rT39Q8wh/+0fv/fuYedVGyvbwn043pAFseynJjLsqxTLoXzAklHFMuipsAVovZwA6V4vz7zOvZu+kP+o3RuSbtpHHsjimPR1H5ZZkG8L3lXGll/zQlYxMRKdbLvE08TUEUynBDwOyGwdq3w3I1idjIRp03NLevTONsYlMKnkjxvdppxs9GK902OuxOyFMvkPqr755/e071pag3zznVhWfgs7SC0N9+nvJ95X71JmdhCL/flKM2HEVe0+iwtibSo9iwtAoH5Ig7ypBt43VY2VBsjfoVeT3G05Lnugub5huZ7rGd5r5OrfujWl8L827Q/LQuM9timxlRjfjieOzyy3Q9yXE/1k9fJks6CXFBFoizaGqU9t5z6c4uGLOfwruQYfWpFU4jeaV6+4AcyAyonn9JZ9bCUTE5une3UxlpBY7ZWEz+5Q6d9ZWJbe9e6GztLT/1zNDq9LxhpLcigI2WCUOg6hVnD6oL6n0x5Pi5K87e8IEpF5Pyljp/Xd8qztG8UxS4kUEigkEAhgVWUQEFYrKIwi1sVEigkUEjgWpOAwMFbVSdcEX1NGYuFO9zw83e7sZd2XfsQhuMlV5VRQ560RV7cr9/R+t7blwPa3xAcLOoAHQ3Ixmc7ALqBdUY2cBnWCmgkstox109mPcHvZrnAc3Adw8IHIoG/cQnFdYB1gKcQI4D9n1R+qTIA6ekggC08AYQpq8Wc4DjXWzDjKe1DACADFqo8G9CVZ1NPzgeoATy0BSEgPu9ZIye0e7L85ieY39gHRGQL6My+uY6y+Btca/c1SwuODUmVbsGNvVwyUltg8fLku9FON1/CEDEQSLQN5M2L1KaHBfY+xMUXm/okgy2sz3obgTb8bhYUF/vIa/U62pQ+YnlK+/Qx2oxx81xl+rj1TYB7CDKL2wJCTTvQNwe17C+HvGzs2Di2gPKDz6LPW58edHFm7s+op7lNw3qCsW3uowg8zTiEkGHssd9zZ6GMlRB9mvGA67M59eNg7+KHkiPlN6cCShfLJb8rF0r1RF4zZEuRqhRNXdnVaKqFhA9O86pfCoBem0k3zQUi1kOXj5cVfLsS5FEtzHdnnmvVS4p44fu4xWJOWXVg5bfvf+ugvJAV8xzP2afy726m9a2trL6oIOijArE4l7JgmUK/IDG3vUcZwgJXUt8mIuK3TgM4aaMHlf+98r/rX/fr2uJ7A8KnSIUEehIguDiBt0X08d58SkPn0TDwhkX+xV7uqQ/2XpqxxhjEhdxDKTq350n7WyCpy9rSHo9yebeXT/0hjbdhzUaM0fPS5r7GmsCTS7papJgeypskv5t6FiuybpTS+ljghbOSYV2T1Zhc2A3phaiYO+legbwnFHMHsjWqlMPpybHawvxi27sCZOk1Jv7LXx1cF/WDawP+Y9nI9zEWgHxfvkPWDa5Uk+5OzxWUXkHyCQZ5EZYqiUh1vcdEO6hDNOeqvqwjRLS7WVkwpCIJSqVaPF2qdfmW5F3Oe4/vWeZ6xtIxvQl45s3lWmfj0GRjq1gOF3f0BtNLS+OxrKDek0T4XnbbKUsoWRrqb4Yv7+mPK6/oDkpXUKqvluudcrkWN3S/o1G1+1C53r1VLqGGo1IchZV4g6w9oupIZ++GXQu3yUGULD/SUnnIm07+oXRHqVr3FdvCdRotlybd5Q9eVa5nfdFPmjfWZS7+gSiqffalb/yXhz/7t79TEOeXv8sWTygkUEigkMCzXgIFYfGsb8KiAoUECgkUErisEgBEBDgFVNvpwtFFN/qSta56k4Jrr5d36wnZvg8LGBwF2AdYBGgEqARs3NtfLL1GW8A2QDlzYWOaXhagz9wKmWYm9wHM5HeezXHTtrY4FVhXkFjIvVgZLTL83vN8FmmUiWvMHdSghrg9f1DjDA12I1G4F9ncGrEFNAUghqhgUWlWEdwf0NX89Rs4O2hRYc85XfOU4xb7gX3uxbuZOlJvI2hsS32tHgBDgL8Avw1Xv7PsKltVxu5x9+R/gFCh3ZAhYDdkDUAwsqFNL4mwoBDnm66XGBTnkscKlhWMF9oQtw4QVBB57Fu7Q06wT5/DPRNtSh+jr1lQa/pob+ycZiFxruJc8O8r3H8ld0lndKGk+pt7sB443++LEHz0d0iIHcpGxkGuYXWwR5n+zZhDXtanmRfWbz36M8fK5XulFrormi6/sSQPGc0kzTvtbuoLAJQyuHKG2qesFDzXEYgUJGI0kk63Ws2CEJ8X8sTfXFRg7txPKzMu6K7P3DGpjjf+f/beBMqO67zvvFX19vd670ajsTYBgiBBUhRXi6IoUZasWJZkObZjyfIiL4onmSyTxJOc5Bwnk+Nxxj5nJonj8WTijLweL7F9LC+xZEu2tStaSEoUV3DFvjV677fXNv/fw/ugh2aDBKCGRBFVBxfvdb2qW/d+d6l7//9vkVsc5o4NtVEvW3gb30DetCdzInNP1LeoGFKxZTHjMYdB7G6Rj55HJwQ/veOLKz4WHwIzP6Lzv6b0o0owIL+utLTOyoLy/4GSERaU4pd07w/pumsRUN6kZntVZiMvamldpEVbg2ZZs8lZhWDAzVpXAGugt6Ic1fsyXxIS6slBTZp2Res1gUNxoqZo3GNJ6h3Sn/Srq+1G7ZXYAJ5cO0FOVETk1ERcDCvUx2y5VGgqfEW+3u6OCrcuiUatdMNkSnYppUKRcDpppDgWayIyWsv1tjdcKR4frhZfEGnUUpyLusZqN7O0eOU0d5+sQKmF9xBk8duVsAZ8J5YMuD0SOeHyJVlUyB1UD7RPktVzMcA8iz3Vi/fQbeYrSydGd0ed3KHqWPOM+s5IUIjm9Fbi3cbcbetYvbf81TgMgk6jcKrbLGzT924a98iInvsoWS/U9Zyuni/LHo91Q+90P7HGYH08qOjSM7zokRVeWtfnYf3ZFGFSHN26upwvh8+0Vku+LC1KIjBynUZRlhPhCZEsxGTZXihHJ/VmnK9NpHuuu7v78U4jnj321cr1q2fk2yrKubAlB1JRIvJCViY9S5PzLqLeJJl8n+79VcmykbmGeuX07awkmQQyCWQSeKVKICMsXqktk5Urk0AmgUwC32QJCGDExB0trxuV0DYuu9E3KoTkjQrPOS2vKqUR1z19yuUnll2uAkjB5gnAHTD1g0oArW9Q+ltKgHIA8/xuFgemsT1ogcB323ANukFCGuZyCTIDzTNAeIgDQN1PK+FWBhID4JOyAIY+qfSu/rn11hUmYSMTTOOLjR1lt1gLfMfyg/LjE9604vnkb4BF8rBd2WDAbXNBZeeMeBg8b+Vgg0odkR+ED4QLMTnMlRJ1Np/2VmZzT1Vz+cKq8yTmrT+xy819qOsaT0FK0H5G2JAnMsvRtgKgv2APzj6/YRKwvk6fBYSn/wBK4+LpISX6M30DF0C0N2ADRAbJ3CVRWIiobylgcIDwoD/i2ok6UF+AHOrKGDYyg/MQFQAt5hIKUgctcMAcxuOeIF6qTXX+slnIz+2S8vfUfPymStiZGFe0265IC8nYa8kH/6Kc8OflJz4XhmHeS7tRIPsKuYeK0CKvS0W8laaVOEq3yhfO9unQ5UeENSn/9eTi1egkRsIwX80R6FhBt/3laGJWIQIOS6l1XqWQ9xgndxyufMeQFwnENK3Z39A9t/X7y36d/xJkxmBwXp1j/sNdya/0ZfZ9+vxlnf/0VXZ1dTVkleV5lSWg8dBUYOg19bnn4iQu6W+IuzSf92M5x2/I3QwMxYSAdqGlcgmFazaR5bquq2G0rD5q8XM8Yjq8GgNvq04vagXq2mpH3vhIOZ8PglyQ82pdj/WHwGfPH5GMpkVgoDigSNxeQUrxFZEUXj7I3eJJ81zkxOlC3kd+w/ouctU7IfdQzPeMd8b0xdYuV7lHZNmbBPpkBWtP1lC8ryEq7lBSh5CVg3i8IJ+XAV/Us6yArNDRiMPOM/rN1z+5e/J4h/UOSIuwnXPLp0a6c89P/teRmdX3iojIy3oikjz1UlgAACAASURBVLunUETC4yISZJXjdZsr5d0rp4e21udrkYiOQmOxUm7XFT9CHYlD+dd4/tfyxsLCNUVesM6wtafFnOpdJu9MIiEiJ7JkQdYVaWmoc2oc908jrbv0vLtPPzN1Nl+KOtXx5mzOj+utemlCfH95bGYl0b27Vb6S+JmxLdfHHREmx8Z3RfNHHi6+rtMou/piwSkwuMiK83GurJxFxbC4OenE36YTuIlE+SI7MglkEsgkkEkgk8BFJZARFlnnyCSQSSCTQCaBF0lAYCIbne9XAkxlk3UuMPW2v3uDK83UXHdpTfigqIKJlgt6imPmLunL+o45O7EeABv/bf/+9eSEaS4PWjrYhmrQXZKBhmaBMRgbwoIBcx9gP3mhoW7ECODnd/TLZv57ra6DAICBk0YicB95m5setJ95BkSKAcVU2qwxLNC2Bc02zTaeZXVZX382lNxn9eLZ1AErCL6bdQfkBflSfp4PWAuhMpifub8aVtTDuivsqLoDv3m9e/R71lznpFmYcA3+kakHMvp+tfFXBSLzzOzYRAm8RIwK2oxxBekEqYZLCSyPLAA9/QxwnrGEZQH9mN8AuvhuAc0vyRXXJlbpamVlFlGQoRy4PUJGRlAw1ixOiskOudF/iXODPPYFyar8QD09LOuJsiwq4jR/z3wpt/VQvZXb05Zf7VCgiQDV4XqzW4uiMAm8uFzOh4mfd2EjyssSw/mKONySicWq3NpIhTRl7DMGjSi8WvWnThYzR67bvOtdErRHgqVq2W9vVQiBmZIwH/qILCxGZ8ven94+1Jt/6AucZ679z0q4I2HOepE1SN8a43P6DXAIkofjF5SYFzdy6XW16prl+8qWAP1J1hTpaY2HUqrgL+pMFbmxEc6eTASpJ+sfrxaHUalHaOgaWTLpnDuNZYb+PqnOfEz3M3ddTaukV6QUR4ZKvgQFW1FV/IpRxc+RZnrktbrpbslH81Ra6oSp5vck1DW8c2sS+EhO2u2dOBFs7Rr5fO5UsRAUu6E3VCrK1kVufnSdrQMywuIb1PIiJjZ6En2a9oCokAKM93ZZGtwrpkDEQs8lk/NyBVlVlOUSaqhHXuioi7Q4KfdQNf2q9RdWc07z/Hmlk95z5F5p+4knt+5fODZ2qFAOR7fffOrxfCk8JAuHqVw+frhQ7bZOHZz+cVlXbGkuV4YUA0N9Sy+G+OLDTMXRus8zBRjWi+Zy1FiNUM9IRE4Etcl6W6TF6PiO5a06t5XYK7yFx3cu39peK+6W+6qa3EGNtptFyA3Wo3Oy+KgFftxziRoErhinTpYhqT80GZZGt4V7x1rqw5W8O/54MZCbQ1GeyTkCRxHIFRvn74qtYS3665L1nyEnWVpk7qG+Qf07e0wmgUwCmQS+1SSQERbfai2WlTeTQCaBTALfGAkQ1JVA0gDzAIk73MxPbZf7J2kMFj1XOxC7NJYu8racIgl+Ur+ze8Lf/qH+9w/r0wJnD4L2g9YURlYMWh2YOyVqOagRZsG2rfYAv5xjA0V8DZ5llhDkgfsmNvvmPsqeZQTI+t2eAQK43WGjB3gMyA9ZA0hI4p3JM820Hi145GPBh9nQDrpuulhdqMMF5vn9SlFetMwBMQFlIYmwsuA7mn1oo6GRv74ulPVc+fycyhM3XWVf1d30/wXukXdwrbmcoj7H+7IBCKeNf6f/7Ozj6kjArHHoI4DKWLnQp2gTrI7oMwD2gPS4mOA7oAj9FoADiwL6tVnvvGqAq77FxXnLpAGih75M/ZEF/RV5QVAAkCAzyDtcSnGNCIyklU+W4yF3MIyjoTEvjUaG/cnFudyNhTOdkWoYFsZ9F+RavYDBcU6BTH2BiquxnyuHPUzQ6wWQl75qezWMVr+45C1Nl8SCCJHR+U2X9z+5jZijzimWBeN8Vs+HhJGbncCLkmqyEk2pvvmwprgbAjQXi77mIc8rXFd2pUbsStWg1xeQEWX7qBKVIA9kBOG5/oCY+HdK36lEP0O79QcJ3p1pbm8grWvzlJHvK0mSPivQsinIvC6N/2XphtdkfbQt9uIDukgRLNJVERN696V6T6bzuqYXT0fnTJO756bu1WhdcbGusWWi6jVbKMW7glzObdPc4Sv4dh33dImMuWrlAtZcnVZHOuq+a4sUCiRHAcGyNAvTNQHCw+1Od6QbFRQzpCdHQhQcjqKkIpMMXMCF2Vj9pg1M3uHMm3yGmouxa7gX909y/ZT3AwXYVrwKfs3li7JcKJ7yg3xZb5tVWVpY3CXmaN5dPRdO646aCID3tlZKzymla/NVrrlLVhb7Fdui5PnJMY3HoNvKF3TduKwqNsqjn6UIw1TrjHNkF2tGc1MKUcLRe5+po0aKOsN69rCsOk7Uxps55buttSo7xGIox0/xrqHJ+rCuq80fGV+T2yq5LfNXO/XCgwr43R6eXjtQyiXT+h1bxCDIu9dWRtPGtgNxV96fjnUashsK3cTqnD+zeKKgrQLxLPp6PPrQV6y3jyh9SelU3z1URlp807p49uBMApkEMgm8ciWQERav3LbJSpZJIJNAJoFvigQEHLLJQmsXl0JoQr3GlWc9t+W7t2lnlrhgSJEEtR8KxlZFVuBbH1dMEBR/oYT7kXcqYS7PBs+sFs5vlvRlvQVFbw81cJ6NC/fZvfab5WH5AtoBZrKBs+DX3GPX8xxATQBgOzdYpkHrDs6jyQ6oj5YoWvCA+mz4IBfIw8oDgMw52wyaxYNprw3WZb0LqI3qYiQKMkOWDysBMhpwy7saIojYEwQkNx/H9g6nXJSBfLpqE2Gv1WNu6DU73eQ75t38hy3IMfdBKgH2YgFzn9r6DwUcb3pgYeV9zR3rLCuMmDNrCvooYwXQAvDALGb4nd8A+SwWCv0P12b0M8DAnuunqx2j4pvdYOvql/blyfiFtIGso98iV0hCCEvkVRYJQWzqWDHni15QGCp6a9vlad8f9ctpszC7y0ur5dQvxbKpUIzbcK2UT1qavxqdsKkYFjkv0tDpxF5uxQum0yDwnusGU4+1gxN3a7RcZZBQKI4P2bjk0uJT8h7zOhdOtFqdXd7OIO4IFzslsuLYRM6tno79var0RBR5Uqz1AZOZa8wq60F9h9xEJi8iLKiDAE/cjb1biTmaAxdRfIcUy45rXAKQC3JrZJaKCqKdLglUryqmypjiQfPeiAUySmNcI01u1IR4MjdBKJ7SgJQ7qN745J2Fxdg1BzwWFKUcB1kKSoFufXF8uDK21uw0FLtCDKnf8gNpeaS+Xyp6MlmJxzQZDemWkmQbSqQzoUwyVurhWq0Syi2cB/kTCjoW6psqkPfgEuoa76jfnOqzzppWwpriLrXPW4lRUayNaKmVVziSTs8VFHh8UCiEQa4w5AdBTScYE2YFfM6l6rl1GmTC+mNRLqKwqrxbBMK9+sxJHWhUo+2t/euVX88V1cscMmNQZDldxPrC4q9ZB7L1BWXZLqOHVG6ofJEggWJTiGjQoj71pnE5BTEigiQUUVFRzIxQv2s9knpyX/U2BeZuD03VT56L591bj/JFPVuVK6crQeSeVAyLTzcWvEZ5NPy59Fg6kxAYnKmDS3u3ieg4txZFgYM1tyfSIrO0eLnmzX7PJJBJIJPANSiBjLC4Bhs9q3ImgUwCmQReRgL/Xr+jyU/8BDYk827ye3a6oNrVJiznms+ccsOve1q7NX4HQGSjhbUBgBhWGYBwg+C9PW6QgOirW/W2L/YuGrS4GAxEvZ74IL9z4Pw5coE4DRaEGODO8gZoYUNkf5urKCMROG8xNSgbwOhhJUiQk0pYNpjbJp5p5eN3vhshQt3ZJAIus7E1TVPKCBBthIbdv14OVh8IE7TIIS0GXUEB2t6sxCav5/+/X0bAIXN1RZ6U49wGOchLrW1L5Ma/PRBhQRmoG9ciL9qNOvCdtv5HFCA7NlUCtDl9gfHAJzEo6H8GNAMsW/wG2g7LHgAOPgEUzMXZphbqWymzAQLDxmkPCBWRQV9mXDK+AUmHFJcin08W/Xx4ct4Vdi2XvbVtSb5TGS3WVoodd9rLxeW2QpJGURQE4WK5GY6Vy37+rBRio7Y8Y7QTr7Xq5Q7O5tInvtL1cn9wMi7dPSyjjKt7UC/5rQ9CFxcmvaQ8FsTl4q5gpZoETb/rDwdS0d4ts4vcHeWgeGPJb8jm45E4cKsKeEz/gtDkQFMVMmdVxIS3EcnSdw2FW6jB4wd0/S/qt8sCmEsfYpq64GCe6zWN0uD3Cy5qfy9TcXa8UiWwjrQoCizvCoTEwon3DAQF7xfauOQSuU1T0F0B6yfU5KE+5/rXXZPB3CvlvCsV8gXF/ais1ru1Vie8vhvGNcWpqIVJVGi105qsLgoiGrvS+ZCVahqGieITh2FO1ivlIO83S15Sk/nKCXmoW21G0VC3G1ewdOl0o1Qup0yp4ZXafV4V5drAHRTvZtZdxAo6K1dP78+VKg+Uhyd6wbU9+UPKlyou6sgzar4Ya9kVyvLiXAw2r2c5xzuE9zzvfRQWsKKEuFg/GdK+kMqQEuaOdFijjXU46z3W4ZdysNZjrJpbw56rt/7zsZRmbf6cyJEwbBcmRUrUR6bXnpfrJ9YorxPpUiO2RmOp4gql8Fi3nS/pmom4G9wnskbWJOm8FyTPFSrqvefmet7B1I06Lau/npTBSVqspe3Zu6MdsrR4Ium6Eyeeyt0VhxcYKyJX4n8QR+2Xlf5K6dOSP+/zF72P5DLqUuqeXZNJIJNAJoFMAq9CCWSExauwUbMqZRLIJJBJ4EolIDBwt+4FoGCT84jSnW5MSl5Dd0xIg3nRRatllxubF3nBZuyx/uYC8Pv9/Q3Mnfpc7xrJNtsGZlncBiMrbENlQP76d9PgTod7AeoElPRAd9CzW5TYcFnAT8BgNmyYxPOdT/JgM2eupYzEQFQ8F7CY/GaVIB4og8UW4DtlZyPFbwD/lIFNGt+pLyAqm1A+eZ7FHHipuvBsK4dp5GPJweaU2CHUjXqibY+LKzabRlBQL8pnMqPNrJyUbVyOlI+7iXeNurE/PeqWPk3w3TcpsWkGVMKK44BSgzYXOAzomR2bIwHahLbCOukmJfoHCcCAvoGVBaAC52g3tNyxZrIg1Nc8WfFSzaC+ypgJ1W8Zixxrftouxl6+Uo2fGYmjWmfNv+FEPS62ZDexXMLTUzy5L4y8cthNhmrpcnUsaDZz5epiQ/xF4orPPeW2Bcth8cSp1J1+ru1taadu2z84mDLGetYtm33IHZQXrdwU+KWzpzw/nlF6o5/UxnJuaiwfblMM08KWmp/kJv24ILuQ7UNyJ+OnuWn5wZd/fKnGFlOFEA8avq9AyOfmOOY2ktcPyr1RkSHC3qf0u/0f/4U+iYFxScTMOqLC5iv6MH2dPMyFHyAW/ds0fK+KDDe7TbL8ehJgbNFuvA9FRNCnUiyaINIreOrXBVMiKLbp+4p+1/supQ/y3gNY7VmEXUvuoBBatVxwvvw7tdrhaqebLGBwobEpr1CCcBNXlv/MCkEpEpEUsrZYk4lqO4zigsZwKo9PcvsUuEpJmvl+UC4U/DGRHSO6viMrizCf82mTNm6h+u1zQVcV4Zh13U2SwCAw3g+yDTHMvLpPBMRPi5R4U2loTJ43871ErAqFTVLw6tJDfq6wV6SUrI/OuX3S2DBrWrOSPKTTWNEyH7J2pF0ZZ8SyYr2HIslhpRuVWEuifMO1ZuX7crVk/uVdwLqdfGeVzA0oz+Uc6xGsoH3FwnBnD03MrJ2t3ShLimBk66osLQInt1BOBIUsSDon2vXizrAl3Ze0V47FIAwOlYfbXwlyMXWk4zHvs9ZlXcO5EdRlitX03YVyuhqH3pHbvjt8sN3wfm3u+eDv63eUi9Yf/7BfZuYR1k62P3i5+ma/ZxLIJJBJIJPANSCBjLC4Bho5q2ImgUwCmQQuQwI/qGsBwnFb0+jFRCjt2upS2b07b9SV92gnc52UAANcCrFBAawCzGCDtZHW2GD8CtOcMndP/DYY54FiGjmx/tPIDnN/xCYOQJ/NnQXmBTwDjGejZ1YZpvVrABubItMM4x3IBg+ABu1Rytdzat+vk7lKIn8jB6gzwJ9tJo1A4Xe0wwYtR9jMDQb7tt8GfTxYuag7RAXlZ4NrMkKzD608NoVosUIocbBZ7JnS959hAcEpM5vsutz2T7jSbOi2/vAWt/KFG13S5Xo0/smffGhjgCbanEC82fH1ScBinPAJIIHWO+QEwY5pT0g1ZM44AdSl/6LB/JQS/c8Cun99pbhG7l5ngdFO/3qtszb01pVOt3Aq8sfyrahaKfqNqXxudbkd1Jbq3UCgSntyrLgyMeW+PBYkfmXFjQdzyW3FtWj42GIyPHc4ztdWE7loSd0NX15LsYphfFyVw8s1/TQujHleuNOPKzKp2HHatWZnCt0t/pY0Lba7neHJXNpUBOSGookvFlthZS10t8kfvicQs54LAvoX8Xvoaxact/0SAGYk0PNj/Tox1zBv/y2lP7mMCtp8xbxGP2f+x4UJxCp9mfmKOehw/5MYPDYvZsTFZQj6m3HpgJUFbcX7goO5irlpQnEYeA8xJmQZdJ7Q4x0KGGqKDpdlsfPNqOdmPhOrJvJrdaK23D+tSsP8VKWYP5Z6XmNtLd2aBnIWpUEu105+GCqEhedHebmDguBQPIuwFSqaTk72VcVgUS5zQhEVrWqp2JXyfiIAvCTWA/lfk5Yrm9lOV5CXrTWZ4+5WehNWFTkF1hZBId9f5qtLQyLI3+i8ZLVQ63whV0jfJLdKE1GnZ1jblsUC8x99xGJYoFjDHIk7SMgKDtYErA2Yz1EGos0tbhVrzUs5KC8KLyhKMDfzHNYYFIT1IXU4v/ZUzArXbcjEsJOTU6gkVNDvWN+H5ZKq96zmShklFqx9Wbf+hVxAlURURHIXRb7M/9TJXBBCakJaQIiggCHPha4TFNLDI9Opf9/7O82//Pfl/01mjB+6SFSo79A9H1dibUqezD3nFZWwfMmsLC6lC2TXZBLIJJBJ4NUngYywePW1aVajTAKZBDIJXJEEpLGMFj+gqpEMs66o2BWTb9/iCtNt5+fLUrB8XJszsyYAiOVgo8KGxTTKDGxnw2EaUwZWmasn7jPLC65ho2JxGAYtKgA/Bt9VZuIOyHuPEhs/7ge0MyuDQasFymaum3gGG382gzzLNKgJ/GeawgSuxSzfrETMOsPqQh5GVrChpGxsNk073lwvUSbutXpZjIKN/BcPkjrmgoD72ChTXp5Nu/A3m1/qysEmlPrzbK7nb2QAqUIdE7VZ5Ia+7bQbffM2t/hRQEWAStxNzSpZ20zT9gKAsQDIjkuUwLqYFeYCChCY9qRf0G64eMK1GP2YTT4bcVyosennE9djPcugV3uMiksU6xVfds7y4o+Rcyx//J07DmzryA6hFbWfXZN12LNFv131C40dI/6JPZXw8AE/DjVuxw8eTV7/bDNZ3Xkm2bmtkfgrGqi0CVZbw7IqWJArowt8WVxxAdfdKIO1ahpVDiTtqbyUcpddnFeQ0/ZEXk+bSdJSWpQ5hUu7vp94hSSd8iPptOcLa9LMrteb7skodgvFQhApmVsO5tZQAGr8ErE3ALD+d6X/1C/OH+v6oq6/lDg2Ro7St+nTaAVD3jLvAFRB0DK/0J+ZhzgH2fo5pY5kyVx2UTD763UZtYGrKqpoBIu56eu9G65Wm75U3+iXj/KYu0QuP29t+PXWf7P65c9V9rmfaT6LnGgvyou1DAd9xEBKUwSgPY1k5/NVbV2hsXIxMad5zCkKrhB4/mKj3T0UxiJ3PG9OQYhjuXcqiuApeM5XUG1X68SJjDA8xeQWzK2BHCZBrh3F0/ozFPHx5Eit2JUOf1tGGWvqLbzfX2pMb1bTZ/n0JSCAnH7OmhbA/j6143shmMQs4QIqVTDtQaUTWVp4NXmEem54qrmIm6VipTu+fHqYoA01/ad2dB3PT+dEEjyteA6r+mTOhrAYPFi32TnIaNxB2Rr7Ym1jwL7Fc2ONwZzLOhESEQJjMP7aBfnIciIVQfERJRRYWBcSDJvrOVAGYn5fUNk/UyiHB7bffOr0+A55fvJT1qCsZa0efHJQfoiOp5Veq3rv1IxRVkDuiQNvCT/z7Ody/6m55P8vis/Ri/nRPw7rc1bp/1JijYoFIO6xjLC5oMzZH5kEMglkEsgkcG1JICMsrq32zmqbSSCTQCaBl5LA/fqRjQdasr1Am27mR7fI/VPiknaoHcYJV7kV0AIgyszaAaYMsGezZBs5APRBYMYAI55vJIS5EOGcxXkwgMm2M+Rh/nJN65PNGOA9mzXKycbS/OhanABz4QSIxrO5BzKBv3kW7pAAWNiQodkG+IZbHhAJNKvRcjNigHs5zB2UERU9gLCft4H/kBT8znOMGMEygvKeIxG+BqL1sz1P3Fi8C86zebVNocmEcq+3SjH3QaYNiOUFZeI8QOIhV7mx4mZ+ZEWEBfIGTKQclvAj/FUl2j4jLKxFLu/TSCbkTTKtfPolB2OERD8ySwrTSL6mtJEvT6xXfnXfJU33I18+Ec8vT7XkAz6fePXaSO7s0kT8qMJArHVy6ep1RW/p6O3Bp572g/HKV5M9hcjVDHAHAALEAUC5GtrNgfPD7VJYH3FxpaQZ6k19L3JJPheW0m6SkzLruJ8PFKxX/jgUfNcl8Vij6RW7Ob/h0k6pUinsmsiVc2nqNwVsQkQwHzI/m3umFwmQeBUCXf9m3Q+36txXiHMxeH4dAUAfZ8+A2xKstJgzAazMpQlEHSSGBZBHjgBuXMN8hBwpG25RzJXXlTfwS99pcyFXMc8xt3MgH2TTUt16blquFnFxkTgfzOO8K2eVsEYxkoh3Xah7zK3XhpYoV5vQ0PNtHsuLtOhW0zjYH9e7N0dr4Xgarg6lEe/GQQUE2tYse6jDq5qseIku16u7LCiI+bE6XCvlmu3uWj5xFblv6yrItgIUu+2yrBAXCUzrycu/DgUuV1CL1BXzsQKcr8meQiddXgRGVeN5Sd+XGq3uciFfpp+kfUuOF5GnmUuozZ1G+mQFcx3A/08q3SZXXa5QGRJZURU54Zu179cerADUSep3gnyc7rz+7JnySCtpr5VOnXhyaz2N/YNyt1Quj7SP1heqp5eOj1TldmmfiItExAXzNus8EgpDzJnMobTzuTX4ue8b4TVYMrB24zpzNcW1rEux1KDfvKVfSHMbaGTE7+g860kCXz+g9Hkl1qg9d1aypqhrVfqoOmlHThMXq+ON4u7bjx/bsne+JmsM5jDWtKwlyQPLEaw3OGydz1yLkg3vhQWJr3P966PC5O5k7vkv5j524vHgnnbdG1Xgbw57d3ybviOPP1VCKYh11FVRFuiXNfvIJJBJIJNAJoFvAQlkhMW3QCNlRcwkkEkgk8DVloC0xQWYubuULM5Dy5V2lgV2T2j3IoCsu6w4FmflnZaNUW9TowPQx0zaISss9gMbJiMgDOAwV0Vscuzdc4GWWj9PA/StyoNEB4A6myCzamCDZXEbABUBUIwkIR/K8wkl3J4YWMw5CBc02Ni8mZYYQPJsPz/ICq4zs3yeAeAMGWHgM5s205gHpKZeFsAbrXqezybR8uB6kwl1M8sL01RlE2xyoS5ca38bScEzBuNWkI+5ogIct40toBxlpTz7XFB4yI3e+6zL6dKojnyoH4Cs+R8m/7vUB56TlvqnyDQ7LlkCtBttRZux2QaohQQzv9P0BcBa2vKwEuPL2vOSH5JdeGUS+K47tvcsLn7/My/EE6Pj3RvX/qg1Ej8lU4XW00G6enuQdve8LT3y+sj/jkop/dsa2zWAEjRN0RQFzEFTFIuLzT6kfR1LUzUcS7zOdVE4tC3veQsCMI+2XTgTx/miwJxKO0oVukLOn+RKJq9AHVLwFZiZ7i4owK9cxRCUtSzgK/L99LRATohW+qEF475YmYlj81tKP9q/AAIDEgL3Tb1jg3gVZlWBVdusEvM+5wCubF5jjjXLMuTI3MRxuxLzNnPgXyphxWaWBRcr45We5/mQtoBo5uaPeZG5njLw7qJPEBeIsXk1yKj1ZWfO5fnMu2hsMzcDyiE/yomcDiuZ+6xen71SAVzJfX2ygjajH/B5rOEF1301N3zwuaB6XOSFt0/kxRtD+KnzBDuyi0QOfkPLeiX1+wbc05vTiWFQLuVFILojIiGuE7QtCNspUo4/pHNFmVQsFHN+qdFOe3FepKjvleQcyqXeogJuHy0WCmuFSr6Z871mQbYatUrBYihkMv4GNOK6RzBvMKflFZ9iPlcsT+ZLZXlDTURaiHqSSyUSoyFfCglS7WbvPDZeG29sg40anl7bV5tofLm1Un5kZGblgSCXfJvm6mZ7tXT8hQd3n12br97cqZfGk/g8/zHbnwOYU83dJ/3KCNf1EmBOYW0B2UFsCNYc9CsGqSnLsO7md+Y61o9GWPyQvv+60i7VpaL3x+2qVztXjI4Rl0bBtReq482Hksg/Ob5jaWTmxrmhQrlb1LWsMyFVeEey3jHLjN/Td2JjUBneDVgoch3Xc+2DhVJam7wu3lkeSZsTO5NPPPPZ3NuXT/olPc/2E9SPd8RPK/03JVwVIocNCVwuzo5MApkEMglkEnj1SyAjLF79bZzVMJNAJoFMApcige/VRWx48H8LcDLrqjcquqtiV+TG6y43mnfBKO8MNhdsiCAuAPvZ1LERAoRhk2TWAGywjawAOCJAN5sqwFw2YOYaijzNJdL6e81llJEYaPdibs7zzBoBrV6eYxYVRoLYPRAxaGqZ6wo2WWzeAI8eVWJTBWBEflhYAMIAbAE8kyfEgrmd4jugIOUH0OQePgEIqT/f2WixYWOjRkLTzdwE9TQx+/kCRHBY3QetTWgHI0hMw4x6meadyYX7KQPP4X7yQq7Uh40esqKsM66w+4QbuvukW/oEsqM8XM99h5UA0YhJQh/ICIt+w1zGh/U5ZEq70WYW9J22os9Y/8s00Ek5iQAAIABJREFUBi9DsJt16Xvu39MDFBufvV3Ruc+c9dPmdZ4LmU/8qtdpTHlzpwqebBfSZFJ+1ABbIEcBjgKBud5ma+Kn4bD8i3TlAUbGHn6okBVekETVfJori5coMIgLcjGjcZy6Zqg4FgrAm0/SSqcdxq4Y4CpmtBslNQXxPTI85FbKhVwaBB5zQW8ORhv7Ym6h+lYWP6vrjLBgHnib7vk9s7IY1OZX/ZmPmO/RgOXTXPcx/0MOGNEBeMYcSdBXQKp398cC7wveK4wNPpmP0dbfbJcfjDXGIm5UaFvmY+Z0nodFHcSJnaMsQ6ob5El7s9tXeQ4eyIt6v6EvP+qNRrIFOzeLPAtujWyQ32bLZ12xzv3ZJyt45+EKEaUFPmmzauy8u1a93KNK0Sm/+NCn8xNn5S7KLGS+oSD6BlYrtPV6LXTKhNxeNM9eZQsVnteTh+LL5JNz1hLPe17RUwDtKMn7pShJcxrDicZusZBPJkRiuHzBj/TWDnRirdONaHO5ecudDWMF7k58+sf5d/1LuHnbsF2zk5cvgb51BWso2pK5o7feFNm0L4m60v3wXanWcZXRlmssVVwc+a461nSloc7Roal6WwTFXSKUd4jK4J0/qr/v1e8ndE6KP24/0S5yE407dt9+zM0fnqiffmZLvr0m33+pZ4oorIdZI0Ms8M56KfKZNQZrN3PFZ2tK1nzMyV9WmlVijYy1CHMedWJ8U8d9sgg5q/r4sv54YXJ24csiUypBIS6ObVuJ1FMngkL0xNBkY0RkBvMCCji8E29WYg3JWhqCgXmf9wBrZ8rC75zHbSv9l2ed0rfXytJiqDaRrE3tdQuFSvqrX/jdwuvCjnenfh883q4/IIpw1QqxnB2ZBDIJZBLIJHANSyAjLK7hxs+qnkkgk0AmASQgzXqAHDZogFFsnNhkVF31Nb7LVeRKuTSuGBZnpVpmMRLMHYhtkPgEPDCSgmzZvHAOABz3F7NKf6GECyIAMDYxBsiYiplpUhnRYUQEAIm5+QDU4X40dR/oP2fQFZW5jWJzZcA9G7UHlQBhIDDYVKF1BtgBYUH+bAw5Z1YXAPsActSJ30lswCAyIAPQQjXrDnMdZUHAAS8Awl5QYrNI/QxYwbIDrbTBOgJU8DfatgZQWOwNk82gJYYu6103eBhpxDnTMgako/xLarsb3dYffVKEBRrS5pqKZ2Clwidtv0RfkJXFV9blnf15cQkYMGYWFZBb9Av6GO5vIOs4F52LsZAd30wJVNpfYc5hrBfEFtDvH468oDEbHPLeXfizpd8If+SxRjx0m0gLxgMuN4xE3dS28/LCpJO8yIpI2rutIZc2k7Tp5zut4lTol3PSzo7l8L6l4BZ+IqRTWtktKfbWmt2o1I1ihbZwI6HcRAkVlRsR70tpNXXVciGVwjZj3wC3lyozffPnlf5Vvz3+nT4/0u+v55uoD2YD8jPnM08BRGGhwTxuFgvIlN8A0AxgAhQzEpt5iDHAvGlznc2tVyzXi1iBAJzxPHyxM7fRjpDIg/Ml8qE+5v6LOXnTyIENXGkhB+rLHA2ZA6AI4AcpRnk5+Bv3LRDpyPePlAACryopABnXl5O5+eJv2pF+dFgJP/YQPshnlvNyF0Ubno95YvW9yoRAX0zn25Fy0i8BbOmTlJFyMQ/zHuZdzzjfVO3sl3C/hMsmcw8pt26BSMhExKIfDlWLxShJFqMofU6khHhIN6p4zW1ZVaxVCrnI+V48VCscDTuJAnUnixrDTUU3bovQoOw9d1D9ZDLIPq+eBOj3rOfoW39H6Wf4O01jl6/4bmhqVYSFDGLkoW9oas2F7bybufHM2tBE41GB/s+ImLi3XzSzisjLKuGdOsc6GBKhqr+3DE/VO5168aQCW29TEOu02yxYTAfWnw/0+y3kAmtXztk8sb7mjFvmi0F3otSBcUEaPJiDGBNPKu1UWaujM6u/J3dVQ0OT9S0jW9dukkVFkC+HYyIykAHr1zldx1hjvmTN+4X+J/2SxPrGLDd4X0JoUFbKY5alEMiQ3ayJlvWGioamktPdhhcWh1wslaj1hAVlZiyzTmUuuiAA97o6ZX9mEsgkkEkgk8CrXAIZYfEqb+CsepkEMglcexIYAEwMbOtt2l8CUPju/ibEYh+wsTgl64qCy02NuNxYy/k1SAnAfcAXNjNmIWHAO4/gO8k0zA/3Nx1s3jAZR3OZw8Aj00y3vy1eBeWw/Lme77yvTIOY729WMuDf8jG3U5TRArzyGxqrlIkNEGWHREAmaL2SF6AQmznAjp6bi/61RpgAiHCezSFywEKDe4ywOVerc8AJmmxs9NgssuliE/dWJTarAGgAUyYjIyEgYQBZ7O9Bqwrytb+NzEADD7CN85Sbw9yv2PVGIHHPbK9M099Xck/9OFYlWIAA8Ji/e65F5mxI6QtXhbDYAMgzVzI965CrrOXcF9NV+aBv0Bb0GzQDDfxEptTtikHZq1LaazzTrpdTIFS3I3Z+KrJi11KuNilbh3jCzT12W/GLJxvJ0JHH6nfN6JrXi7j4Si1YWRPKAzCzmUfeeSlj9qQXtBoKy3tG9IN4CoVv9fKRJ58cYZLE+bwibsfdtU4c5/ycVxZDIRf3aUl+1BtyhE/k15IsK6ZkaTEmUPREwQ/MNZ5pwW9YZiwpBLD+kn40woK59Pt17oPrNLmZG5gXKau5ycPXOoAefzMXfUaJOfacJu25uZV3BXMacz55ADwxfwI+Me+i/cs8eUWA/Aba9jwboIy59oF+vpDWlIeD8gNio7ULaMc7gLIzZy8qP6wsXs6VVj+rS/44R/yfI0+IC4W1HQQKZA7vHcgA3rWUE7dj5sse0A8ZIjNzNXjJD73MCykH7ySLR8FcRTl4Z0O6o2FOOWhv3KPx7oBYh2yhbJtKCFjZLxIDxNYBXEYZ6VtofvP+RJkAxQjKzbuRtuSdy/vX3PBdpmgu7/L+mEJ+DZEOenbQ8LwkrFYK2xWk4nSiCadTjCcLRX/CS5JCV76i5GnrqMDwWCEQVoOcd1gcpAgLX1yF19J/gNW9d0tmXXF5bfF1XM1cxdx1v9I/pZ9BAeeL3Z4lxcSuFYUSGmktnxgvj25fTkq17pqsK+TGq7tHVgiMd8Yuc8vggQXda+LQ/225hdojwuLb/VwyquDVa0nih7ppbP7ImIu6F0AyrM0YY/Rj+sEbL1Inxh9j09bAF6v6Yf3A+o65l/gUj6scz4/vXHpy6rqFnXIFVZFLqwM6H8k65Ig+baxBJjC+eAZji/Uh6zbmK+Zy5g1bSzLumB94VzI+kSHvCOZdKsfaiDm6nMu7feXR9DNT18Xd+kLuiFZIvH8Gj3+kP+j7H1X6rNJmz80Xk1N2PpNAJoFMApkEXmESyAiLV1iDZMXJJJBJIJPAJkqADRTz/HltyPV5S6PetClx1/SwEpuNEVfccdRNfs87XTgvDcDSScWzAOxHoxbwatDdE1kauWAuj8ydBdq2n1BCQ+x3lf5XJcADu35Q63Uwz0EigDytDpw3t0iUY/A3ymcAMWXiWq7h2fwGcAWJYFpbPJtyGLDHdwAPruE7m0SeZSQB5/jOJopNGTI1F1iUnd/Iy3xO8ztgyQP9crKpY8NolhODG0zuZZM8aHVheQ5aWBjwDchG+TjIj4PrBi1UOGf+2jk/6YIhnkGbIE82oJAXaL/RXuTH5vQofULWAIBRV+swLV42r8iJjWy3r+17Htz/BmnsbkYdka/5wt+ovTbjGa7zgfPZWJ+8IN/iBzflMd/ymfziV//2RnWgzxf/k+afv7P86UqQJlMdP19cDqo3t7xiItLi+E3JU0cO5nfMFP3WG6M0F57p7tD4To/cVHlk6t6HP+BGcwtr/+S2P95QE59n6rdLkp2upf00htNamuaeSJPcfrmQ2ROmSVWBelP53ltNCq6dROle+bUvy8qi3QqjtpeXH/W8nHSIsYjjpKUgvwUBocMKzIt//BPFYrChK5yXKBRAEoAQMX44/qsSfsN7Lp761hXMnxAUZrlhoBNavcyJfJKYLwCVmAOpH6QugBuu5phTISvMtRTELXMOc7K5ULsk2V3kIspGnpACWH4wJ0K6Mr9RBkgBLBuwYGCs8hsWJoCL9IteLCTV97A+X/SuvJx5aAOrD4A76groB7gOmIm2Ms+mnDwP4oRPAEHmEd7FyAzLD9qH9xJ12FTisz/f8o6g/oCNPB8ShbajzJQFYJJ+dZ8SWtKUlXcc7U35Nr1cynP9QX+i7/C+GA28mADH+wWs3ifjhFM5L1qN02BWf7dzfvhc4OJUpONrBBIf0LlDIh0JTMy6ZlPlt0E5OWVzc09hQuTD03IzN6/xmffzXr6YeD3N8W7qDcv3W1H2UyeanbTZ7ISuVMgtlfO5hnzBmWudrrlou8izstObKIG+OyjGKeOTNphQu7nycOomZ8/pIhTL3lJlbKkut17tsW3imEphWqx0/XxJljP5mPUT8x9zHn0VIpBDNLM3qf74vrCTGxFpEfu5eE2Ow6QU5DzN6LNDU43iyumhon5hTckBAcz88B39vC5WU/obY9cUVy523Sw/iFRZK9Y6v1cZbj9fHm3lp2YXQgUIX1I95b4sZY7GKgILDOI3Uf49SoxxiF5IQd4HPJPn8Tvr2uuUmEeoM2XmHcH8gAyNjOVe5hLmv4pyOCy5fmXffdHOueeDf91Y9H5rg4Kz4mFPwnyTERYXa9nsfCaBTAKZBF7lEsgIi1d5A2fVyySQSeCalsAgIXAxQTygH9hoAeSw2WDj0XUjd+9x4clVN3xvyZX3AKawUWEzx2Ga8abFb5YIfJqFAiAW1wPSA84AwgB8maauvX8shgPgF4dZH1jZ7dM2crYxM4JgsDzmdok82Tyx0WKnaaAMzyR/c2HFJ4AZm0y0xagjZbUAreaKgfvM+oN7kJNtoMwqgnJwHWVAW4zyQfAANgFamTk+z+J+u8/AGO7n3GAsC35D9uY+xeQL0EgZTVbrZTYIzBhpxTPvd29JH3F/431c39FOpXzkj3w4kBt94QEl3MNczQP5UW7rB4N99RsBLH3ddROpM3hYma+47AOEBPkiDwOJjciiL3OePsZzDBzukWm63yyD+JtraFuz/khEaMS65oI5QeeuuLxXKsANtKetvnwOjif7u/eolwOONyAqTIaMWcYLYHb947XX1naHZ0aWgqF9W6LlOawW6n75+rWh3PunkxP3H+3seU3Fbzzsu/jZdlK+RYDocxW/jiu1p/QM3HQg90QExZXKjvYcVfyKchK0p7pxdVlg0Vo3SOIwKQbyHyNLilChKoKWNLVTT1YWucjvJHEyr4C+Yx3P1RrtsFUq+IsysojUoiVpZAOL1VrtcEXXXJIrHIGhXVlUQCIbYYGYf0rnfr4PlNqcDHiGNQRAHv2KeZ1zzPFYDTAfIRObL61rAFxBGPAb8yzAFoAVwBWkK0A5/fMlrUEsMz4v0nfIC4CNA0Dd5jzmOAPXkQmkBe8fyFreS8x/zLcAftSL8gIoX2A1wDNfru8NlnHgO3MbsuI9xPsIefEMwHcAPIiBI0rMzZDgWF/wrsACA9nP9sv6P/QJYLjZJDJ1BqSEyL6p/3wARkgrrCtoF3NlxSdkxl/1y02dDLDcDNJJ2V20fU2Ou3yX3KRQLWOjuZVGJyl1yn5zfCw//8RCuGXLajT6NrlZemvi+QdzXrhPRMWkOsLZotemr8buQ8traserYhHSK7yOvpUFX23e9XKBz/NLSZJK+UMLkogipKs5WUwVREKWCvlGJ1SYi1zQFFlh65GMrDChfuM+mZcZE8Rb46gxkyjWgpvYrUAjctQ3MpOEldG2N7SlcVQ/DecK8bQsFcqavxk3tB1rPxoY0L8hq4mzrZXSkPKphe3cFl0bKGZEWqolCrWeNLbsnS+NblvxVs4MKdLJznRtrlbA3VR/bDE2L+YKyqTCvLaRlRoEHXPc+UNGe04xNZKx7Suvl3VHS8/ten7S0SvGV/l4DuVnLv1+JazjWAszX0LufloJy6o3aJbfJZ5FhkHeI912/qOFcvgTOi+rv6Qg4oPnMuciQ94NuM/6KxE2D0lGN6j+zH/Uayp/Lgj37Ot+sHPsE79SOiMLpOl1qxHKYtZog1XJvmcSyCSQSSCTwDUkgYywuIYaO6tqJoFMAtecBIwMeKmKv0M/AoRgDUAsi8CNveFZN/Fds652Z9EFNQB3wBRzlwTYY6Ai+Q9aHnANwD9gjPmg5frPKQGMAXKci6nwtXgNBqCaRYGRH71dvRK/D5IXnDctRrPoYKNFOagHIK0RL5wjP7TAAIMoG+89ysE1gyQJgBzlImAgIBP3mRUFmyz+5h5AHDan5jpDX88H/bZysokEjOMaNnmAUGYdYu9dA6G53+6jfFzHp/1uALXJgTwpB3VmQ2puWkwm5Mcx2EY804C5be7m32q6J34U7WY2g4BmgLH8DqDGJ33iahMWVk4jkAxI2jRf8vaAb7FPIxtoM4gk+iKgAX2IfmguJ2h7gGL6MueRH2DJbP88fZA+D3BCnpHICsaBuR4j/+gz//ye5J8f+D+jR0ZQTu/1uR4Yv5HMrhC0vRTxD9bZNNyZN6gb6UpARhv7EBVYESEbtFW3Lge1xZZf3Nv0i/cfKoDVnjsEwrhcGLpOUhaacurOarC2LXX+jXvLT71NPzM3QFb8P0qMtTmRFz3t8sshLvrWFQC9s8p7VGzDattLmgJZn61HYyP5JNiK9m41p/CuvtdWxXtzkXw/dWRNMaLfXCGXy4eRHJ+nnlzOpE0VJh/LTVS92XW5XNAVYXFRi7oNGgM3P3+ohL92jp9T+kUl5hf6CP0MywDGpcUFQIP4KWm6n7yt9oXFH9jyQSMr6D8cvfbqy6UjwJ+5hjKhoU978J6AvDaXQmj1XhL5s/KR0fPvgp/f9y/db+380eLJ0rYd0mK/r5B2lwpJdyVI42fXckPfLpmOqk13KGFR8bmtndPPLeXH9nX84qz+BgyjHd7crytkBnM1dTRrqX51rujDrD6wlADopw9+sV9n5tgv5b3wUMlvLq3FI8znjHFAQWRE32Wc8k7ivu9SWpAcea9u6GLucsdm37qCdw3vO57B3MBzzYIROdOOzDv0A4inWSVIP9w70o7ntKW/Rm5cyTjV7V871tdD5eTZe2UpcbuIwzHJa7QSNLZvKZx46kx3+9Nlv/FuERh37Cy+MBEV8uPEpYnS/OtlIVUUYeGLeHz+5urDBw42b0PGT+7+9H9eu2/kr7qXM2YvKOAl/GFWESL+6PPIsafckKSpwGFPQ9Rv5oJeyIIh/b0iV2+t1AW+CAuuJ+EC6uuW5SUUNbvkQglAVkDMkX6In3AHVVR8oKHJVLEr0lOloWRRQLvWTfH1mrHOrR+93piElGItBfDPmPhYkngry6eGyesdYSu/xwuSYrdRdGtna82tN8wlQT4Zlmuo4WK1myqwdVvkhd9aKSsuxnlohvXZyx30L1vHDl57AVkhosAVyt1OeVihUfLxzuZyKZU7qLJIk1IU5kQspDMiZOZELLR7bqG8lDnwC5AxfXmYS9Rdeu904ygYqi9US0e+vGNq24HTz5Sq3QOqS5gvhY8rMYfOiag50mkW9869MDm0cHTsxp23ntw1vW9uhwgOcxeoZ7rbtuxNDozOJL+wdNz/j+teAryDsPpi7LLmzsbEy/WG7PdMApkEMgm8CiWQERavwkbNqpRJIJNAJoG+BFj/vwgAlsufnLTDI30aMIK7B8C3E660Y81t+wd7XH48cO3jB131Ru4H2OF9YQTBIIHAo/jbXCFBfLBBJ5YDm2+AGEAbi30B8AFYBeDBYSDX4Hfbt5jlgJEXRo6Qr21eKDebQgMojbAYJDuMrAAEMmKDTRXAGaAZdcQNCvUEvOE8IJxpuJvbpUEg0KwkrPyDGvaArdSbjSybLr6TJwflBsCjTAYK8WlAFGWhnKZ9zOYXsJRryIP8AAzZSPJsPrmH+81F1WD7UF+rC3nd6bb+iHwYF0fd4++BGKH+AHq0B8QU+T1L31Afia2v9Mu+mR+Uy9YgyMcscy4JuNzMglxOXhfR8CYLI5RM9ucJo/WxOTawpLB7jBRDAxHtb7k09wAUATxPSaeRTTtEIFYwyO8zSmiU/6ASACx94C1KPPu/KwE0098e7Mua9j4kwPas8m3GXpBvBpXR6c7pua2d6fxybnS1HZQYnz3iQuXeDOD2vHhfwrICUB7wkzkD8BpXPvR/QBfqDCFzVvcbMH4+zwu//Dh/mgzJjzFG/bHu4jzP+e5YKFTTe7EHDYGiruKvOcWs0E2Bu6Hy+IwCcM+005Li4vamGzTxGXvXKSEnSL1FkRAvU64LSskYHhOoWm8llejJ+p1zVb8x6cUlqX57J3Npfm7U8xcCz9sqEH6XIrY2gnxuXIG3V0RSKGZvpDnIC/3AFzGRW9SJxU4nLtaDjqffV4JcIE1t31MA7vUE5oYyEzAaCliFoDDCguuuk6whZ5jHZpWYF5l3DssFzyFpsb92snDm8B21zy0+MPZhxq5ZzVlcC9osklx6LqL+5fPnieq/1N/MM8w5WFnQxyHJ+XtJ42K9Zdjgu4G5zYA5Gs//yaO/5l3XPJz/zZ3vH3++umf45rUnG/mkO3O8vONALap382kIWXd8S+fsF79t6Yun/97h/zJ2qDJ78mf3/5v6X019x9s1DpJQfll0TQErGxEcsHb0eYiCC6w+rsDKgrnNiEbG3Sn1L/qfDGTSuYLfOfq9U7+x8pral3KtpNo93Lph7cML7/m9Rlx7rJuWIMiWZeHTieUeLE39swLiAfkY6xALL+pvV1A+e7cynyBXrDgoH+1zFPnShkqMR85D5vCOpC68+96thLxwMfhrtJ/KcNFYEZdLqCg/rGnow2URY7P6fEBkxaTIiiGNz3wrruyeyM8xBu+Q1UWt6Lenav5qrO/5Zlzdiks33ZdWg3plW/HoaD0e/urJzu6/yXvdQ7LMOKa+uXQx9248e5MO+lbPNRSfIiqQqd7lvclEnt0S2pH1SyiywtZWvTGgMfmiIrxEwO9NKu61m03fHZRZ8piFrUvVUu2655ZP+W5mf5zPFVLmNMYLVhOsdWkv1ozcw7oOyyTmJzn388aDXPwGBdbePvf8ZDFWjIp8uevaq+VKZbQVKyZGS+RBpOucgm7n4lAzfSGSZoGiE13aKsisLHlXvuQhMsLJ9VPRC9KCSAsFvk5nFGD7Ia+QDi2dGEkVALw+OrOyuHh87EgSe/MTu5YqceQfUXyOYyJUxKulKEq8WYTGiqxGTrVWS7MnHp+5Y/nUyP1yY/Whid2LbdWhnC+GeyZ2LZ+WAcbyoYd2T80dmni/4rPsV33WXvjS7t/Q58Mz+8+MyYUW8wpzTxrk05E990TPfOV04RNx2COQ7WAtivUf8/jvKPFeyY5MApkEMglkErjGJJARFtdYg2fVzSSQSeDVL4F14MAFWx8B0KaRBbjwvQLJBOx5D2qjf0B/r7rJd73epd3Q5YYLrnwdwATAvhEfAIiWn8WcMIHyNxtxNmvmIgIgCnCPzZwB0mz22Ihw8N3yo1zm8sbAlPUgsIFw5pKKPMwSwoK/PtDPn7y5joPyAKZRBt57gIYAMGY2D/DRUzHXAThjbpmsTtyD9hyEhfnppaycJ0/qbGXjkzzYXAGy8RwjXMx6xMgK6m51NYsK8kOTFs0yAD02xeQBsGEBGNEW5zxtQz13KYFw9MC3fp4GgnOOcpprFMDHZ9W2Lbfzn97ujv1H5MKGG/N92htwG7D3e9VX0LwO9NkjU9a5QNKpKz5sow34dW7z/zW3V5e2Vb/iR1+VG81KxLTHARWtrwUC3npub8wdicWaEEBrhNOUpEC9A41HaRMLJE7dVBz4uUa1VMlFyb2FbvdAEPVE87DA1duVuJfNvLmTWV8xQHqzEHpAgGdJ4KxUJ3NnG7nqUWmh/6EIix2fH3vdPU/X9gc635wIF74SRbkP13O1sBFUV1Tux1TmS3bXc5mStf5Jf4WQuVdpjxLnP6H0RiXGKeAxn5wDuKDPX8wKx/oS7oG+vd+nyO97lRgjL2Ipimm4oCDcecmn53qj4jcP7ygenj3a2etEVrjVeNR1E2nFxiNuJLd4t+bJu/v1BKhlLAH0EkD6Zd3iYF3RTYsjAlO9he50bj6a3nu8u3vb7tJzW+TJPD0aTS356WgxkHLrzjCer6VxKUqDSbV0UeAmkXgLAtDyciWjsex1PecVBHRWZXWxWCwEq3InIy5GDv4v/3hIt3xQ6QP9Wz/1E9u8W3/tZIrlFXNBz1+56j5e8trzBbnYf93wx4dlXUG/pm0gmpivIFohP2eVmONop2O/sPfHj/zx2fevfqV+78kwKdwqWUOuMUbWRMosDEVr1VvWHjfi2DSc6ez0ba4lX/qJubAj7+tFSgSzzcO5W9YeUx9N7ynHzeHV3Ih3YO3JlfsXPlsSMbC4r/7s4X2NZ4PRcAmAbPfu1lH/F578V15pf6fy4Nhd21dzw2HXL8xoPN2jcVHUmChvb59YevQTt529EndpvHv7QDtzLkTbCZVju9JpAeh3qnkET6YvSPv/S9eXn0S275CVQLS/8mgylp977M/mf1hMYo06ByK09ojYQr6Pt5PKuOI0XK/vf06eSl/vPGnvG+SOPHm3m+s02pJxZ+6JaOcjSvR3I5EAMM0FncW1svf511s2k2FRshmWZYX0271qJaiLrFhtaxy2w7SwS7Fl7hEhMaXvbZE7vkggP0mDSO6hEo2znNxFxTmve1bWFVtOdXa+W2THTcrrrMb1H4jgOKLxCPnIO6g3ZkRgbIoGtxGz9z6YIIf483f7yVfWXHw7b7lzBzKMRWCY9dggufh1y+78Uy7jS/9dxLNf9PxrJDYS45W16g8oMd/sxrqiUNaL+LrE7bg1OjM8nTb9XM9Sj77P2pE12N8ooTDAGgqFEMYm89QugfvKI51cnRsaDtuWZb/hAAAgAElEQVR5J4sEYkj03nCLR8cCEQaTIgQiBexOcsVQJHSi0R522/ViARLjEg7KCZH5cvEres8laLjcUWmqc36+EFHXebW2IjlFsyeemAlWz9Z2qpxvFHFSmz8yPtdpFJt77j7itlx/9qSotnFZVjwv649iY7E6pc9OY7l8q2JyTKycGX5/c7W8o1jtOFlaTHfbheM636wvVN6s/G8ToUFVSmHH+7G556Y+VBtv7lHA8gnfT1mzrkgeI9P74ltKQ+lXm0vemwfIGm5kzuutX0Uq+Q9/9rc3ZYxegmyzSzIJZBLIJJBJ4BUigYyweIU0RFaMTAKZBDIJfIMkwLZ5CBBaoMm+0OW3FM7FGV11+cntrnaL73KjcgU1tOqCccDrN7DZUGJTD7hh8Q4MnBgEyADUAWmwoEDTDMCLDRzvmkNKr1NicwVhYVr/gzszy9NA/EFAn42KadgakcGzyRvQgc0PG0WzfKBOBq7wPO5h80NdzMoCEIx8AWgoJ4BpT/uxny/XAdaQDwmNWTaJ5raJOgB0WtkstgDP4nwPhO5/msa9aVIOmvEbWUM9ADHI/5NKbJ55Ps9kg2w+15GzWXsAkluZIEkAu6wcVm6d6p2j/ZCF2vmOwA0/t+Ym3jHlFj7MefJGhoBolBFZsRmmnGsiK16s8kmuV34gM3OZ0dPkv9r+xa+8qBe9k3YzjX4LqG4u02gH/MJbYPHPCciijzWppwAi5ErbVdWDX+eK3pB60VbZPg1Fvv8D6oGVbil/5vTWiYlCOxyvtNXkilPgJ8mdClTgigrS6pJknx+qqWwLfw5u+oL+h3yjD6HF3pDm+J6uV3AiIpxc5Yw9Nnzr1HPVvfuX82Pe7+x4X2m+MGl98X4ByH9PwPRiKWl/PJ+Ev3zzb/6PRx9+/+sBLjf7MNkBln6PEqTFu/oP+fsDDwPYRoOUcWtEUF0yvACYF/hIHSD2AJRwq/OAks03Fy27gNBVAcgn82lcyckpt1xFRbKmmJX+q5tLt4nAqLsthZOKgF12tTSnJjhvZIUVzM8rMUf+Q6XHcRH1Uq5mTnRmc0PByh49896y3NV3u8WKggcPrURjQSMeObqYlp+puaCeS121kMTj8nkvgikSnKXJN07agR/UdW5YPvDb8hG12u5Ea8V8sFAq5V6IY3ek1QkTiI1Gsxu/5/49lwzs9GNZ/LLqYITF+FLUm/dfK9k86XnJqYLXvU2AcG229MyQCJ2lm6qPjAkspv9ixYObIOSPJR1zESQOcyNEMHPqg2+f+IOzClq+7VPL3zXUTQpbpXW7Q8GRnziw+tSDsnyYvKn+1G5ZPCjqbIe2ZgxBfACS893mOJunbhXJsG2uuKWj9G7147qIh93Er63EzeU7lx+uruaHd023T0c3rz1xiwiRO1UP7p1X/z6ru+7+N8/8bPJru358dDE/kf/C+OsKjaAyvqt1dEbPf+zvHf6VpzRWxjofqDPn2lxrrtIuCigPALvIgvmU92BeLosCyaqmcTUisH1lMn/G3VT9ypAAeMivtyrtEJExNl04WX3f9P/7i082bi/Ph1tvf651oIo/+92lZ5ceb9w1LgLjZuGLC+ozkBad9WPgop183Q+ahygf1kIQEFhkMWYOKzF+IJ8gBpnvjRhkrEHQYWHB+4H7P0XdlHjHUwdibFgMEGR2gZyuwAKkIJdZN2os3iDXbFtFSrB+OPva2hfSrcXj9853pw/IVVu+JMxfZM5C0W+JBoxkIZj615Wf7mi85ua624pH2tffsRBOy5w0j5u3Gcm/LsJwVsTGMcmcgL6UG7do8xq/FndiwzbW2H5JEW9gQdZ7/4q44N3rriu76FDLJW8Z9+Kf2+slGnf2nG8oSTEQx4jysR5jUmMdxZxMP78YIfyS9f8W/5F1EWse1oIoAmz3AxdVx9Lc8FTiapPpmmJArKhXI6svSVKMFcY4bYulIwQ7cxfvhRhwX8TDIREW0yIhAsYxwL3IAEcgbxECTuedrBVypa60FRLxbX7C76meYevPlxPpBW6fNriYfFgTDsviIY+VRa4UtUVa1AuVsC0SY0TEwurJg9OxXDZ1Va45WXzslqlZI439g7KweNNTn9xHfI3nrrvr2JhIiqg+X83NHx2f0OdSY6nyEZEyP6LzO7AK6awVXTzeGFNnfmNT4eNV/2EjXnokROpNiRR5j+p+eGiqXvRLIfJmXjmcK7hTIuNHLjIQeAcgZ/ro5bg7fDn5Zb9nEsgkkEkgk8C3gAQywuJboJGyImYSyCSQSWATJcDCH6CiLoDnFoFGMnhPATifdoWZMZEWdbmFKmpDVnBB/n6dRzOZjbyZnQNemoskA+QpHhsJQA4IDYAMQCw2VICMPJO4CLxzAErYKPPdCBAD88nHwHsDUQHeDNw0ywc7Z7EejuuanjZjv6w9gKB/jntNA800dPkb8317LmUhTysb4Kj9xnfqxj0ARdQPX/gctllFO9yCIxrJwu9GmFhZNqqL7dGQExsz7kHWbIiP9p+Dqyaz5uA35A9whPy4h02paetbfoMWHzzXCBey3C+Vu4+4aHnazf6LYbf6+cdcuDir84CNAFb4cydgrbm22hTXQBdxC7KhVme/3q/kD+RL+9MWtD3AOwQFLm4YMwC1tBnxWwAEaa/fvW/xc8f/j59+bexWHsl7Gm2dcn7IraXvTGv+3wpcMuGNes+eGZ/YFS75biJdnZy7ftx1o5wbbcuLV5y6dr7ghrqt7uSZ5UKxFnVr3Vbs5oTOrcX8/qigkmNe1NOcfKeeNyuN8UcE7pZPFWfcw6N3knIf3P2TLvTytWrcIHTmBTIWuVEQkblVFhfvwwf8QmH8l37+5//Zk//s+f9gGvCXAti+XLsxthlHjEfcW71XCQ3VjQ7GJMe/UAIYJRbOwwIHm9LcZ7zb+DbwlU9k/6aXKwS/qzKfUgYT5aTzSCXp0JYH5Tbmy9uLh39I1hXVkdySmxDAfKq70w0Hyy4XhHrgBSIAdJ5VQlvbF+jZuBhpsRhObummhZ2NeHhKgYABZDsCrQFTvdVo5FQSdE+2Um+5lJeireeq8hUimfvLCqiNqyeFrvAPh91om0JYTMrKYk7lPqyBvbrcCFdFaCx12926rDBao0OlSyYrBmQEufAPlIjR4T6wzfuZj84n/yNMw2231h78pKxAUmmmV/dXHts3lptPSkGTtvslJeS9/oDE4ACMAsA7VnSd9z1Q+4t33uieWPvo/Pflkm6uJjueKfXPd354+h3bnqndcLASNxaubzy/W6QC8jTyFU3gn1FijOEq7D5ijei+XsyR6c4Zd8/Sl9zx0g43Ltfpexov1NR33Wh3yd1UP5hTH9+m9oI8ZA4HSJ/W355IC/eOMx9xz1RvcHId5c4Wpjrj4cLMzatP1JTPIRF8NY2FFZWFORjihPuRUS/GwMAn/Y+A9r1O0beu4Hm36jnXC2w/KKKGPny/3Dvl5Z7oyB1Dn33v1sKJ79M5rjvf7+lXuv7f3j70ecVRKbmthePu6eatbimamhAYv6QHnSn5jRn1m9fI7dELCiI9f7kkb798jD2Ihr1K1ylf3FTVIO/0knhmmxceua67Gr2x54reeT/zw3f36qt7zR0V7cs74atKkFSQW1hoYmn0aSWI0iux9OF5yJB3VUGEwh0ie16j8Tij7+FM4Vh1unDitZP507MQibKY6DWFZDaj686/a7WmkSq7Gjup9IgKuZLS95ITMejdUHlsSHEt7pYl292yUHqH6g3x8tdKxBehfel3nU2wtjBLUpQcmPvHRFZA+Kz+zWJ6SonYLhdMJFfiNqsnsEs8+kTF4HqINQ19gbY0RQ0+zT3lJeb8rX0ZmvuqgcWI4jtrVxEMWiQveCIXfDe93ytVht3xymh6naYdiHDWj1zLGpl5jrUAebBeXBOQ/zG5WZoOCtHd1dFWfvHY15qaV67cRLlTz0zL4qHttuxZcCIO3OLxUSdXS3olX5J1xcsJnX7MuhjSohN3g5nWWkkOIFuy0vOcXDc19Mwzii9RnXt+akpkCmv3YZEUjGPq0VPOEYFym6wvviB3Vsc7zcJ8p1H4vMpYUwyLWzT0mBf7R6p5Mi2LgJkSceEpXsa8SIxdQaEtl1pFl4ioEREiYsb7anO5fEYkx1a5vyqK0BkXUTJfGU2Gb3tH99RDf1T4VNj21r+7/40e8nkl5peMsHi5ls9+zySQSSCTwKtMAhlh8Spr0Kw6mQQyCWQSeBkJsCEBcNiijT1gG++Bc5qT1f2xax2WNlah5ao3m+UBn5jAs7G1eAwGgAMAmfWCWRmwUQKEMcuHw/pOjAwzXzfrCe41104Grpt7pUGg36wpjEAwQoBP22wbuAWhgIacESJ8musq2wWaxQTl43csQbhnfXDfQTCBa/9IiXgC5Mc9aP2yqQPEYeMG0G8WDQbC2zOtDhvVRbf1wC4AQMqGXNj0ouUKYQDYzSYNYBCNX4AQI1R6wTx1WF3YnNIeJo/B5/IMtCexmgCkudf5pRXXeq6tAOs3u9O/bcGcaSf6BXn9pBLnITA+3n/WNfuxToOWdgDwMW3U/0nfiQMAcEF/wD8zbYblAN9vVkDgtzQLlRe+sOd1J3YuH+tMRou3pb7/P3e25t9SLEduYWTYhaO56YNTu6J6XMoN55ru6cqGOH5hR/esm+4uF65rngpblXy7drZVGInqM8FacqMXpTHwU9L2XMsvl1eDoeZnJ+6r/M3kW5y0ySErem0ot09uqjsf1xW1YaNGFdHxXgUpztVz1T98vrr3sb2N57EQQYv6oqTFJXYO+vUDyETp25UuRlaszw4g6Q+UfirnhV9+oXXjmT3lg4xByD3kDDgOWfG1SNobF+jQWFz/a7mDGpFVxXLbK3xyd/eMgvYkWwpp+LmDyYG/kIb23Fo0eoPc8xwczi19QD7ztzWTqkBSONIXHb+vM2hrv0+JmBb4xz8P2ALA3lJ9ePRY5+xdK42xEfnTX379yF+PKt/yye7OI3JhI0OZ/LFj3V1hGBTC6XansVUeN5I0ibthvFgp5aO851Uk9QVZWHhRFK0mib/cjZMjJ6MkPJ3m84fScmUoDlor6lBvXZy/7PaRtnfrc4dX/1slOEdYjOfdrd811f3SxxZaWFTcdlvti/uOtq8fFvj7Xmmza6LrAfmDZAXuUda3I+3BsdPzk88wO+4oH3ri7cGfHD0T7xgZ7ayUDnq3QKpVZV1x30Jh8tjexgtv1/XM6393Azn3yApcmy3lR92Do3e7lfyIU990IjucLCmc3JphReT2NF9wchclf3Yxcyr5mTVdb06GHNjdPOKere5zy8orl4bF4yWRUuHq/udq1/9DxY8duWdZqvFpF8IRcJJ3BPMmcyEa+fY+YjzEAoNXFQQ8OnjqT7zPT70uvyLXVLJejEV8uZnise3qRyWRFTun8yduHcstKEDQxkrslEsAvUIwR+768hNO/SOud4ZHx/NnR3Xek0uk7ygFjdFmPPQpkRoPHj73Tr6cg/pDevP+WvRlXaRmGRH9s0Pf47KXNm5L61N35BphtYAnsjT61Y8ejO44sC2RpQDveOr7mBJjjvHLuwZ3icyFkHZ28C68bOKsT1aMyJpnr/rZ/UWvc7MAzdywv6xA26dGVf+CyBs3nFteE4kx1CcPbb1gLvBkqBY62VfIIipyy+FELwYN5AWWU5CQIg0hMop6ztuUB9rxWPT8uhJz9Wc0hleukLRAvsynjA36DPMT5DHtxDsdYptPyBGeBRG8ace6+EiWryl88Mn6wGIbseZh7cd6AhmaW8nLicmzaWX/JmZkayoIRMil3kH8CvW9k7tvj9PhqdTPFdMbNHEwdkx5BwCdcYALUNZNkYD/NpYUa2erb4m6mszbueWlkyMdAfzlwbcmpIGCUjsF43bdVqFnfSGCA0sLHs16zuaXQbHwDMp4KQcZMS6pzxk9v7t0fHRFJEG7otgZCpBdV4Dv4sKR8UDl5N3JOpPxyj2QxFg/MMf7Klv51NNb3qC671aplkWoLCumRVs9Zos61HN+Pr4+V4gJxu3k5sq1G4XnFdn7WKHavWt4qu5W52q9OubysfNz8V21icZfq/6+ro819niuiA2neBnpl2XJsryME70L32DM3cw7CbFG5Bbqst9vlyKw7JpMApkEMglkEnhlSiAjLF6Z7ZKVKpNAJoFMAldLAmh7suDHqgL0DaAJ1xWCdfalbuTuwOUmC660h80RGzkLuAlwzUaNzaxZLPAJIMRGmBgSbNAPKgGsWxBCQEY2WWzcDTRn08wGnrxtY2bgOiA8eXKNmYCbG6pBIoMS8ztgEtcCEgOeUB82QbapGXTJxD1WdkBTNuxomQK0AK6ZiyIjAKizlZk6gDIZSMcmH/m9p3+fxeXgGQYQGHEBeEl9yd/kb9fxaddRNmTC/e9XghgBfGXDRntgsUI9QZyRCXmxkeM+2sVihZgbIs6bVYr5XaYdOD/vpt971J390E61O5BQ20WrtC/1AJACfKSPfEzpZYM6Uolr6DDgh3ED4ITW/4/06884QF5s+jkA0P+DgNNtCnT9j5+v7O0eKe7+lJ9Pc2nXe3dcC2bmhsedP5q6p4Z2uaOFLWapo45tcelfLNkThUm3LBdPAg3ylZs6+Xh/3o10W8N+PW17K27JC9M1b94VFuqT3T8bf9fjXyrfc8+fbXmXQ7N88Dgrd1DvOv3nrisQ+KNb8IRx4SEg+fsfGr279l1nPvJpERz/XRrrh6mzNMovG4zs50z/erPSjylhMWFj+1K7j/p8+hPyTz93NpzxZkvP7hZwiYwZnz+htJHG/2DedQGz/0UWFVu2hwsrIipOiLR4Qm0zVky6o2O5tYN/4HY2RYb87lo8estyNN5ZjcbW5ErmHYth98Hx3Nl/rlgEG5UVSxEIKwJL5wR4zgF4otEuoHnLfDi9X4N8+1I0OY27GlkrFAVgn5a29yefaN+5s5OWFuT2BsCw87H37E3f+NsPMlcsKi5F1Iu0HbphwcW+/KoH3SipKCg3gVG6a15+6FiSG2opRsmKK7TO+EX3fKlKH7xsTdQPz6eNd015nyz5PTLJ/eB04a4n1o79slwY3SPA/TU7iofuVt19gb/MOcz1g8clgUhRybvZ29G8efXw0JprBa+fjk67idZSj2R4vrLnHlk49IiHdVYs55+jdnIKFO++PHKH++LYPU6un4jL4tQvQxEUqYiGwnasK9YOisToYcFGgjOnn+9rspxwioHhrmsecqW4JUGP9yw0mkHVlzuoqXZQ9gnOLoLkLpWFdxL1xbKOTP+1Em6vmJuNuAn+8Qv/94O/uev9+eMj224d86vf5ueiFYF9+7fkTt1UKdUPFLy2y/udHiFxsfpZRQUIikZcdfcOfzx4eO0NKofv1BdnZZkzKyuDYXWFZbVJeMsnfvOLf/7m91+OCx/eh7z7btAkVlB4X2DSg3lZWVZdvLLLdTs35rrXDwey4/EUwkXkZ7cbtQ+fWFr7zak4lKuxSH0aoB3zC97HgLZYJkE80m+QB8SOudO6pH5BvftkBeN4uwJr18Zz8w2N7XkRFWk7Lu8XgRHIauK4AqvvkCsoFQ/66oLszxMWnB8OlpzCJLuJ3FlX6IgEEnmRaEmzGo3qe9yLSzPqLYjciHiXYyXJwKYuP6v0UY1h8ksuZjG1jsC29QvvZkBi5gPWIcia9/YLSky+s0ooN0AUGMmzKRYNL0FWsH6wtRsvFRRIWDuggf+n/XIxL5v1EM1xLR20GaA9ID1t1jsCnb3unmhh5qa4KLKiqinjo+o+KHMQH4p+gpIJ8wJpVTEfHo1D/165etpVrHVnZW2wKIuFJ2Sl8JFuMy+SyDufN/lDUsgxk9I5BQKOlwm2/XJkhRGrjD3GJu9FyFXadlkWFX++drZ2dnhLfUzBsve014qN5dPDiyIPUGIy5RdimdnaBXKNfvNjIhdOMqQ0L5VzxciT1ciRka2rx0tDbU8xLT4gQrqE1YisKpqVkVZ7dPvKfsWqaBC3o7FUdkndn/eKEX2uKrdTHeWxKBdYWKIiO9bfxTjynpnYlRxbm/PlKuu8SOwL6ytiquHCbVMsfl/0hOxEJoFMApkEMgm8IiWQERavyGbJCpVJIJNAJoHNl4DiVrBxZjODGTuANDslgEc+z7rynhnXXV5zpb1sdtgcmdsmwHI23mZZYSQDILkF5QW84by5VwKghwRgIwTIwxaEPM3F0nqtbn4HeGEjyEbe3CdZPAZ75iBCwfW4S0LLjbzRlIS0+KwSAAR5DPr5tbpSP+QAgHVYCeICEIZ8jKyg3FzDpu93ldicQm4ATFA+ykldyNNIEAMtdOqCw1xKDfrI5tpBsobnIks03CgX8uFv3KAQRJjzyJjyWD6mPUxeZq1CWQBDjGSgruSDmw42h7gv4Jq88/Jy0r8/crmRoqvcUHOrD9HOFiScMtBH2FQ+Qt9RHAvkca0fpkELwPFTSsRfMLdFyGaQZaB9Py5t9EhA6z3yPT+u7/HThX3f//jE/uZduUe3LRaH/Ie27HdLATzSSx8C2F0labsjhWmnQNGu7pfd2dyIm5OGeFdWE2+qP1qczK0U5QBneEu04pJJ78HPt+8r/2nu3fse9M556ZHP/xc9ZDRadpOds3KU47mPTb2t9/twtCpAt+FOlmbcpybe+J0nSju+88b60/vbfulXFd/iIYFjnSsgLejjFIA+ZaTb+vKgeYy1CnPGLyhBblxwqAGmqsHqPvmnn35t7fO7il78nbrgASUbhxsJ8ld1Eg3qe0RMfOnm9pGZXd25RjVp43N7UnV/IRAiJcuLzsLCO9svFCpnWy53TMBmcKxz3RcFNM9NeadiAaY/Ixc0/0T5DLa5Pe/n9IU54oPSfo/2fvirKyc6+OX2bhUZEQjwPy1w9Da5mpKWeLgitzaL0vpejF2uLfAZ65WW3ML05jfc8PycSAtZWEij1XXk2PyM73kF9aQz+j7kO28lLJXW5GejNJfmbpjzCqpC2l728yNyDob7nkXLayNhrD8HsfIrJ1bzqt9v/MhMHlkysW3dV1l8myxL3rwQbZmUSx6FWhE14qSqfo44PS8D4eu+FGzPA8YXeyZAslwkua3+iaE4rriZ7mk33l10nxp5oOey7LbVR52CZmMZsWEWkBP0yeeq1/fIipFwxd279AWneCs9ABsCAjdnM52Tlsd5AlAZMl+fP3AF9dqVR3qw92/s+jEnqwi3KuKkGjf9ueKULJEKqm/XV35GTjNImRf/mdKblF6vBCB4WGmbxsUL7577k7Xl8dro8WDmziPNvdGz1Ru806UdN233DyuYRdcphonL+fbKvHjL9MB4CZXrkTsuyTR3yD3UhHwlte+Xm6hFWW+MzhSOviBg/cylWAP03UHxPp3UGJJFUSon83F3zIsrxTSpjLqocbvXaW/LpbJw8PdqOqirDEkcxY2VeudUXvFSfv8zL7Tec/8oRBzvXt6ZHLxjAEuRD32CuBj0D9wsXQ64yNy6R2Nuv6xQlhQYe0bxY27SuNmu+C/5MCk6xfGYGvPOKl5FSFD19QJEgeD8RIpVheYJd7Kz2y2GUz3XUCIf5TUvwOpFL9jYFUUgiRwx4gPXVhw/3a8PdSC2RbyetNiArEAGzD/0N4gtQG1kfUgJkJX1EG64DKBlvON2Efnwbt5sssCUOwCraRNAaRQgAM0pI8/GhSExeJhreW9BYFislnOSuDYOOhLrHsY083fvUMwKge3+jtUz/pGxHXFNMS2Q6WEl3v3IjHU040AvTwehcSJf+v/Zew8ou677vHefcnuZXjAFwKCzgFVsYgNFSZSpridZ0YtkWUnsOC8vy7GdvNix/bKW7Wfr2Xl2ilu8rEi2oxbZjmRZxZYoSixiEQUSJEiCqAMMML3f3s553+/ObOjOECBIWXFE6Z619tw7556zz97/Xc7e3/cvdcUZcqdFBgwpxgOxK/JypTQml0obyAr7jJcgKBgLr+SgP0EwcNg1L6Qiln/vV2KdupibT99/9KEd/SrX1er0qyZwxvUZqPysoyHMCdRCWVlzsgZlPNFP7Po0o+DdE7tfe6osYkKxYJxifr50SPPEFtW7JAuLoHtkmXHQIyLkrKw3FAPJdCc7iwEBxhXb4ohsKyb0fL3oHMYw5fJ1zbbRq+q7/Wh45Nyz3mP1qkMcqtYDa1/ic7EefiVzyiuRYfvatgTaEmhLoC2B70MJtAmL78NGaRepLYG2BNoS+J8kATZXb1eym2lQIcDDNZJh9amq6X2TbxrFmHZrABBs4tgcbFfiXjYwXGvBdjbDbOKsBQGAAVrnXIcWLkAPILe1yrCbcggCAH9rdcDmj3ysdYHdbFsC4EJkBSKypIfVMEXLEzDNbmhsAGSutZYSFrSylg7NIIlKfJIPZbXPBVxAK5JPrrcBu20AYAteW7lYsqbVuoNrAC6oE3lY11mUyZaLT57NfdvXn4NM2ESSN/dCmCA3Dn6zmrL8b8kdvvM82o38rBY89YN8gIRB7mhgD8g+v27c1IgJa2XTcVO3CAvqSh3oE9xLudm4kucT68/+Yf5ADrQ9CXAD/+2bgWvaBqDgUwIYiwJeb9HG/B8KaB1GijHpCh8yVzkf73x3/VhHv9sfLphluWa61CH3RUZWAU2CArLCHrLIOP/9/vTVRhYDajjX3Fw4YqYTwzd83n2z+VbNhhTY+JSrVp/+dldtKTVSmsgqdsDQDcvfkqZ71hzOXCHgVqFNlOzxh9t/yty4/NgHu6tLEIP/H/3hlZAW62Ap8wXywWc8fsAvdNy/3vcAYLCYeJcSGu3ntUslz5tWG909w+b0E9KYfpv+T15EY515gLHzh0oAc4DN3+yrr5zdXp3OxYOacJIwrWbZXgviUwL6z87Wd9bf21lzjpWjFfncXlbw0ZWzxb1l+b9/bry8O3t1+vHD12ceyuk+yCpc4mw+PqTynJE2vNw4VYsiKHBvc81w7HQi4tQT1TBWkzC5bO0AACAASURBVJb8uWoYd2XBMScLEedUec+EtL4LmwkGkRaMwaqIC8avnWuYVxcaGrRG0bVfiHSXZ/zoQsHxegLHcVUHxizzaEMyJzj5y9W+jyoQcedfz6+uvLEnOzkQjQwl3Ub3Xd0d73lkOWL0W9PNDiCwDvo/gOf5Q35DJva8cPa+cjxyw7mRvt21iFTb5WJILMqL9hnkM9J/3DzTcb2ZKl5p+otzpiLXKMtBp1mMdF/cukK/4MZsNjZw8mDndROnkmPJPfmj2xciPeUDC/dHRLDNddaWFenF9IuUYu7kAFRHg5exSl9otYRrkgD91dkm0TEb7ZNLqcWmtcfz6cvN7vRxxcF4LpWqF0v0k5bqAgxacJDxf6s8nJh61LtrIdVlzkZHzFKjK+wzs/LnlXWnayNuX3TKdMYWjCyDms9cP6z1G2XE9RQy5R2Jm8EDXNOUVfyUrCt6TMFRSHZZBoisAHx/e5c/d6fiOCwqnsWf6FLAxksd9KEO+rssKiTJxtEdpnw8HYZXD5nqxBavsdgfDaIx1x1RTJR0rdHw5IKMfCdL5Vq32LMX0snYTAtpwTzHu4b3EvKm/CgMUB8Ic6wtqcvLtcbi3T2kcbNXLp/Oapz0ykpiO+6bqiIrRBRKfgWVr8y4tXW1FjT8TzsD0PK+nsQyRpYYNZEeY7PVLSnJDXdsuj7c3Qh93ErpJemZnfEjsnzZYPUCcfGAEsTpXylB5F/KUoT+AdjNpMknkzoEwF+u1x/Z8N5Fnigf0H+wxLDvaea7lztWbd0v9kk/t/GVUHAgX5QdsAYFzIbgRW6sj2hD3D3STtST+eWH5liPX2GJpg2uBKXxL8LCeaBaNHnPN9s1xCHPAc1ZIyJf1mCkqKYmX0D8bgWvfkBkxT0iKeKzx/tG1WneK7JCrJ+stS7Vg14s9dZ176UIDDsftebC+nq7kl2jvE/f366yiEQI+2Tp0O95wSm5h/qWYlPEdZ55nXXmZnKF9SDjnHdoSaRMUq6dpPASKoS881Xls0/kxX6dH5A1SVX/e57fYEBNdsdr4yI4jsmiIivrCxRpFhTse0DuoSZUBvogeWPZomlHLMe24P5Mb/DJ0orHurN1rob4Y0wl1GarbbdQPzRDtF3RtgTaEmhLoAlMtI+2BNoSaEugLYEfAglIQz4nTXkQToBptKYACNjUBCbS1WW6bouaem5R7oG4hs0BBASfVvN/e/PaNYCf90czQOX6OUs2PM+mQolNIAA5Gy1rNWFJA36zfnrte8haLdASFoBv3aTZ763bPquqSh5stMgDQJRr2EgC/lBW6wrEWmvwDEtKcB2berQc2TxxPfexced6NvWAq5yjXlzPvQAU/G/JG85TbmuF0lpeAAT7f+v31rrwXJ5n5UGZKQPtw4YTUAiwAzlzWJ/sm61e+A0ZIAv7TNoIsAT/67jostYb0ouOKV+vZLK3Cmj5A4HCTT/lNrA38qWv9NN31p/7w/yBTAGeaBsb1JIg263WQoDxS4qHcHZ3/dhCKsiPzru9w6f9bU1AYcYdJFqwebp+TbQnOCet67qJhnVFvf2OWwgr4Ii0zGsKLpxtFCoD9eVYTq5wli9hiTEeHWxqELvCHs4GO5Uv3eQ7x3b3dE7ajUsdwcrH5hL9JbnCuTzeqOTkQicv7fbOD5356D2PdN287aNbP7Thvm923yJ//3vMDbVvQXhCDBJr4JBIi5IsLS6sDr+xp1BB+hV9Gd9TBNrefGAZRQLopL/Sf9H4pE9yPbJvsjsCaXeJBBiRcmgcDfmLEBb4pQfExM0FgAdp8dbCs3UF2GZu6hfhUQlDd6Xs9GZWw7G5b7s/nVTQaveeWCMolGszTxbctED3hN/oKpyQR4vFWv85xXP4S4GqgC//ZF0Wth6TKstQLYj+24nKzoo04J+VRryIitpeaYbHi0FSIdKTAjGd+kx1eLBJACjSyKnS3iZZIWLiAiJpnrKEBfMFsjivol9yPPkBN9MKIrxaN4511QS5wz1xLC302XSwcbGgvjf87Ve8mepkn3z7XysXVXu/PO/f956B/f97dyQWubnjMnO69IAAcvXVTa6M0vnSw7KqyAms93YdO/v47qNnt0Srtb3leNSbGpKsejL+XL802oVE5bLf8fyF5UCQbshSoGjGw50ml0qawdU5BWaNm+ezlxmIs4TcNKlNkTFgKtq4qwvRnsnPDL27KCuh/EBl9nDeS/eKwHjLTKx/ZTI+9KTIinrRS9RHSueKup76Mz8zZxIzAEKavsdYBVDmfbFdKdtVXfrWlauHrxQBctMVuWe904mtjW/03ll5ovM1fk91Pr+tcca5mMUHcoWsKMbippBMmCM9e81yosOkk4tO2Fv3xxpHhPZvD+uyCSD2go1dEavUXoiXKl+uRiPZciKaUR8DIAcMZb7HzRIEwIhk9S/kGmpXRuA6VhaMbdphNHZKeQWdK3VxSv7sN2UFcPjnT3z0vOaxbesWSwD7vuuUXMd8E0QypjFadbwOWRmle6JBI+uZjqAWDMh+JtBbINmoB91hGC7E41EBmaEARbdRVuCUVMKd/uLBc7V3jTf7IeMIiwI0+NHSB/jmHKQFxAHvomZ07FarBMq3yUqBiWqryuYrqPbcvuRTQ2crY8MQNVvjJ8y2eMGk/RXTFVmQtJv8hwVzmZMhBrAcRH7MHbQzpMBB5dcQ0XFZX3T6ivHyntdLXnqfhYuyeLoi4RXSM1UFa/fnDYTSpjmE8nxU6V8ofU3yPSkri/KmMlMO5NokWpRYJyATykCHtwAw7wrWVCiBUG6uxd0i15xWarrwWSd1XwRrv8Jg3KwvbKBvgOcxJSwr3qxEoHd72BcD1gL0N2SHzDaY/2hu/0E/WG+xxqOffoehV6sCoG+/rv6Zvh3BjU0rhO9YEDGHWEIU+fSrVaddBZCePtp/QMD/LgWWNiIt1NrNJRhGX6/0YO3NHGatjV+p60TuhWTgXd2qESG2L0z5MgAUyeCkukpX+7HapGJpPDhzvO+ArCLu1vrgQqVlLsXqYUZBtCcXznQ3sn25hu6/Xq6h8iI+RGCYLpEfp5su9JzmWnrA84MhBfomv4YIjYKencS6QtfYNTRjhHmjoHvGi0vOKclyRN83xPzQ7ygHQBgxXr6h1LayeKU9qn19WwJtCbQl8CqVQJuweJU2XLvYbQm0JdCWwHcpAQiFe5UAvgEX2NznTc+bssbrqJjikZpxOgEAAL1IAA9s6LjOEhxsNtgQsTHmk03u+HqebHrZ2DRNvZVsXAhADMBv8rEukixIbzf3bGzsZsmC7XxaIsCSBfYaS3pY8N5aOlBOngHoycaJ8635WpCfTQ9EANeh7WhdZHEtmoiUC7CFstu6WgsTSwgARtj4HPra1OK1ZW8lXuwzucZq1lqyg3M8m/Pcz/P5ZANtZUJbUUbOW8sVymhlYrVYuZ7fLUCFzC2BhCZb0y+3EgSN4sJ2PmXiw7eYquKvmoC6WTcAyIS22q70RQr4v/oQeLa5CFZ+rcTWS10jXPCCm/EXVe0iwBSAO5tmfICzybbkD/fT7wHGH5SrkYX35T516F2NP+89GR1bcVec8KODP1Z7xrn6PCtRDNJGWr+mNz4ntzPs1TfWTRYA49rTP1yTpVNvfbWjt76yX4XvHvQWZycifVNlN3p9wY1DtG04CHwpLX7zlcgtpuL1mK8UX7/h935nNnO5d8SR9vItT/nXPL7SyH4qXcqf6G/MFgXcVgTQ/hfFA/ig/Pv/pHz5b3Ch85Gt/8hsK502w6VzGT+s/5oy/i2lgyItZl+GeyjbHwGQD1ygL+FaBxcyjygBsgeA+GqHKWn1z8qdFpZb54EXAhfLt38cdzmjAjTXNf9bs2WeA9jA7/W4EmB+E4zrry/bMSSrI2c0kDRqXv/Maf/HyzVzRUet1ui7O1mtF2KhwFGnc7rSSPU59VMLQSZSqva4s9WhGZERuHlh7qDh7l7zpu8MifyQ4/+uiNwe/XSu3vHHIivSOp8tN5Lp6erookBmX5rx+0djJxak+T0uoSy0uIG6gFjOn2qCPiI1NmirP/Cj2yvrpIR1cWctLCDILHHJ3NEkctdB0Wam9rnHi1ekFUz8JvWdG1YbHdc/kQvTHxyKnSfhbum8xRwvPNWUcbRaP97w3IFksXxi/6ETJ7Orxa2Ram1fz/zqG/SbCVzHpHMlk8qXzGpH2oyenjVeIzArnSnz+M1g2msBr+NyLbUtftzM1QabbnrSA3PmaP26Jz8XfWtJ7sj+x73TX3xMBATgVKnkJaKPdN3i/sXQu4hdcdNctG9rLKwMK75Ktx/UJw5nrzz7dPaqr46Uzy79+JmP1eWaiTmOOdu2M7JjvmtlBemPCcWy6Fesi3Sqkd/zaNdNoYLTx5X/qaVI987p2GA4VD53Mt0oVPsqc1tUbsZ9KwM4pTG5pRKNmrPdW0RceLUzHcOR+f4Os6wY6Qm5VCPIczxSVLDsXDNgOzLcdexcbfjs3LCIneu7Flefnxns/sTzV2x/ROfCYjLu5DKJcj6TBPTepWf2ith6y1j86LW4NlJwdiNAv+nqSFY/BJB+p6Y0LAbe8+GdH3phs+uiTcRFRHreAgtNTK5cChEn9AfdekpuoS6rh950vVHNOtXaYK6uMCVqRsVJqUcibk6q4a6ib0e8iNsXhGE+4nsVz3MXH7nBrSoQN+8/CCEIIFwe8U7CygF5875B9vy+wXpg0/zatHwRmRPKBdbyTdmvK7h27gMiJnbWNJdVgkR9S+yMT0wKAr6vH3bOxzLlF5UmlJivmF9sHCze71HlMye8+XHFvJmUzLZqPC6IuCA2TURkRn0gejbW5c/fuMnKwj7nP+vLnyr9ikiLcWM+tCGmxXrcDd7/lIf5ie9/q8S7AlDbau1jQYEFA6QGawfiREEmICPmJcgMZGZjCdjnN4mdl0la8P7muYC7rF0AvX9CCesiDtYXlMG6LaRNIHRRZODz0r7Kzpfq1f9l3bqCPkO9rSXxvFqy19dMkeoJctn+YF855zylGBb7pTuAXK0VFGvi1gP3T74CSu9bPCsXjbIYI7D23+GgH9m18+aMeJdtfv7mR9kFhXXjycBhvTCgsZ2LpyuOYkzk4tmybCG8Idw1JbLlLyo4tywwnE/KGuJGES/EYWk91G+drYrHMVBYTOYisVpC14fphvMXya5SDHJQcxH9i3URY4G9A3Pus/Q7/cacNqZP5gpkzrqU9yjjgbGyJPdbJyslp0uzRut62ZYB2UP8MQe3CYu/Q+dq39qWQFsCbQm8miTQJixeTa3VLmtbAm0JtCXwd5cAIDgbIOseiPdA3GRuiJj60orpuWfIeFE2ExAaAAmA5GwQAO4BsQETt6//xjlLXnANGrHWNB3AC6CMTde4kg0+ycaJ39hwWAsFCyRZywg+2Uxz3m68KIslAKwUKHsrKUBZeJ4F29iE89y1On7Hv3UT/Fu/lnqyubdl4Fq+W5KDjRf/tz6LsvEs6gBAYAmGVtR58zlrgUHZLQnTuhGlfhx8In9LXFig12r02fraGBX8v5nosfeSj409wqaQOiN/Nrx89siDzEFTmdwr/c5us/VfdZgz/566UVfqbS1kWv3Arxfze/9xEUJi84NaSQrbJ6xMWz8tYWavaWqnrz+jKa+XS16sF8DKBIAJrVTa44zS3vXf79PnV1Nh4eF3FD4b/Nv8r+6vZryfGsye23E6M7bt+o6H/cWCXN7Il7q07Y206o1ASFOOHFcE5bzsISq1VKM8L4JiVaDiYaEfAr3C8ctKZ+a7G6v7BLLdL4uL+S3OoqdYC5GJaN8nZX1xs5xN3CoXUfvrjtdsI4Lz4r5HgLr5Un6jG2h8to9IU36f90J6yJm6/W3+F/7bFnd6tTsjg5Ct4WLq04WyXELlziZGPzVcnhx4Ib0HFyLnj89ueYd519T/aMYcUGDkA/qBcfE7Sg+LtJgRaXFBPdJ1kJwxhsY1oC8a2ZsPiApAR+aU82C6vlYy3vITqtcn5Dbpn9ubIGVEr5jDhevNIP7opVAvwATwkn4NefQXSgDeaF5zrgk0ysKM/tD0sS34XTYOyULoRPoafs+o48WrgQAYHfFKsRzLK9pAV8TrrdaCXoXs7ck4gQIamOeXj//jxeErfpmy0hfvV9vcjYsZtN85VWikaecBxaq4djR+8qjc95zMNzpuBqjflnzmmwrgPT8UPXMk6y+dlsuaV+QGhtgWrWDv+ndLdPIJMWGtpLCiIyYIc19B1/I7Y785n+l/vifqYfUaxdDYIQIlGTVBJuEs9D6Te9rsz6wZwWyNX2UmyykBx0UzMjG7okYuyLqid3Bq8QOdywLhG4rCUZeNhwhFb93Wxq83TDpfNg1f/VGqygMzvtl5/Jw5vH+Heebqnc34DIrFYPoEvjMmTpQuM4Vs7LIFb8vRrw6+btU3tcIVy8/lRFqUf2XvL8cUEL5vqDxZGE9uD0RU7NTgLUvutGVBn8FEYpT56ujv/8uf3SBP9Us7h23um5ZYnpyJDfgfHf3Q2ce6btqjAOy7+yszT4n3qyxHOjun41u+piDfM5CFqh/WHgByzKsQlwcacmw/l+02j267YUX1mHy26/IxWVPImibVHItqYwV9nlEfPWuufeqIqSX8aRE6g8lCOTI8MXtbsljZv/X0zMl9z5/5ajpfTDmBgNHQzLpBcO7o3tGjD99x1R/ICuMv5Arp9QLX3yTLAH3mjcivZj9TrBSjGA9XJvzSnfR3gerliwSJpnMCnivMr3lI7qCG94Sl5Pawuk1NF0uH1YGIaeRV6Jjq6UtYXiMMq42q0yHt6T5fDIWk3amm9MvVIBKElRfKlZrItq019SMICYhx+16kFxygPEo2rgnnLjQ/0A7MrQJondv1uf/ZwnXFy1NPNl1wiZypqN4xEayb3Wnx87uVuJ91B+sS2sUyGvZZTRB+4Pi7Voqp7s8VwvQd+ren7CQKCrpdlCyfvip4fFCWHMWeyMwB5pELHD+mc1jO0fYQIs0818kKwFfeAaxlWA+IBG3G0uI8cx7KH9ZNFuWkfLw/kBnjEFCYNQjvEsYt88oFC3GRoNoUhXmodf0AQcHYv1upldSmD7TGWMJ6BJKYddrLsZLjWT9IB/JnTNCeyApTvV5mFS+m0eubk8musFNRFgrquZ/X78wxJBQ5mFcsOcxc5CteQ04xHHorCmMv10jfCzlZctSuh2lj0qXICp7NuPumEoQF7zvIRM2YKqkX7IrE6oaA2JViZKJ/x0Kxe3Tp+m3XnD2zNNmRV2DuG2dP9F5fXEmuubFSQhGCg/8VJDy2dLZzQQG3OxW34vLlyY4n+nfOP925ZWVc+dOXURKirz+i+wYlkydllXF/NFHNyMqCsW6trykbY+qUEpaqyXhW3rOqDhZBX1HCErP1oK2YZ1yRTU7bLdT3oou182hLoC2BtgS+/yXQJiy+/9uoXcK2BNoS+AGRwMvUEGeLsEGj6hUCq5eSFpp8aEFakEubZCdvYsPyY3FF1viZgvF8qzHI5pxNE2AAZVoHFpqgF3nwv7Ww4B4ACjbqFrzgGjYwgIZoSFM3tP4A1dgksvmz5EHrppuNvy2flYUF8anfZksLzlmQnk0o91BmNkGWBLFgPb9ZSwwABTae/Gbfh3bjbzeJ9lk8A0CB/62ZPs/aEOjzAuXmPupriRBbH0v0WODMAix82rLYa1uJHL6zyUO2rQCQJUEs0WLlaTeHlAEtdu4FVEEDPW789AGTviplaisR4yaQMYCx3SgjF55Dn/n7ODZrElrZUCdrlWKtZ6w1CDKgvJaAsm1EXThPG/OdduY3zgGsCY9rRvY9r7Fux9kFrCsoB4QAFkfWNQT9HeCAvq0Ato0HdxePHbu39qWO9+c/Npwbin9goafjjogfyL910fW9glNYxQd9XVrC5SbQ+ODyPaa/tjR1WeLkwS5n8XGFLf7mdLw7LQIiFw1rh8eq06Wy4iwrHY2HtbCzka8u+FlntDYbSQel+Hh04DG5fPqYvm9V0O736Ld/TCMJiBPqWJam//mwD822a6jrvtb/pnm9d786cDU+6M78TNRU/1KQMvL9lJwuTWypz1W+vnJgIu+nvq5zGwgL8jiZ2iGXPY8rIHceggDyAbAO4JC5gj52oQOZA5yR309f4IK/pthKBNRctnEXBL5K7h8yX1j4B7n52kA15gwekUY+YF8TrOWQ2xj5t1c3dupPy1XOb+sUhBKAB+QFoA0AYROME1lh57BUw8QTcgc1KpKhp+QMZkph70Cp5nXUFcQ6EY8X9GmcUsPriZpaJRHJVqv1vYqYPp32zHwqnprJP/NvC+n9vz4uAPlv5F//9pnq0D1ogxMkGfmXBFj3R6bulkZ4VGTAIck4pwDb5YHoucWtsRMlkVTUdfUi4PJFxLh2+iLa1jYQMnVmXmUOZayj2Q3RjDY3YxmglDGBHBVjozYgX/5jAsQv6/emvMH4WQXOcN2Z6jGzL3y73A+tuRHv8HeZzHOHivsPHW9q3cZlxCDSwvg1EUUX8HfCOZJbXRteMV1fi/jfGpmYmzi5a/jOfCrRE3UqzYDSi7Ve9dVurA/iNd8vPDhwW+dXet6wrb80d2ywMlN7qPtWyr1jKdIFGX6DEu8SNHOZq5h/GZ90iNh6MOg1QVHudTL3AjJrAWjP1a7+0ytPy5Ljt2VTM+SGjZzcTl0lV0+3/PudPzd5f++Bp//Nsd/MXbvyJMQPz0qIwFisRv2HTmzd2v3UyBUHHui4NTbjDo3FEvl4KsyZLmdB9WmY3YnDCjK+aPrkaXFsfMokS+UMBE52pWAiNTnxCpsA3290LjUJwN9XIuAMbfXsnhcmnhg7OTVbSCfm/vytdz/Y6S30yLrnegWb7yJODVYboorMomJaZLzV35DmNOD4g0oXimfBvOmqV/dp3L5FT946q1GTDRreqKlMd8jyJ+K6KQUAmRdg2yWfUIJsySfsdQJnR02u18T2VgTe+qVKvRLx3QU5nkP2Ncar5A4oz3v/dUoA5pSBdwyu4x5Qwvpss1Y045Fy0cm2C9y8U0Tk1qV6b6hxPQgB2BuZifVFprAk2WxFBcGJQoJ9X/M+yNvg409OrDpHx+edTCrmTM3lTEbOce5ezBU/F0sdUo/sDUMvKgddg3It13vf4tuH9iSfOXVl+okHFFPm/76Ie7k/Vf7vUfqG5qUFud/ivcP8j699NMohSdEoZ66zCh6MPeRAP+UdSv2RGZ+3KEEqQHwD7vJ+AejlWgiEDeRO8530xQ3zuX2/88n4gAwmD/L/8HoZ9HHRA0CYNRLPY+6tX4xwfqlMXuW/8d5jLuHd1Hx3agxp+asFWETkq2dOxVLhvkTWJB3XOaO+f7he9ccVv2GP1B2Q9TWK1ZCq17zy0rnOpwXyj+jTVAosub7rA8KKhm4lJVi/2P5gFVgu9QDWelzbKXIYy51eWVOUI9FGWTEmZjsGVh1ZVSzG0pV619DKFi/aGNR1vd2jy2U/2uguriRKtaqfiGpJKCLG1EpR06hLlUJWIyRZkJSnjgz6Ii36sv351+v/EY3fkyrlovL5AjLV/92KjXFIhEVRLqd+VLLKeJGgSzEs6HO8n7crYbWyU0m6F45bWk3Xy/lQgYyCvgsE/cDFFSajkPAvJ2bPpWTU/r0tgbYE2hJoS+BVIIE2YfEqaKR2EdsSaEvg1S8BgaOtmuG2QhagtZpTnAdIsdfyv6t7rRb9ZkE0NzECWl+JgGwgWkArwLwlE+lImrnPEceiZKIjAGmAkGwO2DSxMaB8FpznWdaqwLoxgqTA7BtAh006gDj3sCFmo44pN2UF1ACgYQPGpsySM60umywADajcCr63uvOw5uIWpLf1t5s5G8AaoMQGyybQuLVOoN7UDWCAsm8+1vXKzltq2Hcl5y0xwqYLkMyWy+a9uS7kbevE9w1tu/5gKwf7advbEi+WnLBqe61kRSupQTlbCS/+t24FkDl+swEs6QOUH3D3uPF7fFOd1cax4ZnYtoypnEbzzYL9Nk7JBcT0yk5dhLCzbWZla+VL5ta1FZ+WxLKWP9SLBFCDvADLAGq5n7riOoD6U0/Ocw3ADG3Gd+rV1ObX0ZShLV8rQbhuHYAsyIPrAJX4pI9Zq5dn5MYm/ifHPzQ6HD13R24gfnUjk7x2KZmJZeuFoDdYbgyEc75iLhjFLjD52prBisBu82x1//Gt0fH/cX38saM136FMz2rnvvx8fGtdaYP7EQD33gOr4IjV8KuzxW+krzK7K+dmcm5iXC6ijguE+9tykHyLXJ184EjxaiNN7/XqrX1Im9+MpY6YlLy4dNdzIi0q1wh+sO5CAAL+8x3+Qw+9NfnXxU/U/gHzAFq/1Pf88bHRD5q75u83iiFg1v36M74+pJSWBjDjLd8KfK3Lj4JgqXWx4379ANkBwNmMtyBQEBmD/CSvyzy8eq6y/VknFfzYZ2b/yYY8BN7KNdStZnfy2dPD0dMjAokBRik7sqxbAJObfhod6bXxgZum7sCJR8pmoDAd3hSWgp3ZsunMyk8//Sce8dxy0ql3JZ1qw00mcmXP6UzUqytl42b0kI7kUE/jt4/9Qbi964Ez2+LH/uxMZdce1zTGZD2hdo0ZxbEwXdH5WHdkrvJM/jVRkRXT0hQ/LjdgB3fEjzBnUL7vtVYzY4Q2I2/6K0AQxATjGfky56FJzIFsMxBbQ/7EtZLHLqWdIlhc+uXicqJ8Kv5sfE9qLWD7WORNZvSp3072zC7h+krI95pFxQUOyBGrxQ2p8P8q8R54nVxDTfXPLJX3PXf60UPX7HqvZs7riR1wQ9NiYMTMyUWayDxPGvZ31Pzo4vHULk+Jcu5Wwgc/7yzeL8x/vIM4T595Qgl3I+f9BdlyvUxXOuaF9F7GM2BvbNXP3KA6os07JuLi+S/1/0igVPz5Yx9e/IVjH24Cxd+8ff/cTEfv4OnM6JVTta17y258zPWqW5quyfSqx3VTwq2J7UFAOQAAIABJREFUFY2YzELJDC7Pm2itZkRMqF2kyL1O6LTID21iCEAOAOwmSStSo6B7jr3nL+9bLNzd+cChyE0780H2HhFjHXI7ZqYqo0Zj3gxEJrviXhE3Skc0dnKtRNj6GKSvbVcCIPRqQmAXTDQxKPCwMxqcidarOxVgu0/OoPzABCXHbRY+K3f24u7CHicIUhLQEaGV3W7D2RGPxeeTseiUYlmU7r1umLwhhAFJMetiguN/1gHUifkYEhFyo8lgtcyrzC+jmoducZwglnLzkb3Jp8dEdXWVg4SRK6hmcGzIn5aDeZv2vlMJ4BOiAPKvaV3zkb854h187pwM0eT6Sr7kqK8IR/dar95Y8fKrjzZS3eoou9SDu9TXCyJDI7lcx6LmkvF/OPj7vym5/l8XIS0gy76yoOv1ybOoI2OLtqJfUhbGGP2f9Q3jkL5P+azlD7LgWsYmfZd7rRun7fpu31Mvcg21Xn/6H/fwTqSPMiZQzEDOmy0q1m/Z8PER/fdpJauIwHsz9zJc+l0or1f7OSYw1kTvbFZEkm3abMnEibeAXEIlYklTa9T9juXp9KiA91CxKQ5keguDjhvUy7n4aqKjZHLz6dXJZwc9WRfEq4pb8UrjVbje2nKzSQYYZ1l/GDetR6sbOmsB+1Ky5/3HWGTdLYIg/HymL18e2D1bU9mfUfnmNEcFya7icCRew4LKV93p0xE/Uu/MDqyu6PxZ1a1LlhiTIi9uzM+nI7rvkOociJzYrbL2UddaxW9ILgcll8tETnx1y57ZSd37euXXJddSDZE3b3TdYGhlJhOZeGbodOfQynM9o0uHYunqV0Vg0AfH6X/Kz9O10bPP7OyMpZZl5VJ4pF4pXhc2Q6ptOFpdZV3wBfRq75Tt8rcl0JZAWwJtCWyUQJuwaPeItgTaEmhL4HskgRZAtpWIIHcLsFsw2frN5TeuZRPLJhRNQ0BVqwlsrQrYTFjtRAta25U8LkyaO56XSVwQeNG6OWLjnzGpyyqm50eiJiJ9Yi+N1h8bCZ5HvpTJgsPWMsGiB2yq+Y3/AZLRMmTDjqYnm3HeMYDi1JfyQg5QtzW13U2WJOvn+LDa9Ba4tzEvuNcG1Waj3qpt1koE8FwAazQf2aC/TQk/zQAD5Dm2fi/loY52E7hZe83m2QqmW8uPNRXvtbq91GE1/lvzskSLJWXYJtu6WuLD9iHK3MpI2Xw2n6MMmwkP/qfv2HYDnCB/C+JDJvUYLylZifXquSdiyidKZvo0bQj4x730FfrM712ini/3583lt2SYBYEAKPlO36dP8b+NXQA4hJY1/0OkIT9AGwAi6ka9aB8AP0AcSDd8hXPQXoC5gJIAapZsIw/rE7k5plrGk5Un+VtXUPRFxiggKWXblgjKj75/9RMr27pOv7Ux5N6mAMMdx7uGE6sKkq3YE3L7FHF7zVzYH51yTsoVlD3kxz8Xd8v3L0VSL/xV9W3P7U88Sr4byEmBj+ev/48q2n84tPYv3/k8FmuChYzV6fHSrlOL9d5T0uI346XdLyIs7uj8kjmR6DdxkRX7zUn5AtqAiQF4Iav4r8f/3cknGtdHng/2ocm4gbCQSx6jYMRmT/6oDYxMMT6ohKYqGv3PiLiAtGhFGhgjAHTWn/v5OunLt5ToAzyLeA7BOllB+9B+A3IbNNfhLd37fPGaHvmaN9LAbr3fiJw5LmLAyKXLt5JOAbAGtzgXIgPsHCtFcr9WdzrURvsX5pwDsVI9Gi96vZ3y7R8tV+sCcdxlwUeRWq0+2BWUFyu+IhK7gp9dk6/U3cKj9bhX9SPJx1bv3vZM4TURkUFHpQ3u70wcGQVoPad4AxxyNfNmWTF8Zjg2fnAodvpgT2S2GnUrjK2Lue7ZULfv4h9r6cL8yDyLzG0QYv6HZFuQT/9Z9b3Fy/1DXbJyGKsG0cGOxEInAHFOsREakTC+VLtPl64RFvHoqEn4Q8Ly5kRWbBAt4weSgrmUHwjgC0BLm0MeAdry/6dFckwp9kWtFvFkodAMiHyPLAX+NUGkkRmWKbJWuVFyPJRQQO5T5d27BMYjK/oB+dF+jGHmEOoFGPzQ+jNXLRj+XcgMqxUsVOizNYGGzH8MVN41zJFNq5UP7/75SuebXgjV/zzFpvCeWLw9KkuKkhurh4UguVWWNJJdZ9OCaqviczAOFU/jsNzETYycm3Wyq4Vb3SCUrEJI1gupYdt3Cp+8o96nxJj6r3LUsvqB+z47e+K1l3/jG8nXbe1PTN4soN1Uwrh8N9WbnwlTYLL4Q6Xx9bawokBevA8hDanb16QrfbXvmO1yXDVZD8JGLTDViKNmUDh0Af1xBRAOA1c+00IBtoG4F90gd2gJz/OivufmYxE/E4l4mVyxwpzVWI83g8UDJBXPQmudOdMS+My5yLHVCov+CIFSlyumRsLNH9YY6c16y0O4DIMYwzoFq7QWAuE3dT1Wbbwb0BwH/F+BrJBVhTsxvRJdXC7FRVRkPJGMnhiYRhAGlZoir7hh6TXlhdyc75aOO/ETVeP2yz7oeT1ntBLEYuqDBZEWJ5PJ/J+rDbEa23wwR94hUvLpnYnnl+XGzK6RGHP0UcaWJcXtuo53UaubMvoYbcq8x5ihHzB3WqKCeZ13/nRrf9acaq0NWdvwLCw7bl+v/x36xPrjUsfp9efynuR9ifxWfggtKwwuhVR3ZMpaohnvQyfS0YSCJ2gWq5WdiWrROVhciUZKK53XNhrOfrl5issdUkJuk5YLS8lobjZdS/UUsSrwBMCHiusgq02RkU54Tp+sUy520Mb0nbisDUw0WVNA6ponV1LzQeBUFT/ipdrxkriN8uwTeXK5yjGqcnQkO8rvTHUXemVZMaHnxGKp6pzIgnnHC4d1DWsf+gHzaUYDrU9WEIdS3cXCFn92UvEtwsE9s8dEVPi6f0YExeLRh3aeU92HlfdtYd0NcguKYrEQXrs8lb1XY+x3hq+YGle+V0ieHfFU5QpZpCRSXcXK1JGBrauzGe/k49tOKxi3s/+e50/r/JTkWn3hoZ3Z4lJyuFJIXBHPuJ3xTPfTK9PjsmgpX9nCAPEeYby3rn0v1efbv7cl0JZAWwJtCbzKJXDJF9+rvH7t4rcl0JZAWwJ/nxLYTFSwGbAbVwA4C9YCgLJxJwFOAKICyHCezS0bKDbkAEGgiq0Av3VR1PSjrIPNT1Mref37perLs6xm4JomZOIKua+WS6CgGjOuZ0kHngkAxeaaclJ+Nt8Aj5SRjTaJzTrXAYQAIKHZBdiCxjabYggQnsP7xhI3lnRpJRmsawcLEq9Zf6wBAIAf1JH8AAXY7LUC39Yigrpb8B/5QJpwHeAyYANlpSxoe9qYGlxniQyubS2bJQ9snhZ8ob48k/9tuS0JYUmPVoKCfCzRYT8512o1Yl0YUYdWSw7+t4eVTavc7G+t5/hu+5QtI20FeIhVCRtUK1Np17knTPlUPxtv48m70Vr7Ih/kT18hr+/F0dR2Xc+IsWHlyXdAVUuSAOTYvkJZAMAYG4DagDXbW8pGfwAYo5ynlHgGICP9lyi/9F3Okz/jCr/OfJIf8qR/WbdZtAdgTlNT+1efKzn/z5EK4/O1Su9XAsSkfwMwkZ4VIPnUTcXHGm81f7X77I6+zkI2nj2eHPbnogxfY55M7XITQVUuoDz5jZoLe9358qKeWgyTChQTmT1UuX7vM3PXPIk//o/P/9MNZAX3v0wN8eAt9/9J6YXS/mlpzM/Ip/0nBfS+rRCkU4DBuI4ZS7wgAiMiRnHA1AXKbK9Pmy65rEcNuQUM/Ck98qd6nIVP/27iZz731uJfPK1yMo43HAURMevWFa3ncXHypnWZHhXAttAChNHOdi7YnB1txbxyUqkVCaeNAOX2CfA/II3WN+NuCdcwmwkLAbcdRwpXH5a7nMkrUgerv3Xj71zMcqFJ8gSubCWcgUTZ9DjzkbsVNmQg7RrNfSbWk0rEpFxuop7rpVzPqeRDNxBa2yskd34pcGrqZKnna5H9Jyu41mGOdvcKaFd/cUpL9Z6pU+U9oyOx8SZonW9kFRw5Z+SPf1BlD9P+qrIO6GvMsa8odsVmoV3o/5a+gosexizALvIdU3uh8T0lV17TfdW5kuc2tvUmJzuv8A9uGWqcLU+akWwg8CwmN00NlRl3TeVgxsxO/1Gjf/AnPTk+N/N3/pJJfRIMfYN4GT+4MuI9Qaf/mpKde5jzAZkog2XHwlsffCb/9DW7sMjrlDyOqv/tKUhWyAxwWnELLhfMfJdA7Nv0+9dFajC+KT/zBPM4pBRzGGObOYFnfy/kSX7IDPCO/shcwjxJvQ5K874m92Q1kWbpY6UrxlSuNw74Z39S/W94vjZYTik+dcIrNGPI6H9keUjWN0eLXZFPH98z/OzYqUlrpcWc8kdKWIhc6qDeb1U61VHIvfCPDv63yeeuu2ph2e+ZifhVyLxm7BSCeysodVQWHj8leY6L9DtrLQ50L/Macyjz1zZV6uloGExHw0aPF9TyddNIJMOwVm+EC6IJuqX+oAZ2y8qnqHkp7ctHFjisXELFBFsuigCoVSp1ZWFEWrguRMG1o1nmLt7LvGux2oKIgLVjLiUx35bUL60VjAXqX6PnDIpA64i4tQ6RBnvOVHYqLse42a4YP1iFtcxPgPxfVGLORykCa0HWSA1ZenizC/lYvR50iJnorgf1ThEs3WJbpCEvRiYwYUzBwrOuSRwIV4LOsH7okEndUDLurYoUDGnxDVlO3PS5ufdnzma3f+Te7v/+gmT5i5sah773V0q/Jbl/QfPNsxr7Vra8V6kbZdu+LgfmNbtOa80KWVFuNOnpx/Rd+jj9jTFjlTGa92guZf6k7yBDfmcNw7uNxHoMhYKXOpj36G+UBZlBTLOeqv0wkhXrgrLrpUf0/y80z+mMgrmYiHpmoiN8JJ7xnKkjPenCUldWcR+SUukYUbwGvakVRscLRhSPoVpejelPJCfXSYs6B/HQqJX9Mwo/3UpYMP9tgYQTkSCXayHtG8oyQcttYmU0QgXBXpa7pnG5X/JLq7LQq7QuDS/atBCEKBRMKLEuymJsLRKgke4teNF4bWFlNpNUOdMKqJ3Xs8rRpCLixGr7VVf6EVbH9C36KX2SOXpF5RwWmZFJdRZzIiWYW7vlJqqo8kblQqpzcPfskdJyQhX36vpd0cXN7apZTMTD2OSRge19iokRS1W2uH6wk+eJhAk7h1a90asmzZlDw3tq5fjbq4ETPP6Zaz8rec0qcHef8mZ+UllwXxXK4KssF1XOlShhtSiC2XUh8SteZHpxiTHQ/rktgbYE2hJoS+BVKoE2YfEqbbh2sdsSaEvg+0sC6y6fLFjN3GrdEgH8WiKDTTpgBcALOxI2oFgzsNHlHMC5DQ7NpobEJpbzgO0AAtwH+Md3C3ACGqEYDpL0ItBzk+WFdclk/Zxru7/oGy/bMGEZgBqwhk1Mc/OyXl5racFzAHV4NhsMnkedrIsnykrZ2OSQPxsMNtfUyZIKrUSD3XS0gv1WY5xncL91L2IJHZ1qytNaCdj/+bQH8gQ4QW4/pgRgbbUYAdPIEzkiU1sGC6RbUsB+2jwt0cCzrXb+herC9dZU3YI4FsDjN/sc6/rI9o1Ws3/ut2QJ9/Ddgvv2N5uPLR/naQe700X+thxcQz9kEw1w/7tKtDP/A3icNPEdFVN4VjGId9q6IX/ysG687HMu+nkBl0+2vrb8jAvqSd3pF5ZcQLb8RnlsMEv+Z6PPb7QdABhyZFxxnSVUcHuALKgPv9FHKTfPwcJmu9K3lein9Ceus3UELKIMgILWdRb9lzI4W+Kuk/KdaKEeAkZRXgA/ntuUs0Dg+dsKD596v/PxVH/X9HVzsfTYuURvcimS3oA2pIKyfCIsnD5aLB/b4Z6o5sPMtkIjtV+BmneqcjvVSgAPFnhtbTOdvvjRGmvjq3jqUZ0F/J08Wd734/KEoqLXyiIp4rjdEQjc1FYGQMdtzeezN5u3rjxqhmtyVRNu0GAGIHzvte5TtQ9EPvHYR6o//vW68Q+0luKLA/dOvO/cp0YJvu3r3pbjl/QdkBLnS58h4HHsXZ0EibbuiNZYnI0HYAvWT1Mf3vmhwKxZlNg57059B5S7l2C4kC6v1+cfT/7rDTkInul7tnB9EHErla8tvVUiJQ74d471QNvkGQ3cVKLs9A9UnJ7sonttbr7S2x849TGhRt2uFylLITsqd1Cler2RTsajdbceygdXmIr7rrdca3Tm606s4rjdUjf3o6GZcBsmo9ggT8v91hHF0njPc4VrlxUk/I3IGPB6h8qsoNs7BcTvEvhOOzPn4Gv/ZbfzS3aCi/y4bjFgLY6mRktne25cfmzltYuPlM6lhrbMZbq39PpTN/eVZvpikdJtla45t6oA2YBqimehgNhV07W4aLpO/7VnBn+y+ZTiztebWseIiS7C9zZBss8oMbYZp8y3jEOAZN4j51kNgaIvIhP+w79oktuAp7+ufvoxLBIKjUwzNomInshcdXCPxkdZ5Tmlns24A5BjXDL2GceArg+sP8u+a78bUW3oKvqHdy4HdYCsAFSegPirhvGbT5X2uN2Z2SuvSn3rhq7I3LsFWqt95UzMX4w35H0IwoVDwPuJXJD9uO/Wj1W86OHJ4d5zy53pmoJtW4u8e3QZLobeq/SuSxQcYmO35ps37l4+/ui+uaOPzZieRHZoeqAiy5SpylZzprKDfqZyLLxXMoNAmhZp0VCsBd4vjDvqRdtkNdojVfEPecdLrSq6cNxtTMmUIl6p1nxZGMnCJPRloRA0gqComxu+78aCeliTeY36kyP4P3ALpVq20Qjk6T/CPG2tP2lzNKBpH94bzKlNTXKlZowRJUvws+5hrkiKnHIj6m8iybaI2Nui+C4iWVexmLLyJF/e4X+zngfuoHjOksZRDcLk9ORyIuJ7XSIsRFI0xlTuUcXaGCiWq+lAfvV9T8Cr48Qd01gYdOqF13n5iULNPXHSiW8rhe6OquM+KtB1VUTv5SI/Ywc6v/h5leEdegbvnfMHVh+r9c4DE5Ud0xrzvZorO3XOrkXo/7wbnlyXtVUkuVDz8hvEJdYRrKXo39ZqKLE3/8KZx9esKji2K9EXIYLoC7zDIZKt5aHNf/OahfO84z6u9N+VaBcIucIPqQuo1nZgXCDvjZZOkmC6JzAdW2QFFcaWiyvpZH4pKWdN4gMj6ob6XSD9CERDursYLa7Ee0VWOIlMuajA0g/EI5Xm2nKTa6jTul4AviInpSsJP9KoK+5FVq6VmjEzGlVZ+1W8GT/WWCzno5dHkvLGVvdk6WGb/0Xdx1oEW/eYjCPWRodEmgxlB3LJ7pHlcT3rjCwajoo86Mr25X0/XsvJxdOAujCkGuOTB9APGcN85900psS6eU7XzWku4Vy33r+rqn/Tymdk/2SytBr/o3PPSkQNhzkMqypP1y7IOuQykQ/WkjEpsmI1bLhp3eslO0uOCI8eyWlQsUC6JMstsljhnYhS09p+IzRiWhLMFUtyB6Vg52FrH/9znWdt0bSQaQfdflG/aJ9oS6AtgbYEfiAl0CYsfiCbtV2ptgTaEvhfJAELQlvrBDaQbCoAdaxrJTa0+BVnI2/dIwCYsgnhHPMyWlNsfKxmKiANmt3W7QAapmjoAUJYzXzub7oaUbLExYXEYDe1XLN2b0SKrtoiGTdFOQAGeA4bBcrM5gMQmHzZvPA/GyTu5TubC+rBxgdQFx/WbEKQBZsfNoSUDRC3FYSnbFZetpxsIi3QRVn4zr2cBzS2oBUaYeRLnhbot+QBQBgACc8GfEYm+DXhWZynrBAq9n/AAurS3IytF6SVtOAU/1vLllZLiVZg+kJ1sYAFAIPdfXI/z7HPa7ohWa8LMqYPAIqfUdreUp5Wqw6uo31aSRTK2PpOJ39LXlkiDZmCNpIvQNy4EgAIFjYJ08gLlPJpc7uRtfe9LHDVEmMiLqwsrIwtUYG87Dig79KGAIPUl2dQPksioP2H6xT6FBtaZAhIRXta8oX8GF8QEvRJ0G7GBZq4AE2QMYCdyAF58jz6AnKjPzHO6L/0J/oKZbIEY3V3xg2SiixbqDeBJWvtQx86KfBw5rLakYffV/9kes+W5y7PJWPXL4uoWIh0ROqO50ACRITyVdxImKqVTu5cnPqjFa8r94x71XXLjS4sNloPxjp1Rav7pUCuTbdt+Je2Skpfs0Ma0s3orAoqXRNIHoGkuDr9mAfoisayPT7fcbO5unTCXFM6aTJBsWltYY+oU33/+yKfXvib+hvK4wGi/c5xsOO6zIM9t3/pDbNf+ZGM3Ett8vf+AV1JmwFoP/EPfu9jxc+uyZS22JjRmqb855Vo81aNSepC/6StDtgnC9g2Clht7ur6grl/6c0byqSYAX1yrAEQY10i2SDbjFvmiA7FC5aLjMawwp77FdPRHTqxRNrPDa+ajgE/2ummY7FGpR7G88VKp0BaE8pPTKFU71bE9HgjGhFv4+XL5TAdqdfDDtc3abf+RCmITKyETqYcpKue471QaURTi/X+cwre++bB6Nn+pLTuBfZQrn+iRN9Eo/fvRTt0ZS1Ib3gitXNxOdKZGi6dG1Rc0/q3tl+9ODw/me2YXXrvaibtPnjH1RJQ3kSkRh+RZYWsL0yiVDGjEzOm7/ScKU0fMvXO7aYR7zCzr/vlr4z8+Y8zhzCH3qdE2zJ+aEPOnSfNX0p7W0BzVYA6faTp/od4DFgAQUwRA0T9uCZAGBCOfsCYsKA17ckcjhwBhptk/YbO8N3/Qz7UBcdrEGXk/VUB6jNy4zWqGCVvTHjFMVkC9O9OHn6tyEFzSi7eFmp9BksHgl8TT0IWGM9pzD0yFD3zBWU4qYDwDLrq0Ll58rdxc6gDcxDg+18q8b76WSWA/IsesUb15n968o9ufn51b34805ub6xJ9ItJkVrFxsEroaE5TQVOZ4Zn8Dcy/zGmA3awhmD9FSJic3CFVqyIe/KAx54qGajhuVOhpVHO3aFpHxGfoC0zt05QgLWpTxsM+Fha611H4i7JsLsJqPXDDcj3yhW+wNDl/8C6jToDjPJM+z7zL2Oc8B23IOJ0QwbPtsuShY1l/aVDky2V90WnF+hlvkhWStZ1b7BrEWmMxl5+PAbOiCDOVaj1ZqtT6RKL0imwcUdoqZiUTBgI8HfHOnjso4iLre/6snF1NJp0wuMYvTeca/rEFcY9yDTWqdJnIhzFZWjj3L73l4/f2fPo/qT/CjmL90HRRRR/V5w1b4ye+KXKtUAkT6bXwZE3ZAoDTxnynz77UOOc3xgwWf/Q16pPRfF2NNqr9IoSHioJ4o0E1LlIYCxveh7x73rAuwwt98P5gnrXHuL4A8n5ZCdljcVpukxVN8di160YSXa0X1BWDRqEpyjnv224kfq1iPKQhGBpFLTc0V8lywcitUq1reDmSHXRTcntE/AniQASK45CbO9n7uMiIq+SklXc6VhWJeLa07PtBp0iDVDJTXlVA62o06Ucr+WhJAa2Xyvn4KbX1hOJKdEcS9alaMbIswuJibW3XeayH7cFkf1gR746pLFtFTNQUSLuS6c89ImLlilRPYbuIFQUPD5mLuJ8+yv2W0OQc71vrDpS5mXUmfa6Puumzqagkd07JHTecuX9xouvril2RUP//ms7jDuvpSjGanj7eVx677sxR3dOtaztlYOFIHo4sMBQbJJxQOXaI2LAWQigrMFdQLpmvOLLwMMuNei0vU8fUpomdfdNtSsz9/1OsFFvk2f7alkBbAm0JtCXwfSKBNmHxfdIQ7WK0JdCWwKtXAuvWFYADVgsecBWQDPCcRT6bVzYUbGjZALBYt4CPdf/Egh0AlU0D3wFqADJZnHMAZLDB5Tzf2VCMKNmAquRLanUPdSEgB0DBEiprrgdqy6GpTGt78SbKD6CyXYnvJAAHgAfKhFYr9SIPS1AA6rDJYUNjARI2zcjAAv+tlgj2O3Xi99ZrrIYmAAf5UT+eZy1QuJdNFCQGYBbvMIB7PsmH+gOWsnGnjGiUkhd1ul6pqS22Xk7yspq/1JN8WzVAW2Vnv9vnIz/yQn7WXdeF6gL4RfkAp6yliL6eJy9svtQROQMqUCbkB5CLH23aF8AE2VjZk4e1SiCPViKI/kY9OL+ZJKGd6HeWPEJWlFF1d1dNYu+QEXi9/rvVnKV+F3JrwXUvOlrGAmXgXuq/FmX6OwFJ+U6/oR/TxmzskRHP5DukFwAXfZyDa6gvYwNgh/wYSxzk8XYlxhfkA3JmM05fhYyC7EA+bHAZj3bdw/N/RInNNgQbB30DAGM+Xw+nvzZb7xDINSxf7zfW17S86V8ZgXmxVFAoX195orfPn965HI8PBBHHjRVr+VSk1ChHosl0vVRPVirzhVh8MXDd2YnB3oV4JXewkEPh1/nR9efZD8YS5aFsL4uwaLWu0D127gGAQPO22ddkZSGnFvVTAtYmk15ht2fq/ZuC15pDiZ1Sc1xSRIeGSYXl8+QDJMQOd/yn3+J/8fTvVv/ZhuJW3Wjnn4584PitCw+fTDfyOy4QfJn2oH1+6+alR7/y2S3voF3GN9WZf7GcoZ1BPOn/HMiAuYPxemDzPXLDA0B8ev2+1p//sf4BQJ+XbCZK2SZYz3ghDYq8GROPtkdkxWA9FGrjdSi4dGy760cytYrTJVwz78v8Il+s9kqYsUw6tiy/99GqLC2EOHXIimJFkYijMb9ueiqVWdmpzMidTE68Rnp/wiRH4u5gh5f0jxZXzxzonF9NutP9HjHUhWNJlKU1z+jNAOe0EX3xewWyn5eBLFo4mKOYz+gTjL99OwsnGD9XKwFc3/7Wo9Nb64rJcXr7gHnqtTuarpg2H3fd922jyptUsfbJxtL4DZXBq5ug7eoV7zxQvf/X/kN04Tia2rQZz2N+ZY4IXqGLGR6sF0/4MyLSfkcEj9wolc2KYrEqjsEtDyy/6b/MVEcem6qOTsjt0c26lrmLcoxfrODjAAAgAElEQVQrYZ3BeD5vyfGiSrzCE+txGBh/5NsE95XuVL/ZKyKiW2UMFmt90adyN792ud7dJFkmq9tkEZJpuoESqSGXZYtndyWe/1sFL39Iv89JtsiG4O/hP1trH9vufDLmcY3FpMs4ALy+VYl5mrnrg5urgCu24dKkOVndkS4udJlCJqP2K5kVlUcB3Y3ikRDQ+2fVdj+nuC7Ug7FEPZhfeY9zbnfdcfcLzP9cf6O8LCbisoYnOiJ0ktJozqrnVDVH+SIuVFiZh4m0kHu0qhzYdMnFUigTJAk9UHyXBvEsnC19GffX/tu3gl9bqxtzLXWmTqfW62ItLniP8+5hcHYr95uV042Ku7NTsuuTvEYgzCArsnL/JvDeVh9CGpICwoJ3ejNmhf1xtVBRKdRVS/XeRhiM1urBFrm36tMAcD3fEwga9kR8tyoyI1muNBKNRiPiyyP/Tq+6cs6rTsk9zQ1yjne7OrKsqeStzzjbnsjddtO+5NMLO5PP4bKMgPRy65cgxooRAWXk6uvtzxeu0RokZCxDcFmrUt5ZrA1eNL43u/fTPEW7HFebKqaLU5dHoXhXbSmFi7Sv9d7V+WMTf1qJBRXqyzsUoPYlySz9zrrhD5VYR5I3RAVWKVZxI3yF49OK+Af1k3HGO//8UZUjtIJWXOKjB3rHgpGgUVAMhmBQVhFmdS4tiwLXdI0s15KdxYisFkLICBEEFVlEuALhd4mwSMia4EZZOmh4ec3wC7rm6lRHecJP1HzYrsxgbkFWCHXFgdgiS4O6CevRSLI6ou+FRLS8GNQ00QQe79BXeuwXuXJY9NsTcsW0FEtWw503jW/T87tEFHTqk7VVkyhUYj7g3cj71sbOsc9j4DFG+cTykznWkoyM4XQkUdvXN7ZwUi6eJmVlwfulua5SHbadPjgS9G5d/LzcUp1QfV/bqPk9sqToxNVcz7bFUOTFMRk7bdV8QxnsPsc+u1ukxbIfi4d+NKb8qpLh+aGONS1txpj7eyH9X2kDtK9vS6AtgbYE2hL43kugTVh872XazrEtgbYEfjglwIIekJZ5FdCTzQBgThPkVAKsAoRAK5RFP4t1rrPa/xbkZwNlLSjYYKABb60u2BRzL5pGfFpQimdZNzg23gD3XAho5jrKSl6UyzXL3/ZN9+t90yhxPRsVQAWAb/IFHB5f/w7AiE9yrmOTw/Mt+M2nBcntb3ZTYS0XdMlFrSy4FzCaOgMaWc03zrNjoRxsnADJKDsaqTwT0sBqglEuvgPUcT+yBzwhPxLXcw3lseQE9bQAH79Zlx2twJK1VrDlR8Y8w17LeQ5rWcC9lBVwkvxp01bSw1qNcA/losy0J8AOdbOEDEA6fQY5ch3twbXUmTJbKxe+W9LCWpxYqxYLYPIsZEF/a5UF/aTT1FdlYaPqBDnKSVnID0DNkg7c/5LHumWF7fOWtKM8to9QbvoXMqGe9BNkxKaY5924Xl/OUX4AKtrJurey/9MXaIPt63mQL3UC2AKsYRPMM2kP6mC1UwEhAfPJjwToSlkox5pLgvV+t1wLG1+eru+QOvJrVLBbdB6S0R6x0erEZJczP+pkqkMrsWS/7zUiXSZX2z19diHfmzST0R4vF3P9qKlPlbzoAzG/dt/J3N7ZShCnnADrrW5g3qj/IU4AEpD9dwNmUy9IAgiL8yCMQJNgud47OV0dfno0dgrrh83ghPla5prq7flnqrsqk2ksQwAKgSpTEvHd/v3bfq/6U+AsFrRABkUF3i7c33vXr7xn8jM/oesBWe0B+QC5c5O0+a+5d+ZLZ//78I9OPdlxbVNDedNB36NPVuQOyhKOgKq0Ia4m7IFGf1plGog4tUcUxwLQFYC39WAMNF1l/GLswzyI9sWygX6yTfd+ULVSP3EydZM8Xg66nLzpGc4HyXipJpi8Wh2S5nhYF6ipgNtOpCAFfyG/oet6DfnziASN5KCpz8hjd37Rb8yUG7WTjzWSIwIaO9/Q7fTf0eXcqkjex0WMyPX5m15bD1+bLwUz6XqQN8VgKlILViOVYOmeuNv7exE3s3D/qV+YvmvsxvNIzGbBXOj/dULiYpdSZ+RJn6fujAnmyLuV6Bv/Jzc2PM/k03EzNdRjju7bauTR/EX5bRufbnQuF0yqUPqmlGMfKa1OAhD9zNqFTuTcO/6wOvaR1wOkMnZeNgjaGkB+/aH0KeaBB9U+j8gC6Bbcl3UrsLfGibmt82/foeDlT3x18Z0VEQSH1+sEEQlZwVh5WeTey5GtvWadtKBPMldAkuzCQkLuxjQ5hiVZTizWFKcWywqRKnJdtNJ0X+Q7VcnDOSOrikJXZP65qFM+XAzSuX9z7ScvRfYiA54HWc18hHUY7cW8x/fblbYrMY8C2EVS9YJJKm77eGW3mZ/sNosdHXL1tirt/2gznoXrNn60d275919IK+KE09irc/foPsBu+hskgryZma4Vx0/nA/e4xu8ZB48ujlymheGOoBYGik3RUGDtFf1flm+oZfXtqJBDT5YLNXW0WVleyF2L8au1hju3VNg8X9GpWKPwDqaf0H94H9Afeb5GWCMqpzeZjL+SlRz75BKsd1v8uFMTIUDMnU3EKu7GHlJi7WSteGyTGQXfUJGceD0IeuQGqg83O67j9sqSok9EhUzAZOamKBYiZlyRFgMCSmMKyJ3SeBeyXD68WnGm5BZqbNV4B0uOl1FlXqP+N/LAypuOeE7t0GDs7NUEUV6SBU1JFjSrCkov12BxWVsohrrHuwhrPogn2hEFA+R8yTmcvrb7488spxqFYzOxgZ0iY69INEpOzY3UTie2DX2p/0cOaX4dEqEBsX4psgJ5oNyCmzbWDIwNa/XEWpNx2j6+IwHGHe8G5jAIHWJ4rQXc1hmm/ExfySku156VxUMslqz4fqzeke3P1RV3Qd4Dg7pcLjVEUpxq1N25xbNa1shVlOI69CvJOCDMa8w016WyyJiLd5TKih0xoWvmwrqnNVWYVeyLJb0SS7o/5dW9K2ulyEB+IXVWlgjXigT5btpKRlPOsMgS1uhLIihSIi9Q/mBtxZ6C9wLrC/oocwn9gj7LOKXPsL5ifKLEwjnWUXwyF7IuZz7kmvtlFdevYNyL554bnJElCHuUtTVoaPoUf6P76b+57PgN/9tTz8qaosOL1EdiSTMqkiabm0vHRepMaDyx5mNOaLUIWld6cuJSJFiRa6gX3Ehpr8weW2XBfbTXJcfXdyPA9j1tCbQl0JZAWwLffxJoExbff23SLlFbAm0JvDolYLWcrWsmFt8s9q32PpsIgDhIAjYJbN4hAPjdmmWzGQds5H8W8mgusajneoBXQAw2rgDl5M+GiPOAUyzguY772YhZbccLaaACogAKc41vpGRo8AJRm9EGRrFEvxPUms0ceVuSg80K9UNLy1qE6GsTJOPZljSxwD31sJYXXMexeSfWSgwgG56JdiayAvgg2R0L33GjwUaKTRfys0CddRuCbADZKasFpgFp2XSRPwmZIxfKyeeaOfrac0jWXZMtL2W0dSF/5E4Z0d4nL3u0bqJ4v/Ibn/Z++8l5ey31tZqwtBtg3F1KAFWAdNuVkGErIQRpA7lhLShan2uJDduvWkkj2/eQC4CflV/JJHZ1mtXH5DWnk/uQH3Kgrsj55R6WQFuz3Fnrr5TfamHTBgA89D3KxSYYcI42IMAyY+K0EuAPmtRoldK/AfMAxdl8s8kGBKN9rauor+u77XuUmQ00+TDmuAb50maUBeIQAI16MlYYZ5ARgD2UQ6CZSSxUw63FRtij75AAbOYpB3Lf3hMsjN8bfuHgcMfJTq+jtm053imfaqGRj/q6kw67xqrTQU+4OjEb6xwve7FvB47zZ/N+x7lHJmnSptwfUAJIRl60Cc+nPanDd3vQx5kvqOP5QyTBTlkk/Pk3lt78V+8d+C9fklulv9r8gKpcotyXuTZadGPfvLI8/lqChENYCL9vkgyDzoyZCgdb+3ky76df81u7/tXX3jzzhV/J1lcBw3FbwgFZYY9fKvrJxP7Vw1URFpAlm4/P6cSEtKvrM9XhyED0HGOQ9qH/MP7tQRsx3v5EHf2ghk5O5btaZaO+tDGy4wg6nZXqvf6X6QMQGrjUmNF179Dne6xBl+rVHfUaT/tBrijLiYwICjfqeFUxFHE3cCLSLHcqtXoqm44Vso7bKNaCqteQO5wwiIq88Et+rGPJRK7OOua53XETu6PT3Nrh06cdaWcnzwrkVf+MzdSDwt3SUCeGt+87aZOKjJiIm70n5nZ1xt2e5+R7nzmT8jfNQXTQx5oEDnXhhIIZt4jhRV/tXErbtL5rGCe0A/MkYCdjQCVxTDEZM+VEzOSyqdy5kT763osOkRoPPXfF9i9f8czJ1exqcTYxefAZt5rfF0TT5GVKwzfsnTvwC18bef9v/F21XC1JzdyGj/1b6HfEgcB9WdItDAxEJ+/Zn/7WmcdWDrxQDWOMecYxz70UEfBScnvJ3wQkN6T9zrz3gMbLoDT+h6X9n1QgbWntyxLJy4UCqx1crfVHJ5uB4MtB/Eg5SD2g74BpsrAoTyptQNpeAjBuEtwipJh/rDUEc8MnlZgL6d+MgWubNg+OrIwiUkRW7tJeFiGmgNsqA1YfBKSH9PFq5p1jx6a+Hu2q7C05SfoB7wVrLfmAHliUlcVZPWS6CeXXw6LvefJ31Ay0HVPQ+WGNfrl7MRk5+HNEYjgyrqjoXC4a8c8lEu5UsWzmuFf5hr/0/huIVWPlShtRbp4L+Ml8D2lMnR5Uot+lRbJ0iKSojMVfqMm6JoHdhpzHNPNocTPHXM/8z/zMWGlaq9gHffrBk77iVohadMoKrl3Vl1jE87OVes1VeYOyCBYRI7KACTsUN7whb31yZxVUBOzWg0ZjW0K++S9znHMzYSSpmB6Mk3WFCafjTHlH7aGVe04OxU6vipQaVqwcyXmZGBZY0qRv7/yy+/DKG6Zz9Y5RyYwxyPvtRS7KNltWqJ0Zt8gitvTQHT3PZS7b8sv7frVjMdqTev3cV2bjjfJt2XruFlmvqa1fFnD9ceUFIM044vm4frKWnXYtaEXW/vyOBOiwEIG835vWEDVZWAQaV34sXMr21TOR+OpRWQ1oEna65AYqTHWVYrLYySnodE5kQCJoOMcmnhk+qUDbOzsGcpOFpcR2WRM4IiHOT9wiJsLSaqLUiHsZuVDSKGvkM32FRCxd1fMiHSI4EvQI3dMX5GN9iiOzonw3uqp6ea02J0dQ5fnT3XsUQ+OxbddNzItcgUzj4J1In2ONZd0+sZYmQQLwvqWvoBzA+okxy5qCdxEkRnPMIqZ1eS0qJsVrdt1y6vCJR8dOq/55jUEsgm/SFXnJZ+TI13c/tv+e5xdF3hzQxPZCKRcPl6eymWopynoHQpO9DO96ezTXs/CNyst3XG8vU5IMWFoDb7Om5H3JHNMmLVqE1/7alkBbAm0J/KBKoE1Y/KC2bLtebQm0JfD3KQG7AbXAPWAHwAMaviz+2WwDZLCBZ3OE5jwbCRbrALAAb2iOsggHqGVuBkxmQQ5gajXu2TxYF1MAstzPpou87QaJBb3VyLea960Le7sDtoC9tmzdUquOxYybZFPTaplB/oC91rURGnuUFSD9TUrU126E2NC81AbCgvU8n2evkSVrWu0cbLY5zzk22wImm0AbG0rqRKLunLOyXL/1PGlgNRwBtthcWQ1c2qLVSoL8IV3YFLJJAxCiXCTKxfVW9XgzYsB58gUQtSRGK5hry2Tz4rm0sSWVLMnA74AxTVcqStZyAtctbCApk3W1Za0nkI+12KCuyKY1P8qOnKyMKYsljyAhuIe8AOqtFQWyGjTydtMkK6SWZyugT0t2XRI1WbeuQDbWRRb1abr+WD9nCQI+OQ8RR99mfAAS0Y8oE+3Cb2xm+YTQwB0IMidv2h5NZK4FnOF35Mhv1jUUVQCwJU/aFzkyhiiLBQTZkKPNDxFCPbEMoGzCps2y3EB13Njtd0ycq94kIIO8mmRXT33hqVsbD+cvc48ciCcWcguxTC5er+aKkXgq8PyKFwTVBS+br/newcBzHxTg9ETFiUwJZAvif/lR634B0uJPlXYoYfHCfMC5VmKLOhhAwM2AV/OHjQf52jgym4Ok/5mCF392ud51IuEWGb+/qMS89M83Z/JCfLSyrzJxUoXYQYNHJXIRAOYm/3Hz2drbNl++70xiq3uo4+pv377wINr3yBqC4PwB2aG8fq6/MvvcOrmw8ee1Nuvp8BY9aarTb+k/ACrvU7pu0wOZQ/9Awaz7L089OS6g8CNS+P53OmfJipmIqV0+5EymTgVjR6/xnr5GmuMQf1eqLmJhmxSMXLrI643buCpnhg8vNLZP5YJkV83xkor6uyJctiRd7SReb2KeE5f2+GC1FtSrpbocfjnpSCxSWawZf15gUiFwJ6uBifTHNH855iFxAbeprp+qNCqfkNLsNaXG7JtLwdS5fP3MaC3MCTBVeBg9X4Dv20YT985FnHSfrC3U5g7jnT5MX6YfABjRnvx/scPOVVzHdxs7iHFF/8ad1k8oWSJEQLDCDcu6YrUjZURUmG/fsPeCZEXnUu6BUiL69Vw2+TfKOCcAeLnavXM1iCR+U/k1CQu57PjNuTt/QSDpb5xHqF+irOd/0hhoft9kaUG/Zczfby+kpQjCTBIQ/24RWU+Oxk4eUqyG1b++S4Yyfz9HoCDvp0RMfEP988C+1KH8fHVwoGH8esrNLaw2unqrsmhYqPUbBYk+NRQ7s1xqpB7Q96MKuj6rul5IUeDllLxJXqwn5IuVBWDiuBLz189Fgpq5ZuWQ6QkXzFe23qUJ8XWQO01XSriGwlWVUwn31ZaTtau8Z9JPZa4pCKmXUYS7ILID8JF3wrKCb88dNKncnqAg7D6sRCJOzvO8RRF6feIhouozHaIysuo6cXF4C3o1zMniRmUK5bLGWZVlQ16/v9if2No7hvcKYxlNbuoBWcJ33t9JjYTZnshst0iLbrVzcl6xgHt9xUwR2UKsmvWDeR6CFeuKJlm1OVh9T2fSaLz6jXojUSx5Sbms0rsk7NOcLWOpsGKqjZiIOrxbpSWAsl5wJc0FCkMTiKg0CZEYtVFTca52/bPVwC3J7dsxxbJgvj+rto9NlMc65PJrtTcyuyqSItvtz8qKxcctXXrAn/w3fZGpTxcbqed0LSQ476aLtnsrUbHeltvkAqp7Z+FkVq7zYs9nLhu+aenxD76Q3mNOJ7eZ2Vif2VE4afavPmMJHFxPMV/Yg3cgdhMk5gAEx7uSdwDytv2o5Zb21xYJ8L5HQYQ5t6npD1khF0dm8axXLOcaC3J7dJX6ztXq7345Fz8tciGayJYrXm8hFEh/WO6NurpHlt4pAsyRtUUGskLAvGJa2GVZM7/+4lKipNVmKPIDN1CeH61nFN9BY0umS0kFu6+7q6LWsrwwm67Z1tYjreT/SzUc7Q7xIJ9Vmurlpirdm/8xWVp8Xf+fVudhrY71KnOLtcamfzQt5JR416AQwLoAKwq7PmbNxXuC8jAWGc/cQ7keFPHSNbBrfjQ/n65OHe3fqfozT7EOOENcl9mTvWOPfPI1D2+/buJbsqzIzRzv65d89ouMYR1y57rMW+dzylKSYsCxeqXQqag5vUo6ZZfSzbUc/3y3VqgvJcP2b20JtCXQlkBbAt+nEmgTFt+nDdMuVlsCbQl8/0lAoKywmo3Y7brPfltYC9gCxLGJAISDmACQYuXNnAsQy0aJ3yxpAJCMhhyEBiAT7lA4Z8kCSA7yBthF25CDPLkG4oJNBAA6C3nr6okNzIUIBDYj1mqBXVVZ2vVJU8+VpFhJGQGJm8Dtev48CzAJjXA2wtxP/XiOBactKM61raCrBdY2kyTkTZk5+M7G6FElwEfKQH0BZ7jGunBCFtSfzRObKGu5ANhlXULZ/ACn2ZixeYJsob7kAyCIZpe1GOE6nmWJEu63mlvc37pbaq0LZWCTZ9vUXsf9tq6tsrdaZFZO1pe3dbllyQM2qRAtto4AjwAhbCRtecjDEjHUDZldiJBic9eqnk29qDcbVfog95AXMs6ZsFo2rsRUPkm/5F7kay07Xo7mP3nRllzb1B5Vspp8tBEbYTa6AGa2P1Mn+pDVToUMg0CgvZAJRAQHY4Iy0V5cQz9suj1QQjZsyMnLukPjuZAR1h0VeTEOrdYgz6ScVkMf0BSisOlqoBqEuVOFIKsoksLjTFIAakEqf/yU7Hdm3f3O0/LyVNtRSXpXog0u8M1TzIqgr7ycn/a6ZFURfbYryP2xXCUcL7iJ2j+77q+tpjXypLyMpWuVaDvKxJijX1rLj1cCytLfkB99BkuCzZqZaGl709VR+gxjCKKEPkZ971E6fyx6mbvORPrvu7xxmnEmME8BPJxz5k7vQZMP0+ar9dc1r9V5xtI5uS7p+6V9v7byjYfvJN9/qfSUkiX6miBbWu5rRspn0ajcfDB+piW/JREQgeIDABgdUPrwen02X09fx11VMeXmI5L54iYhDUgQP/GB6Cf+U9ZZ3SZw9g5d26wfxInV2C6HmTOlIDMiX/R9QaR/2jPZk/VGfFgNLdf3QV7IZpfcQAUlMRuKWyLXHr4jf1BCmoR2ykuWbE+W5J58LuUEz3dEw2d3xN3lrojzbj17BIA/6SUnDuX+42w1WFGw5eRXysE8LlpkNRBX2X2BscnR1dqx9+j7fUlv+IT+Zx5nTFq3dXzSX1/qoL2Z22hrS5LTd/j+s0qAQRuOuoJtzPd1mFM7tpgjl/OqePERrdaOiK073De3/O3Lnh0/Xfe85pgbef+vB09O/Dz524O+doMsRO7T53lLEJFrF5r7zt8E8aZ7HFmNhHzyg74HIjB4DmPg95X+D863BnKPOpW7L0s99Sf/9dZfeCXj4qUleIlfcdfzTw+9M1A/mZMFw7jcQp0Jk4dvqwbRxVKQWhA50YtVg/rYqtxFHUx5+fsz3srT6serfweyYnOpqC9zE+8t5rTfVXpIz7yuu7b4y12LS+Z014h5siSjJI26vNthMnINVVashdO9I/dExut7r8o9XeipLMx8o+dOt+pEtyiA85Ri0AA+NuN09MnYQMRDKRLxQrl7KqlRZH0gLsQN5U0qHJPrJMV+MCIyNNEFMhmpB5WqDKJqtSAnQq8ol0sXWmPQtnZe5z3A8+jnAjTlpsapz9+Uvf+YHvDuuFseVcDyLGMUooV4KuttT93/Qom4Hk33Y5vJCoQFYZErVlPFYtCVTkY7xFLICsSJR6P+alipe8JvsyITnWg00pBrq6wrayq/ESzp/JIKWRUeWosF/z97bwJv2VWWea+9z3zOnae6NU+pzBMZIJAAYRZQmRUxqNDarT2oaOOHw9cK2k3bn90qbbfdrWgLiGArpgURQoCEDCQkIXMqNd+a69adhzPvs/f3/M89782+p25NCT8k4exfrTrn7rP32mu9a9hrPc87hMmLvPLMEy6rOB2uT4uBpoWWiIn95bBrKqjJ577kLxFcuqd8hVsIerRgSDrFBnKKc5EQWXH7wcoFgN5V+k28EZskxU8vKxUwPlnXAOwymb4W2Yi0ePInD3/ijY/0Xn1DXcET5qXQL4JJzGnZPdV9qdtaOuC6gwXedyQILObKsZZsvqRPwGbedbzLzQJptXaJF+37/Tv9izUyxwozNl71i5N+o6wpSt+7ZCFQ8BOuJKJivwiGHbKwGNDnjAK7rE1lg0vkAik9e7y3Up7P5udPKp5N8AxZQeaA9wLz5+QKKSmSgyDVZT+Z3ZRKK9S9emgi2ShXFzMiK5rP4+AdijLHuR62N9D1nqssZHYqvz65l9qc7a7eKeKCvkb/4N3Ce5fxRJ/hO+96U0RiXcZczLqKPFkfsVbgOt75jGGuYf7n+zG5yfI2v+gwlh3p6UP9D4vAWVD9mgonInFeV5zOX/Hk7Rex5qNmkJXmJu6z+m77HbPIZd7g+6gEI8d0ipTTUIiPllB0nj0HbXVWBZpzFVznuo4EOhLoSKAjge99CXQIi+/9NuqUsCOBjgS+RyTQTlZQLJ3Telo7jaXDCAubW9m5kNAixyoBUP4HlQDwuIbNPJrVbBAAWFnUcw1EBIt8QF7AWRb2HCz20cpGi46Ng7k+AUxiM8Jin40FYAS/raala9r3y8BiE3MKJhtu8eETrusifmcTQ7nNfRLq1eaWCoKETQPlMwC2Vbzmh8mC38jDngfIxncjBKgr12BJgQzYhBvQbabq1IkNE+UA6EVmZonAs8iD30lGXJhbBDZhyJTzyGGLkhFHbPoBjOMAGKCyldHOx+vCd8oHuWHAPNdZPexeymUH95iLKc4Z6QGYQ7tiSUG9jTwASQSY5W8AdYgFwB42kYD23E/92HySL5va+DO4r+nWSMksKsiHc/yN7ADAkAf3I2fIsbtc5eA211hMuYVvt4OClh/lP9th8kDutB19ELnQPnFLGZ7PNQbk852xAHhv44J7yY/+zMaZzSr1ou8xfhgTyIeEbCgnbQ24x++cp76MFerMJpr2M+08rsc3OoAPZQRsZxz2Hq9E1fumG1tOVqMNIix6c1F1ursxVyr72bUbUof7E4V6lyDzUi4ZKcSFsGwnh9dCtEVUHE56jVunsz3Hp7yeMVlWFNtANuoDKUI5sSCgznZQPuoWt3CK/Xzar8iEeQHNW0iI9gOSCDI0+NC+Pw8VKwJNZfqZkUE2Tpv33dN1WXVtMP2RnkZph0ia9wMezisOr5EVXCNAMJV0cuguFz5H+9bfJlc3JwXMIWesNn5caYsSc1FvKZFPP9ITVwpeKp7y/SulT13Tfe/hm/u/mBV4iUsw7l3NWolb6EP8NjUbDE5K7mgbUwf6RvOQTv6WbrfwI1cknuiTIcTFKqM9q0laCBoC0BuUYcQxYSDz8toxE3pdg7mUL6fkGfnjj2qlWjBbazj57XDZJOr0QV1hs/0FhQaoV6v1RNbzyxvSib09fkCABj0AACAASURBVPhY2vcOXNfrY43CnGwEgvdTl360IhCeccu8/GdK719q8qVjzu29bKL+wKePVL708I7CT073Ji+iDbifvk6ho3ZXUC3tbOpP/2AsMdb5m37zcqV3K+FOy94Vy8/DuqIsN1ATw33umKwr6mq91Q5dd+tid+6bjaT/4Kax8bnNv300ri1O+zJfYfnHATFyp8pZg6hQMvLRyGFkHfz0eq/xz9ZJjZgmXyIpPJEVRmpDYESPLnw0nK/vFS3UUMFWxVmvl4uoDZIp8jxFg90sN1at1LM8qWdR1rTclY0ozYgAa6r9F3w30ONmBwioC4avfvUlOZH53wLhH08pXu93kKywkiMQns3cxDtj0o/Ch+Q26HgxWXjrMX/967H0mGyscaG0uutRqmmhMNcVuMroyJa50oArJ3KXXbzw9FP6HBfRsUVa+19WzITZL4+8oXLbj24Pb9M8q6DZgYJo14TnRyIn6ikv8bDiPZTknka5elMscRTloqz/JjQnnpAFRkmBKGqVamDkebuk6cfMNQbSy4NapLA+lWp/cjK3Pff05Yeq27cFUVLrmChLPJCcrERiRNXtupcxTmI9sypZNbdQ8aq1RlSqBNlk0s8Vcml/vlTtU+PNJJLehIiVrAgXlm4VWV9kIsXckBVJvRkMOeHNKwB3SR625H+n0bg6Kh485tLTgZfs18/MpTsU/6Mn4SVOyHJmr+Q6knDBkIKZq6wltyEzhkuwC67uvq86URutfOyGj55KViy9d02rHaKCee7NSrjI2qL0WgXWdpvKB5uRg4rJLvzhuDXVcVeSpyAsLZ7svvTuF8098te6DjkwR7Jegiz8ihLrBcZaSfPwd43Qe5bD6nvmtofu/lR07U23mKUs44r32fJRLXqDR57InehZ4zbkemsnZA0h0iIckKHSrKwnhiqLmSG5XYKMiOaO9yRP7hvCzdgjikPxSnSansHYm1nulWXG9ijMlqTE0K3rskU5KlN8B5fKaJwuZOVaShT8yqmPtQHzXZy44CVi68y4K6XlcpOHyJENcgtVajT8nv71c70qN+7ZmJdZQ92pxNzGGoA9BPmjOEE/Zc3Ey4F3CgffuY93Cusq1k585/6m1aq2Pw1ZiBxSPIuCYnqsO7Fn+LjkcqVImwtaQbV5D8YtpZvvBaX4mnAlAaGI3IphEXp6CeOUMvZOoM6s9VjHU5cOKddqqM5HRwIdCXQk8EKWQIeweCG3bqduHQl0JPDdlIBpQ7L4ZlEOiAVYCNCAZhyLfTRpP63EBgGt8K1KaNyxUWgCJK3rbPNEPgZIszjHuoJNy8NKAO5sHgAFAJK41kBa0xgD6C6JUGlArLSEwTkATub/JYKg+FjZrf+5Ltd7/Rb9DQgIwMs15vca8J9NnVmOUC+ezcaBI+7yCDnYpso2IvzN87mOclq8CJ6PmwjKzXNJyAagGSCfzRKbFNs4kZ9pY9nmnDJaXdjE8J3ycR1yH2vlTx3Y7LBRQnY8AyCIshgZoa9NEJm24neeb3UxtTn+jgMD3Gv1WwbiyEhH/G8jKzhH/pQTYB2gkmexiWOjSJnNsoTyYXFAH+E+rjHLEiszecWtdSgn9yGXOCBufyNfyss1tCHPBijMuvp83qWGuc5IDiMgzHKhVa3TflA+2pi+Ql+GZKJ+9FGeR5swLvidfsx5QBwIMoBI7jerI2RgdSUPyBXqStshi4NK9D+uM9CdtjQLIQpJf+V5aBPybNP2hTTgHs7zTPpGU6tQWvWNvYuNtWPF8IL5WmNERhY9hagYXl9/6NjO1IVdg97JsDs3kXHZeiPRCKeCVFJeloMnIt+bm0sUdi4k8ncK4p6T7iRyaD9oM+RAXSgL7ijwNw5pBPBurslWufWZUzFf8Zy0PgYJh/uUn2u7mXozroKm9q+0xvUduf+FEv3Knt28reKl3/T5nhuevHnxsak1wczBrqi4uVduobKyL6jIM4zlHbjkNsW2uHitf2LjxOdmJ90X+6jvXyvRLmgOQ8wOK6Cs6w2eAesV72JmIdld6K/NLATpROrywoMjAioZ67QdIF77AdH7eSXAOvrmhFwETee9UrgYdX9SgPGvxm94LLzigldFdw6pTWQi8oy3GtxBSVAZxdm9f7qx9cmZxIXy7tQd1mtBvu5n/FxWnu3lLVta5imBnEkv6dcUMj0p9/gCmYIgm03NR416kJGmbSLjn1yTCA91Jf0Dab/Zf/5BCQse2tTmBx5O375bSYTFSmxFBh0fKjaOPvDI/H8wK4XSz/3XJZdJHLEA2zbODaxhzjDCmP4C+Nne5itkSBQN4lbM9nfvmunvAog9hRQS7f7pIJnYJdLi3momNXvph1aQFeTH2PvPSv+zlTnvL8AuiAwjGyEemVOYP6oJURR/PxEdUGOcfMtw08c/15nrP0Oiald1/2rj2/MffqLYOHydXlX3KkrDy1ZUYAkc4xwWaMwdK4SJi6nvBGnR5qrK3uM8+x2yanhvs0w6K8diTRdbOv67AHbeyd9UYo48hUxpq8cZ/zxLUGQjoxfVN4qH8ps+MZPq+/qe7h3vaPjJD4y6Q4OpTKXpruhYbVMzaPnJtevcJWP73FBw0r3t+K2X5oPi0GR6OKW4Mw/3BnN39NbnAjVIk3AgBoVIi5piUixoIFRlcSQrBHfcj7xCKuEHyjiS2yj9i0pCViu+79VlYWHKB816xVzXyf3dLO10jxKuaC6QnPbIguJJuc66XG60Lnh08SVXZP3Spv7UVBP8FyEgLmRZfMyPzMmApBNq29ORIq5UUZQhyb5UrR9PyZ1VMuFLszsS90JwbWJuaL6VSygVvLl2kXOounDQhEiMdapjv9qznk4kRYBG7oqoFBwMkrvuS/ZDAtystE3zi+alKCtripriWEyJrBjakt3tRGI1iSGRVlfnvYXrRtN1gNn5GLFoFoYonTDmrO8zL2I5ueJQDGc3UJ/RXDnnCsGim0n3u2/3XuMe6b3q4a8Mv/72n9//sa+/avLr3APZj/tQFEiQMbLpALdnHFmn/ZEOx/x1f6uNli/0vERl+vDopXu/me7Vyyo5sn2iX9YUmVxv+aisIuQOKpWfPtoXKiaDH1RSZZEEE3J1dFEqr7lBAbMbtaSsA5ZJiC59V0BsH1dlS0eYcBVZYsjqommB0UZWNK9QardsPWNAo2dq6XVj7REeHHhqeMt0Y2jLFOsd1gDm3ok1CHsPI74Za2ZBwTjhXc7zITpYI5CY29l3GCHOeon1WZ+fDEsKRj4vYuQKpZHidCEzc6w3KeKiW/XaomtYk7EWRN5HW89quths5fFM0fWNcRtUSqmGjH4jWVjEjjF9/5ZSh6xYIbHOHx0JdCTQkcALWwIdwuKF3b6d2nUk0JHAd0cCpgXJBp7FPUASIDwbAgBJNgCcR9OIjQDgGyge39kI8DfzMRsUNqIAYIbygYwAbALCA/qwmUfzCrCVA7CETatp8qE5xd88czWtf55ppMLS9qlRlh+CB2suMzrjctt5LhsMNsOA+2hhARywScblDHWkzJAv/A6YbNpeZn3Ap4HNPIPnASyzQWHjbuA/v3GOzRP1Y9NEvkaq8Mm95M+13GfAjQF5ppkMoEa5KT/y4R7u36KE1QqAMIAXGy4DFvW1mT8gAHUBTONvyk454ppmBgzbltPqF9dQN0CXT7uOMhvwz/PMnZGB04AjAO9GBkHgUB42mQCCyMSewTPtu8nCrHjIm7YxMNJcMxkwaC4BaDvy4VqAa/reNS53YcEtPiX/RjkDFMnPwNdz0dyMA6sWH8IsJ3gOO09AaeszbJIhEwC42fzyDDbVlAswFHKJzS1lQD60Bfdy8Bt5I0v6p8kbudEfOJAfMiBtUWJc0S8pg7lYeam+v0SJ/oKlxcFA7n7++ki9ePt4vVfKg1eg4zfr96y7N3tDSpYUnktGlZww64Hy7INBNhH0hpXefFT56oHUaI/A/p0iK6jDnEC2pkb2KgfloF7IhP4JSA+wfZMSiPXpLAxOk12z7sgHl1LkYQfPR8Y8C/k2y4PFh4BZZAxI8wkl2mrZSoFr5hP5NxxOD388G9X+e9Vlr3pJ+MB7/nXmj73fq35gRRl2+HszP5z6wsZfTv/+4wJbmXPmBNgBUk4J6Ht71afLqdEEwNkhdyfMi5Jg/kf66rPSAk3h8gULtI+sUkFk+SdKjG3muzHq8pvXfrzxhr9/a9+D0TWjxWglpnNb8NqhFycecC9P3OMGPYbw0iEteD6+WQl7/qge5fuKjf7uYiOzPpVOZwWQJCu1sCyXMTIu8MrppPxA+d5CMuEpvrA3XqxGkRS3vZSXrOn3E6lkNJ5J+VNZGWWkEz5lZIxRryYRKauB8Hj1jnBf6dMTCg0AmfxJpSXA+5mDec/c5tgYjf9uBCfzGHMWRB3zAeDna5TM0qEt21P/XOjOfWz/9nWDMwPdEyIvcN3VfnxWAPxf6STkUHMsxsF7yICWG6e72m687s13zB396rT8hT1jvbaACx5NSr1Z3+3IeG7DwVK092Q5mhvKeJ4087sFIDeCWrio2VyiFlrtucXt+XfPPrHw+/fJFXy/bJZe1qZZy2OvU4JkMyu3s9b7OVyA7JlHkDEuqt7QnpcgRtwV8a7h3dx0nfWdIE3Opcwaa+ovTxRf86f/MPZ47+XfSvuVh/1iY6sfBdsE/Xv5RNEpiLUrK16L66+7N+38ikI8pBN99bkRkqwsvFyjTJvt1XjF+qpMni3SokkA41pJn7iDyqnNJHNPxgihgeMyhmm+zxvcc5oy8ztrBvrsqCwrDqtMi3JXdZ1iQWQ3Zfe9RDEs3JDibhDIOkZWkB0yxYqAtc5pyQp77kKxWhNDMV4u1w7ok943rHG5VT0lIRKjV3yd7CcasK0pES28I5asPryomk0nxojPUasFNbnAclcH8w0RFrw7WIOxZrtIZFWfgoOLtOj2Vf6LSmFX07pGrsqa5VZfWNcfzIwe/5WeipueZ1zzbuegD6FwwPzOu+pnTte+ctWlppppuoPa1X2xe7z78vqBwrbd+ntusD51USWRZe2ItQkEKO8Q3qfxdcXpsu6cP70EWA9ANEEasxZgPYLZtPMTqVc16t7Q3HhBbsNS2zJd1Ubf2rm0AkbXkqlgSjEZRo89NVoU4ZAW4cBL6DLFdAgHNszq3tDJHdNRuWZKNBTMSsG0d+qaXoH3XLf0UtShc1NSJTKln/ZS2pqadmYs0SdZq51CdrXf2CQ/xL3LCmT2ya9euPuSV+15pG90fm0qV/8B9dVhvZt3Sn+JvkR9WUvx/kdpxPoU7zESY9csWykPewrKQJkhIJquO5XX1bIWuaR3dKE331uZLM7k716YLCi0V2KT4nIwfplPyY93yz4lxhVza1yhxqoBISrSR9ZQzYos60jY78iB9Ut8jd0ugs7fHQl0JNCRQEcCLyAJdAiLF1BjdqrSkUBHAv/kEmCFbRr/Br4CCLLxZpEOGM0nG042Cyz8AazllaEJvAJikgeaVGjmob3JQh9wAWDXwEw2Emwy2DQAeLKJ4Dry5gCpY35vtwbgNxb6bJp4LptrqYHJFUf+Al27tNVp5cczATxNe/9H9Z3NC5sFys/v5GUa8eRtgLqB+Wy0eBYAgYHknDNtdzZIlNFQR64DiDaLBUDq9l0Lz4uDJOQLCEEegBymVc91bMZwOQXIB2BrJvDxPHkW91ie3Ecb0jZG+CzrxbXqQrlNA5frASZsZ2UEg23GDMhHPsiWZyF3ztPelInzbP5M1vHyWD7WNsiI5xtRwX1xwBP5sjHkHLIxgoJyWmwI6kUeACu0zyFX2llQ9IY1rjpOvrSxETmU5ZRdI5VpO4ykMkKF/mikGb+NtcpC3vQjNp7IjTYCzOFvwAPuA3xH85++DeFHe9DfyIf7zd0U+VBf6kOfRPuOMUadKbf1K+ptVh7cT7kYl/xO/8CqhTFUrIYus3cxnCgHDU/RC3r7o+LYvMtctMaN17Ym91VeG3y1sr58sDrr59xCLl+eTXUdrCeSUvP1dgVeAvBvmgDb+lztoE3MJQLPNGsivpuGNn2DuizncQ6BtxlP71aKWyhQZ+SLrMwKpVmmFmlB/owXADDaF2CteQjQuPLbuQv+8Hhy8Bfmwt4Ta2brJ/aF25hzVhyyvNhyfeLBylWJx9ZHty9ZkdU+05Tto4vJrvcczm343SPZjTc/2HdtnNRr5jFcmxi+fvFbXVese/gmBf/9tXjMgthDGEvICBJk70gwO7e1dsLTswr3ND7a/99qPzv5d23BwI8p5u7F/u4VZIVq9EXF5f2TStjd9XDxh3Z7qb7RSmqwT97s+zXj9QqwLAvIzCT8ZFW62CUBMEVFrSinM8lcOpmIqvVSypPqeT6dOCxN7WNyhTOdTCYbuof+yPjB5xXlfJ0SwH+0NnPz5tHMy182WXvwxJ7iJ/cTeHuVgzajXwLQ0uZ2MG7p77QrZM4PKTG303cBrOJkBWOAa9vX8zMiIZ6upZOl8dGBXU9dvvVmfX/nKmVg3KG6TT6muXo6EBryBdAVEokJ5s35RNMtDSQgoGwoSo+JaaEgF1q9SXfpUDLq6024vr0lN+2Fgfw+RcNq626B3/O+71eyMllR9zue8TfUh9M3HJuqP3wocKWjIi3WLxViuSgv1x9Y4kA2Mr+tOL5TVhbKlPmPQkGi36zEPMJBX0TjGLdbEBWfUuK9fkDpOVlWtNflXP++Z+BGxnaxO3JPJXK1fDXKjtSibDeEhYLYO8XTcDMjisN7opGozSXdXNTrLlnY6eRO6sZE1GB+/ddK9L0uERfUr+7uuD6EfJS1hVnqVdXn1arLawOK13wXnYGswNoi0rw1JcuJ++XOy13bfXdZcT42Ha9uHNmW23XJ+sxYs3yysoC/iruCIn/K9JDS8bO52Fo73B2KsPCG+vKNmfnKcQXa9kQkZkS4eLVaY0hWFAnFqaAOE4pRMyACIydAmiDclUwqOcXY17WyQPXnwkgmKKHMRt5OGAs3q/I3LVSrYe6yqfqaqD859X/kAuqS3uTMJZQbCwvmLT8Mf6BrsVJLBg0swTi2KEEUY2nG2EUZ46wHpIViV9x+IjMaPN19Se9kevCRPYUdvV2NRW9N5eTMy6bvPSmrGPpetERadY7nIgG5hQrlFgoLC96TjO0lwkJHSPyEoLYtqLiKgkr3K/bEtID4A+lsXaGMXGnmSN+ICIG1sqaQpzTni6SIeoYXa2sumJgXeN+QS6RFBZ0uKrZDVJ7L7p0b79kvEuGoRtEmERWs71n3nE6pIV4t5nVTZrK56KzV1jMyvMjlomp0771b94xedDLoG53b2T28SBDxbeq4ZcXOkMXRcjeiLLykWCuwFmIPQTnZJ7AeszUW73fWxqY8wlzMuyul/JJ+V6ioHArvUk+kFFj8aeJ5qCy8Y1gboYjyCiXWG6xP2teVzflMNyw2gvoIU07TvdYztWVMmWvITv8/ay/oXNCRQEcCHQm8MCTQISxeGO3YqUVHAh0JfG9IwBbggMEAWWwuceEB6AQAwOLegFTAJwAPAFn85wN6AZJwPYtyNgucMzCeTQGLdDYQpl1PrQEDIRbYRLDp4BpAMDYegL/t4KlpmrNhAgynzIErPikF8m6LlWAWEQC/lBFyBMAMrSzqYgC9WQdQT9MUi5MYyIC/eSb3UG6eaZsNIyysHnyaDFfbkMQtQ+w6NlCUm3yNAADoY5PEBhSZQvZAWnAP8jTXWVxnFhyAFEaw8GwjmdhYmby5HxmbdpfVhTyMuGn/bNcEMxdQyMbiUrBRA6hmkwiIzAbRSAuz0OB9TV5mAWIy43dzdwXwT3npU9SddrPnWx14Pv0Q2bNJ36xUdoXL+hV4XajWA9Tdns0mFfnGwVSee7qDstGvSciJT8pD+5hlgcXmoM/QLtSbsnIdwA7yQ64A4PQ/2op2hWCg7ZAZ5QK45Dx/AxZzP255uIeDOtCe5EW5sKIwqwt+G1NC7pAcRoAcroRubV+ikc/4Tk6pvbX5ZPnRgWB8bMifyBWS8wternrgYPfIcMWlUo1kIh/4vp7tjUlo5EOZz7aRpixYC+Ba59da11N+0s1KtD/5nOtBv4DYM0LhQX1HG52D8co8wjPb+yFyRqOefsA8sUxY2IOPpQb+UMGF77jfu/augiu+q71A9zZuWK9M36IEsfplpb0C0gIBfY3f2fn/7i00Fu8vJgo3P9R3LX1v+dhUPuTeNvG53E1zd72mPNy49WjPwIrfWxeiickYfErxQe6X8/nSm+fvTyi2Bv1l5DL/qavenryVeh8UaUEfbh7dUqA+GQ07ufFyF3p7CIrM6Y/Vo9zOctjXVwz752aCFy0OpPOFRUVPrsgnlAiIKJtOrUmnhW2G0aQsBPDb3yVtbaFWYd2FUUl1lH8KNy4/+Sfk539egYqledsIegoZwB00yZkXmQORN/O3gnAn3j+cfskFXYktf3+o8vlfGK9+8w+j5bAtzeL+mBJWX4x7gDOzUGNugACgn6L5+g6lLVbHtk/6f/ygLLxP5oqF7BfvffkVtUOb19youBUA/qeQTjpH21NuxugZ3cvIyqIh6xGsRT6ktF0yef/Let3vfX6iOa4g6G8QxjQieJsyhV2+m+tJuhMKYj+0ezG6eLHqRq/KNapJz23Bt5BiMQS1QGrqYfR0KpWe3pB8+7zA5W8XwwPvK4VH/10UBXGLIaxMcKfzx0rtffk0ojnv08wrlJ0xBTkCOQTAxsH8AlnBwfhk7iIhv7ON+fMuyLncIGAd10s7A5f62vr82JziaIw8Vbq6eyHolXVFwcmSQaL13eHCBnfTifvchdP7ICsUcafJr9DH/r3SWKtufDKfVkReVDK3XG/rBsgL70zkxGplXYoB8j43Vrlw6ptzr96pYOAvl1XCKyArCFYO2E/MipS/bEBhczVk2J8rQQSd1boCy58vfvtoVMiniUsxKcKCwOGKieNvEteoOBtO8Wm8gkiJI42yzC88eZ9KeAQPl0FVuJhRcG7RFSk1YKh5wNZPzSpJvsxl44pfMquA6iMv7vl6l8iKA7IWwdphmWSR1dKLfZEe5XzmoZ75InMSbrCwRqXPnsvBu4O11N2zqd47bpq6K3X3wI037y1csEmWaAoWki99esOPTR7Lrl34zL/6qdOR4efynM41p0rAyEbeu8uHh1mO5xXUSwry1uUq87mBZmBsSF3PjckyIiUgftlaotkfvGgh31ceE3lRkcuo1PDWqdlEujEu0D5STIkJuY36q8XpfG5+vHtILqIgflmTnuuBYosdvOPpg+0uo9rzerPK+NLSbG7fwYc3PD072nNI8SZmeoYXLm4EiROKn7En31t+ULEn7sv3l3C5x9qQdQj5skZEgYQ5jnUV7zT6KXMwB/2QNZwpfrC+m5EMMqlMvTy4aebY4lS+JDn0SVas716lxPuHuZVxtto7X9YqekPWKifrldK2toDbPJO1Cm1QJQZJe2U7f3ck0JFARwIdCbwwJdAhLF6Y7dqpVUcCHQl8FyXQCrzNAprND4tqFvIAp5wD6ABkYzMA4ArABcDGteYahkU4wBSACZugprsFJTa/9jeAFnM2ABcbBzY7XAdITf5cZ+QF5yyPdnDHtOy5BzB6yQIiWBCCsBmLDbRtb1aiHqadDZBMnmgLAk4BUAJysSE3bXV9XQZGDWS3TYkRI1yDTOIgOs8wbSuzXIhvyo2Y4N74JsfAcZM7smVDRLnQ+OWTTRdAIpswABAAUCMuqL+VhbyRvREQfEf+bGIBruIa4lYG2zDxaeeQEYfFgGj9ufxh16HJbMA65ab9zf0Fbc5zLQAzZbHymOUJGRq4yXcjloz0oF/RV2hPymKAtRE2bH7ZgAKSAFQOuoZUcP1M6Gbv4loS7ULfAJCjfc54aAyERJ9vXWvWFUayQRaQH+1gFii0D89B8858M/Ob9UsAayM/qDf92UAFZMS91I825jrqxHPpmwY68p3r6AOAjNwP8QaRA8BKecyKBvIqfawcFidr0eVSt6/kGgs7u91cozcxuXtzcu/6etIvVjOZMZco9ylGwpPSYBc4nFBgiCZY3ySB2oJs69QpB+WhrXl+O6DFxp7y0HbnorVNewIYxC1yIDlxgcZ8AWHBs2jHFaRTq5xVAYsmL1ygEA9h+UB7WMDizbVM+OlcPfhfGxtH3n843LC8bpyOBiRc/2cVmPZXNaKRf0nWDydy867++9t/sfbDJz7/hZdPfaNPrp/+xUSaYi4dF1Z2uYmhfneoe+1VqYHptatZVyimwtOSL3PdXYqnURwK5nyRFYxrgJptIiZednniyfdNyw09gYafCC8VQ3CU8rh94VZ1+qJb7x073uUtPqX812T9+YeqwY6TIi0UabcnlSgJB0z4BwRS+vlsqqJQJN31IMyqLeUYJsrpdG+lUk9XfX/STyX2BGEzwOh8yndHytX6SWlqzy1U642RgS76LHJ+i9I3WrJGQ5xyNueGXGLNWy8q/PRb+5KXuP3lz7paaNNEUxw/KQ3tXTt2HzHXH+RHH2CuhbRg3GyJt8sZvt+u3/5RaVrxKPZ841VXHzyycWRTI+FDaK5GVozpPBZGX1VC1oyxswFBzGGMu+bxkl7vLV2J6CuLjWZ9N6ERm/PdsYIfDYr0m92QjmZlYXF1yoXX9vrhpQoqcCThKYq7gsNotiiCGktEXQLWjkjsB3q9KycarlaruqlvRK50k+JZxItEJ2KMf0cJi1aAbfKkD79RiedQx1tOI2tkbNZj56IlfY7N96wum5Me8qM7S1fLc34kUyZ/o6waMrUw0yTrcF+0mMq7fL3sCO6cEv8WG2/Uk3HP/P7PlHBzBcF/lDgZLcGHsrqIPvjTejn+6XmXL7shc2DgrcOfXBNEqbfLndIrIFCIV0HcCtwqxcrCPPW/lLD4gjjBUu1sfbFZoDdds77xjacn6j1dmZpsJ3qq1XpaxGK5WK4Hi6V6sRGEG0SiyduYN6EMZQREyz9GbwAAIABJREFUQC/PDxrRbFCqz6nPHteray6XTVUVEyO+3mhaikgW1Y+96ydOFGqzT4nd3Edw7PZD1hVdGmc/pDnrZzR3nfV9Gbv/a/oOcSRl97B7Q/nowrf6X1y6b+CGI7OpvjWyuGiuHRUw/dpb1771KREoKwaE5ROLH3LejfR9fgN9jHc38RmWjqZLooZr1CuKQxEwzvOsbCIFi9F31h4rsBMuV+PNi5yoJlONYble6krnawvqZWXFu2CtP9m3bq4gawxP1hbzT9+5I6kYD18l+LZ+MxCfJ/NiYO7n/OnwGeYbU0g4W9PRDxXLxcuLLOmaPdp3VGUamTncxxo4HYbe7ky+Nrfp6qOXpHK1bDLTqOh3ysAaifnPLOdsXcda2MrFe8D2Eqyb+Y011iG5xspvv+HA5O67tt+9MNHN+pN5xtZwZjFy6iDSRRqLmWQ6GyZSqbGgWtqytKRsHswPrCNZO5+VyDybYDq/dyTQkUBHAh0JPH8k0CEsnj9t1SlpRwIdCXxvS4CVNZsJyAojAvgEOGSDAGgKIAS4ioY1wAugAJuDNylBCuByA40myAu039mcsqEhDzZU/A0Yi9sbgG4W8WwG2DzwnU0Ai3rATgPS28Ed+5sNBBuOJYB6UUq5lSMABYDfgMhoVRk4ZVrv9nyAnaa7BCXA0LiLojgZoZ+aB88xIM42KnyyMbMNOM8yKwIrO59xUoG87Fmcjwdg5TybScBb8kS2gOJcw8aLTR7PtOcZKWIkAuXj+ciVvP5eiXZjwxnXpENuVhfKQz7cRz7mtsi0+u13IxrIG7mRH99pb9ofEoh8OA/oSPua6ywACyNM4gCOkRic4zubONqe/kcfQebUI94PaEfKyLX0PwBRgEpcQU240tNrnOIdUujW/VbuVTeXreviH9xraCz9nAPZ0M4k2sG0Apta6EoQE8iTdqPfXaNEO0KmmOUJcjFXANSRvMjHNAK5zjayt+o75APuByBC+A5JuEUJgoJ+wTMhL7iPT9IOBdzuuneiGqZcI31J48h9V9a/8XghOTM843pKV2Tun/cVa3NL42j1sOurVL3ksYbz75dwGZ+0ZeUMrqD08/JBW1I3ZBUnnbgAeTC20Gyk/ZcPcwvVFnCb9qGO9HPmCA7a/QYl5gWsUOJjLJ5l87vKDGkBAfq7SmNK/yp+EaDimszRS/dVr3xC7kimDrsNyHD5+FLwOndV5tGP6gT96GNKt91TuPngje6O7Cc33rLhLze855paK5aF3XR7/+vcG6IvuLELh9y6TGmknbBI1+oHFO3aV2TcO9eVpqYu9Q8iYwAR6onWe0Vg7PuHFKOiTwHBMwquPSPi4mC4qQmATkRD4SuTd9096E/fdZn3FPPpXUozn5r+H8he8mn45Up9fnigsDuoN7rk2qkmLWzFLPHWZpKJoBx5i3IzkxcK5SWSrlhQBNZkylWSqeRe54XT0s4u6v6aSA6bS6wdX6L871Birv4/SoyFv7F6r8ncqNKF7mD5/yqq8bS+NzmprYkgfElGfqdqmdTj6Wr9Sp2jv/+GEm13toM55CNKtAv9+K5KNl16/KrtycObRoak/Q0YR/9f7cDCB4s+7qP/ngtAzLj+j0ofJkPFqfjFrTn3+OOLzXfaBuFLQ0L7FhQYpJAPo4s2Jold4Q8ohkWuXAsyJ8r1gZ60H2SicH7JRbnXELh8keTeI3AqTGe39A6nCkGlOv1gQ913ibBYPt6nb8R5eUCJ8f6dOpjfmIdpP1wlMR8xB692AC7focQ44/13LsTid6qcp+SDlYX73OyRk/V19Yvyj926MXNgs9wVXSYrADFvCSd3TNX+/vH7Nywe3ZpwjY2rkIMGrn9cmTP3Qjzx7kOLm3cVfYM584zWN/GCtQgg8r1AhOdbla4TQfCKQkKvJrU5dAFHW1l4JkQf1kakFQ1/NgEulmqN/p6cjHmiRfWj45VqXZN0kCmVFblXc2k65YeKSdOo18OutOIQJRV4u16PxnXtzkw2dUQmFjO1QBZVbc8VWdEEZm/56q2pxe5c9MBLLgmmB3oeDVIJiOHlI1OtDfTOLv5LAtwT0fscDogK3gMmW+bPxjcGX1H5dxd/OCuCl/EE0QiBxvuQNSHzH+u8f2qS7Byq97y5hH7GOKZT3qb0ekoOYRGINhVonk+mMrKUyNCfbe3CfMEczZhorv0E0mNREYmo6Bd5wfqLtQ7vHtprl/p8j5eIrpYFxhOXv/7psfG9Q/973/1bviwiASuyH27lh6LB21t5riZA5nKeey6EmLlvtfVJVrE0mD9l2+Z1ZXsqG3sHi0UFy+6TRcjw/ER3OddduSfXW5lWWel3vLsoC/sWWyOzpkBWdtjeg7UKCSWML4h0qCfTijJeTu8VKbKlVV7WYba2PN16ktBFEn3Q3ajXtoSBuvkzhAWyZo1DO52rQsdqMuyc60igI4GOBDoSeJ5JoENYPM8arFPcjgQ6EvjelEDLymIJ/F8CMQBWWaCzUGfzgtY7fwMishlgA8pmBY1GAG4W/Gi7snEFbLXNEPng5uOAEhsENq/kA6HBAaDO5oQ82VBx3wqSgrK1ruWD69DsZqMM2MmGvubKB/Kucoi/uZYyQFgY2M0GiWRkDMAqoBGABs+ivgBm7eQCz7Oy8L6JgxBGRnCvgev2TrJ7bGMTL3+cYGDzZEH4kAvAHCAfMrGyU4a46yYjBvik7qadjvwBgLmWPIgHgJyQNeXiNw77m/spn4H6VkbutWcbkGlygXzAXZMRRbQ97cEzbTOMaT4gIs/hPEe7XO1ZJi/kQP8iLzTmtygBfJNnuyyRH/kC0EEQsLmedMl+bUz9jGssGgnFNbQ3ZV2hEt4q0ykfLSsLZGpaguYCDbdO9HezpIB84PmUhb5LPQx455lGbiBjwCsIAfoc9eZ6+j7lBFyjbIA7aASSx82ta5AfwA79HM0/viMP86fMOcYV15HQoj96+4lq6tBCLRoRb7HT39Hww1Il7Zev3KEQB6PZ48eOp/tmF/xcUfEqqANpTKl8Nl/ruiZ+UG/KBSgISGoH+TFXWByLMwHItCuJegHiv6ftGVv0N8+BnGGcnumg7yNTyLK3KSFL5p1R3wtdX2ry6sVEplz2Ml/RuRVa539Tf7t7f+ov3Eb/yEUEn9XvFw94M6Io6utrXup9KiEA8IrjzbVb3YaBvfKzT7OuPEbGZ6K+2cXpnrmit/HI+OBodvYCOcZ7pXrhq5QX/QFQ5GbATtw/ZTRtKr6G/PMvdS0Bo25PeIFfD1LFk+HIp/9T9lePbfYPLXqvZY663sm9TRPsU5DdlNw/Lcjb+N65xermXC7dpbgKuWI96jvmZzKKW1JNi7DYmEvMBlFQloPuqZKfmPcrQUn3yS4gCvccnIp+9OXbIrlJYr6kD71IibH7ebmqWdB5wHXFm4j+TE3FXK/owy93w+kXuyOVf3RHK1+RdUjRBankzy125daXcpmviLD4T7qs3c1Tu5ggGwGSf0+J9wIWHk3Sct8F6+due+OL+c4cCBHOvLiChGplxruGsUb/IL9zOlrBt9GEbxIW6oBrbuzz1u4pRQ/Lndol+ns066LJHZnGzEjKJYZSXq4iUkgutPJ6DaXkCsoXtlxNJL2spCiXXPLy7vnVIJscEAG0LRtlFpNuaHw4edOThwM1dSSPUcueDpvzwm8qfUCJ8p8TMnymirXAdeYf5jkAMdxp/ZbSahYpX9T5P1TinWEu786F5Dkn2Z7LRW2Epd0SzAd9x9448Nf/KO9mm2VxdNliY2k85P3FjL+mnJnY0POpkcnGNblSdL2sAZh7Vzusn7xaP/6FEu945gTmI8D1OFi5agYteTKHAXQC6vM+u1jjdUapv2Wc0P4+A7yH2GMeb1rMnSN5tlwGrCzkGqomonFKllMlERNFjdFBERVqW2+uryeb13BOzs6WE40oLCt+RU8m5U3LB9wJWVbNeyIq5xYqgbm+ahEVjCPaesPA9PxCvlzpHT45WxchuH++t7CCsCh25QblU8pVhWvnyrLBeAZobZfTH+gEIDbj02J1NN3C9b6paT3BnM0z+YSgsHUfMiV2DdfwDlvR784hztGq7fX9frIVx4IXkc2HvK/6FfSZwM8uqJRdVOhlMMWte2kL1jmcox0qcoM0rSafEEBfTywRFvQd8kL5ACKCtUe3yIwbM4XqNRuvOHaHSI59u+7cMSwigbUWbQ5JeiaijnXUuc7VrCWYy1gH8l5eXouqjJVsoRp2Dy3uqJVSScXj8HO95XrXYGl6bdeJBxKJCLdXxJDB4tLqzbhkLWZuLyFOyJd1p1mNU+crVZ+HJvYPLhZnc+wJKAdzK3PImSwj+C0QZ12slhY21cuLsm5ZMb0zZsaU2D91CDsJoXN0JNCRQEcC3y8S6BAW3y8t3alnRwIdCXw3JGAbcTYd5rrCrAtssd7cuChhyQBwwCIccJB7AXXvUcLlBJsdgEY0aNlQsUgnDzYMbIgAVADvAKghRdgsACgA6BpYS57tGyA2EAA/bH64lo2SbN9L8y6qy+m1nFz7CUA37jPA3LTQuJb7KS/kCZvv1ykBcPB8nmtAqm2o4xtrIyAoJ9Yc1J+Nj7kJQi7xwzbwnIuTF0YsmPY+G3g2NIAI5GcxLXg2m8v4wT2U04ABazOrK/ezMWNjxHMMWI/HRCA/Iyr4Tn6m9UY5zR93XJPM6oIGNSC7ab5zH7Iwwony8h2ZADYa2WJyjMuXPHk2v0Gu0BdoUzaX7dYRVk8+yZuN9JIcw8YxF8wvuOoxI9zM0oQ+wjna/FwP6/v0ETb19GlkBzlAXQFdeC6bXPo1fRjgHmsWgAHakj7Od9qCv9m50qZmPcRGmHOUE1nTRjyLdqNduZ9xAwDJtUuk3FKsDH4jX56HnAF7AW4nswlX2lY6kH2kWnjKBUH/U9ltL/YSwSuHvJPzj7krj04muk/0ZU5kBOJzPeOXNiQP0xzU13M6bCfeDnYyphnLHDaeljNsAyvpB4yXTUoQnO2HgQsA22cEdrEMEdBIPWgHtPWJE0A/GoUYSCvMwNbs7pceqWx7or2mDRUT64b1UgaWBverA5dMinJYq3t6alHqFM3+rCtX13cfyGT6FlxBhIVpWcuqwl2885C75MkxT9Gsr80GNcWhqJ5IjIT5qKZxLQxQDjReqTIZGKTOVHcXJvYcfH3y9s2PNFbgh+5ouG6b3Fetf7R0+dFrEw9Hv/Opy+JjsSFvTonjE/NO4OZkI53Oj9eT3fXIDVai5Ma5MFHw/GRqwA9r84E3OhkmKvnQHe+r1hZ6/BDXMbXhfCH6iddcaO3HXIG8OfBfT7+sC9wPRVrsTZTn3hxkch/w/MxvNRtW8VA3597aTI8v/Bc3XX8sMznU+65qNvWuekpa8fUzNtcHlQWue5h/6dOMD7M2CFtkBX3iXUq8Q9DejYNt1k/u1hfGGKQlhNv5AO+QbU1XKWQ2mm4SI8ck4AEFqo8UiNvbkQqObMhq9NS9m6XTu359OuqWXxUvqQjL5XqYCKJEMp1KlDUxeAonoF6TWKe2yJYqjX3igg5V08XtiSj3sOIlQwLFjxv1B5q/jG1A9PPSxG/Liz+Zk+hTAHvECsEV12pkBXIGnLtYie/nbQWwyrPP+9QZXP9E+UffNilXUJ/J+7Vfzys+BIc89aG0/JKvv+6a+y/eefAvL3r60MeGJuY2q5l+ST8zB57u+En9QF9mHcP8fUQgPpZKs3INdYrMISpafcgsvOh/5P+KVR7AWLT3IWTF/1aCOEOu9Gnmo1NuU/5nlBcBuHUBfV1BtsPjqVRCEQPSPXL7NiDLi75qJcj4Sd8vFWvzUuGYyudSi7WGUzyasFKrN4IffvJXfVxf6eCdy/uU8cE8jNZ9b6ZSu/mah3Zd0D1f7LnvxpUGOBPDfdn5noLIiqrLVmvOk2O52PFpff9LJdZJkEDU8wtKaLLzrqbcdgPfmYvpa7yvmEtItAFl4p3J++dcgeszyqzzY1MCvL8hhmjUZau2qFF39WpJVhZlP5lB/CsO2rCp/JFIhuODm2f8vtF5LZ0jw1VYYzFHsoa7WcliQ5DRrIiLxZFtU6mDD2+cLc3kFH/F43eutSNufUletr40SwPm+FMK1VZG5mfWR1xnCje8clPzJ7tn67VkrwJjB5UF2cl5LiWXV1f1DBcOdQ0tyuIwMlKWLCESkRExfD6j9Hmln1BifcgYZ7JpTjiqxzrld/zwE+uqsh5hb4CVCX2Z9Tlr23ay0orc3AfIumKyVpzrVtDt1qXLNaIuZjl8Pu+qNpF0/uxIoCOBjgQ6Eni+SaBDWDzfWqxT3o4EOhL4XpdAHBhmk8CmBkCaTzabzLsGxALiAsQC7AEGsFEGXAWMWSISljam3BcHjnmGaf/ZNWxMTAOS3+MpLjPArl9UMq0x8uZZ2gjplnBxwvm9bNooL6AswBgH5aasfLKxIn989wMoGTgef6cYKMF1polG+Sjn15UAqgHC0TBnM4ZMIHMMXLN7eLadM9lSZ/LneZtb5QRsZdNkZYsTCrbBsU1bE9RoPdPKyb3IgTJSLqwfeI5p5vNp7pyMCOL5BpxbPcnPSIZ4XQzk4RkkCANkC/jA9WNKL1ViY0h/4TcjckwDGFmYDIy4QG7kQVkBsPm0/hEnLeL3sel9QglARKpsig1QO1lxk/9grpvoE0YkIRf6zDkdLSsL6kB9AfX4DmlBfvRzwFVkb8Qa4Ax1QVbIEtlwL2WgnHyyOTdSB3LC5I/rHXPNwIaW63km+fMsSAvyZqPMhhmACFnySVvyPIAy7iv/7dF6dEfywsxMurJuIdl9uVwNDcqTSD6dKe3dG20/4MLa8R43sV/uiNiEU27ubZwn2Ktbms8DqELDFvdNdlC3n1diLjiXTTljGHmhoYuM4gfjAQ1L5HHWvLAQEUgImcOzAbNfbpkRGLcvOSXrgMPvPVbbNFcNs8sk4Fi42f2X2s+738/+iuv3Zl4qNGSDXDXd+arEnU/d1njtZDUyHnApt3Si6o0VNrtLvWkn7Hq5vBsOT7gXPbR7yZ2KvMynukSFhI2fajzlfkpExZf9ze4NbfXDmmJMbbEoa44x/bYl/nvdpbD4+IGD4eY5pYcvld1F63cb77VqrZEMFVDh6ShV21fPZv1kQtr+bkNe2v90xslaUOpveLvW5xK75Hp/Pp90C33p5GytHtSmZktx0Jbxx5zB/LUjuXA8J3B3SQv0wz1NkreRH/jswRveuXfhhg/+51RqzbJbrcu6/o379vxvuYXe426ut8v1zhad3GGtpqFNe/43pX9QYpwaaEk/DmVZ4URW0Le3K71VCXD0Ne0ya/0N0Yy1DGQF/XCF+7HT3BM/vVgN3S8oRsWfcLKQaAbg3q5OlpVQQk060ajc7mzNuBPFICqKDde04M1pkk8FkZeoipGYK9a9XNofHEgmFgUoK9p5lBJxkVOc80Hf93tTme5ixht+JAgXXuRpmLbFsmDeYm7jvXG+ZW/Wo2UJwNxBW2BNx3sI8A1Cov1A1syXvBuYz2wOOwdRfVcvqaX9KuOd9/KK8aKoDu/aedmWbynGwtEbZp6spOrBH+kaLCqwhGCuXM3q4hKd/3irBn+lT+bQverbUyItlknaliwz+qT/MQboe/TB01lykCVDjDF0L3kqMZ8yL67K1p2NrCDDlvVPeHxiwa0Z7Jqr1gO/VpMCht6jik0x7if8VE86lc4p0LaCcNcTiYTcREULl+7/bG3T2N8n1s0/jkUD6wfevciPMjF3YlW2AzvVVI24G6sfT16+1W3bd8x1L5ScgnD/lK4C6IVgY4zSZ7BaQYZ8Z36grqvNzciWdxSEHHlwPeMaOVEfgOLTyuo0xeucPo0EWlYWyJU1Ke9kLBab1nr4BCSwArEUNIfFc+B9K2A/nOjfMDs+sm0ylemqEufIyE4jo7BCYF5hfcJahvFJH7taVhlrd9y4/57Hv3zJ3zZqCQhCSFMO+gvta4o3cTeMvFBNyYW1r61p22vHWGSehCyg71D45roJ3jioJQoLE115ERZOlh6HFicLkeJrdI9eNL5Z1eRdZoQJZaa8rC3ps/Q9CDzmRPolJAJlnVO+RysLmcTk2MBmBfo+2agnIMt5LvPL2cgVZFySz7bJoFq5MuYKyurFmIAkelbzfbtwOn93JNCRQEcCHQk8fyTQISyeP23VKWlHAh0JPH8kYOAwG3IW65AOgCN8WkwCNiNsBsxNDcAwmw9+N+sHNvWAJGym2KhwDRsJNM3Nbyx/2yKe5xmQHdfai0uOfPiNfMmfZ1FG5dMIXW38QpcUerb0TJ6zrNGs7wBl9jyArvcr2cY5/tz489q1e6kDmoKAb7yDPqr0FiUDOEwrjE1TnPzhu5EDlifXmFsngBf+RsZsbkyrjO+rbepMY4182XwBwlIH2gnZALKzQaKNrN3MpZEB7NSTvE2zk7/5TjnN2uRb+o6mqgExyN8sBiCEyNOIEGQJWGLaZGwQyf9MVis8z9w3AW4A0rNRZDO7moUH9aVsgDOUQzFuT2x2Xl3xWtM8n98BmpAByfKnbud0tEgLruU5Rk4gVw76De3OMygf11BfzrO5NiKNjb0RLsgHMB2Sx/oFsuFe/ra2pqz0L36zDfYBfacPkzdEIL/RniTrU/SnxNdOBuHexcagXBm9NvDlSyVZ9lKCV0Pf257wg6gvPTkp2ALQCKLRLG7OSgYsVXvFQTkpFwAW5eT5aHdzAG5sUQI8OaOqfet6ABasstBmtON+fflVpTGl87H+4HkAap9QwsqKPtK0ghhMnXTrM2PZdelD3ucn31OsRRlzYeb+uv5Od7G/2/3z9Medglxv7PXmbvmh1Bf/+vPBm39kRa31x0t7b09vyu53/f5UXX7fXT2j6BA6LpJ1Bb0hLPgukw9cakhFUc9BX9UbPJWs4B6RFVvy5eJ/3h7sy2/yD//4oWijjc/mY9VWaJFD2jz2wTuuD/6/m1Fubh6eXL803vGZ3Yq6nQsPennaoNsLvG2yEHiJrCkURdVzicifTYduYsD5heFEeGRHzk285vi9xcTiXPSjt7w3FHDbHF97Zw5M1vq3Yt0E0HVx9sTjjHfINA7A2/WJ0vTxTXf9+SsPHfvG4wdveFsut/5HenqS20XapNx1vf/ezZQfdMfkUKl78Q43MDkrh1TLXi+Yg5iPIQ0Z36ZlTX9m7gv++N80tdEZU8xZb1QCUNoE4GZHqHgGMYJIkYXl9kNjSkDwebvXeOkDofvQFu9Lrx7wvtydcG+4qc+78pc2u8JHx6ITjcjLbkw2DvQE1YQXpnvyLionnSyS/FStEUTd82HUF/jJhsJ/FDKJRDqR8roVP4C61JNJtbSn4AK+O570Nkw1vKsO1aOFv6pGJ36sLZYF/dLIVSN1l+t6ti8C1hlv9BVAR0xzABkvUrL+yjxo8xXZQe4wB31WiXbmnXA+4+psRfpO/W7vdciVdoJvrQKxXy3S4tDg1NyTlz4xRl9iDsI6hn57JnKB8v2YEh2N2Cz/D6TF2Na1yb071ntj9SBbTyXRTqc/Qvi8VqndstHqaO9Kno0lKXNX04r0PN3qrSozSAv90JBlU3MtpFgzRcW3qMuaJ9EII688O+3lk1GjVi3WF1x//fL7P+xdcfz/9qUaZeYAys78y3oAmUDYADgvH1g/bR47ocA2WffY1Vz6zLFvx3q5d0t8rmux/D9Gj0/RL+ljzD8QD7y/IEB4p57LvM57k+sAqyHI+WStRnlYrzG4WZ+dbp23omydP84qAcY8/RDCnrmgSz6hXFjXO0ruidK5LuctvariR1KEhdzbNY77yfApWSUwN7PWYA3H2oU1qa1/6FP0CdqNz6q+LfSvm0119Zcm5sa7ee8aYcH8ZApLcasLnm0uT83ShnHWvsbmOsYBfZryLK3zltaJTctNkQtjuuLKoJqSBUlqgy4vprJBpryQ3VHoL58UiXGXEkQu/c20DlgzMUbof7z/WbcxTzIfzyk/efeL6otThZzIChSZ7AXE3MIY4B21UoOBki4dorGD3cWZ8UQo68pVjq/qHG4r50QwPZs112p5ds51JNCRQEcCHQk8DyTQISyeB43UKWJHAh0JPC8lYFrgfLLQt406q3EDg9m4sMln0W9AOdc33SK07jNiAiDW3I5wzjYDtmHlPksI7HSLekAtwGGzRGCzA+hbd7P3LLihN/fKRZAwuoRZQ5APz+N9QRlMU4vNFe592Ihb3AZ7ptU1Dpjzm2lS/p1AbbS40apiU3+dkmmIIwd7N9lGzIB7ym0a9uTHpo1yPqTE5ok8zJacTT51ZMMWl4dpRiNjM/83cMVkiZsg8icvwGncOLFbNeKgleXyR7yc1gacoy64ZTG5sFkzmbC55TwbSOoEaIZ8uY/v/GZyMOLGZG8Ptr7CBhKNPuoP0KIN6HKMkni/MBIFmbOBrbkw8BS7JHSlg3VX2kU5qKfVh7Ihc/rMeR0t0oJnUycDACmnWZ9QR/qVWfiQP8/mdxsXbPLJgw0x7cymnr5q5Qd0BeyMu82KEx70CdOGJi9AR/KjfsjWyJtm3R6ebXg1KbdznTbeX+tPT1w8FwzcrJTcUBjL9iRmZxTEFtAJuVCv4FlYV5gcqTsEClruxIthbICAATK8qvX3YX1af7X74p/MHabRHD9vbkc4d86b+5ZrKOYYgEQAsl9WAiRz0tx2GzJjTrLIyJVTSfGTlwkLfv9I9dfcNv+AG/Im3e5oh/vb+lsBQk85ConFprVGKllNCaFu/j40OfdgtlK9LhvVXUIxhP2soHaNWj+uV7paZrPR9PCe8fLlPY/vfnfvZ3v+U/7f/nj7ZX312ZGbpu8e/sTG986KtCjvGn5tdPfomxKf/O33e1+curfv6MhrN8sV3pIrCz/9M37kOfWBptgE8ff5nkvPlxpdc161ODx/rPKy+z7gp6f3OQG2jG3aKtr8Fz+Y2Pcv798Vpruamrl+beGVUSJ1TCEkFCiDAAAgAElEQVR+kd0rleizU4kg+Jl1B/dLLfcz7r7XTrpLe35BcTyWpr3+nKbAqz7ujjZ+0dUf/5Jbd2RclhYNAPJvKDFGxpRM65q+F0rLPWqB7wiSee4VSq+X9K5W6q2H8vamrl4PU5XpYDib80uuOzE3ITdBXH9Ufz9b0D3zuZPRqAgLm1vdzf3ee//gUPS79TCalLuhasbzkgulqsQnqiIhWC+q5xS/oiGd5XK3iAlpImc0xmqe5wflusZioz6e7s72+H7UpbJvSkS9837YdTIZ9R+vunHcNMXd0mE58qdKv6WE5YlZFq7WS1aciwWERusYQI53wA+2ZGfXxskKXPkA0kMcQZia0sCKfM/FAuCshXvuFzB3sdbAwoKx237820bCf+Kem67cJcKCuYX5mDmIsco8wbvqTAeyeq/IvBOlfObjhzavyc8M9Iyma8HWIJm8SEOH9+hNSnTq02l+M/dSPuQKqQdxQsyKM81z5y2ZlrWFw31b4f6PN7rn9yerya5EcnosWZjdm8nUZsOoWg67q+O8WygzfQAZUAfIWvrHKQexKbCyWHd08hTCgosVi6Y2NdTjK9bFmKzFeOcwzzfJ9dVcacUfkF05Y/J+Zu2BGx7mFUB05Er7IsPblVj3MF+fN2l33gJ9gd/QsrIAVL9TiXXQT2BVQfDteqXkGgLR5SXQpEBfZU2j8ePtVvyHyWoxvVvExZHCQOkanedC1ky0E3M36xYIOsYEY8yIxWIiFa7ZdPWRh3Z944JdsnrYrveQpk7Rsw2fuZ53LH2o+Q6OHeSzPPeepmmYC1gXMccz37crr9Dv96uK1FVrJk8esPzazOH+nnxPpZzvL3WJsICcZT1l63nmRVu3UE/yp/+R95jK/FgUeutFWOjVl4C0jx+QOFhTQQK214frJurl0rfqpYVbVgn/gi+425SQ+XkT7KeRT+d0RwIdCXQk0JHA80QCHcLiedJQnWJ2JNCRwPNSAgYWmvm/aeYbcMrmc8nZ9DMuEsxdDBtWc5tgrgP424iQZYG0BdU+m6AMBAZ8YCPFJ8CnvDnfF7jFXUWXv/iEsDqeY9qFbJB4Nhsx09Ri47JZCW1K87u/GjhqIDvgCOAsoOw6bQbJky06bpBepmQgMCCgWZ6YvIy8MVdD/E25ARfQJkWGaLNxjk0UJIq53GGDyKbMyAKTKXlRXtN2pG5GgnAODbetSrQH5aacRnDESYk4SUS5eA7y5Dt1BlignsidcpBH/N1LHakHwIQRE/p6ytHUGG2djW8+KTegPJtAXAAgO8gkA4xM/lZvPtHMhITZ6cJy3jWKCVd83IgFs2KJu9ei7Od9tPql/DNHZpVDmag7ZTBSDlm1W5GYZQXXIE+ABGt7xg4ApaEH5G3jizIaqce9XGNys/utvZpjSmVsgrYqoyfCguv7pH3O8y/pF7AurfS54dSJEwkv2KvEeICkgwybfY4gG+UifZNnKcXVdX9dfwMU/Aclxmg7sGzEGWMQDX6A6viBTAFM0Bg9ZyCw5TceuSBDgHK0z5v9XjIZwsqiHqXd5uze/pnFdsVP536n+iHFu6i5YlRwB8NNcYC5WTbJ0fWnFN/dqy/HrsjVqt8aLU7vHF8/sH8gXOhJDzauVasN+6dmv6KCjZ1qsxmn+N7hb6w7esRtHd2/p+uiYmMxIQdFsWM21fd7O7suvfHquUcfeqjv2i9cOvPN2huL+5LHsmu6fqJ0qFdkRv6z6380/Fbf9ch8yTxKPUTAerOM3Y3Kl/Kuete7D/357PvG/qQnXTpG/6P/QgoyR0wkSlOXZsefHCxtxKsQTELPq9WhkBvuYGys/zhgp4Jqu/UiI6669y734MvKblv+XW5tBn5q6chf8wduovd/lvO3/97T/RMTd0stHFAXzVIDJWsQFVyr9qKuzCeAmWi0MhfTH5LVMOdmgwGRFRk+w6n6iFw3yfub83cfrW7ePZI6Fuoa9aPzil3hFEelCYSNld3g7lL07Wu7vWaluxJNkHejXD49kQzq49m0X8inUzOVWrAoomIuqQAncuyk6siGwpOH/0bYqAVhPao36qlMajCdzdWTCpbMgFRAAYWQSVW60tt2F8OnXClMQBi8b1lIS18QGmTFLqUmYbFa3IPYPfG5k3cMFgGA1My97ePHblMvc/9VCbKCZzDP2ru4rTjfE38ayQ5h+SmlW1Yp1bCsAHpllTPzc//173hX0Ld4T0GOMee8X+lfn642IjyYND8oS4MPjozPPHp0w9DD+WLlulo6OSgrC+YcAzdPl8WX9MMHlXgHMZaqz4H0XfEMs3jSyaW1yod7bO5jnALwmqUjpDPvFcYw1zCvn0J2rlIB+kFTC35qaHUDkpmB7o33vfSygcev3D757r+8vWhj9Vx6B/FJYnGKKFfcqnCL/obUxioTOaPpzvzP+4F5vqx7TeFixePOEPfkXIr1/XQN71kINJQgSOshLBqysggVUwFrCy+hSdTzjohoZR7oUoDpnrkTPQnFbXhF12Dx4Jb+w7iFYr3E+smsaVmjjimxdjBrUdotp2v9NRdMbElmgiePP72GTjVcK6eOLk52Pai8tzeCxIBm+3ZrqfNpk8/p4ncpxd+LjA/mQNa10yrDD4o8zstKRAue6FAi3ZAnrJB+jrUJJJlZaLAuoF6s++lr1IXEWruhPCg/6y5kyN4Gwo15lv2BEQ3I9RTCIgyC2yuLsxvEEInYOGUbwTxFHp24LefT8p1rOxLoSKAjgReIBDqExQukITvV6EigI4F/egm0+bi1AjVX3wJEbfPM4j8OOBsYaWC1AcumCc7t8XtX5Pssag04OqbEpoNNABsnnlV2jbJi5kqpa+7ejBtcVvdjM8J1AJC8MwB12UDwnbqY2yADnVcjLTgHaPByJTbhAGv8jZY9IDvy4G/yJB82PuYGC/lwD+fQOGPjA0jHJwASsgGwM0KFcxAN5sYJdyoAMXGrDa4lryY+2Xo+ZbSNFvfwG0A5QBwbUOpvQLq+LpNJZo3A/aaBxqbtiBJkBcAl3ylTnHBputtplYPP1eRGGeLEg5FY8ev5HcCFTWC8nMiPtoq/5ykrZUCWgB2DrrIn7apHp93JvwXEQSbmioDvnBtTos886wNri9bNDY0DI4rMmqSdiGknZWyja/IxsN42r5y3uB08Jm6FYi6u7B6T2ynADuQKYKzcDKX1VcrC4ZWlsOBdWXjg0VxCHtDDVD3jV8z9mFlMnZdMVgGkLH4HQBgHY8nIP9ykoYVMO3FdnHigzek/ACCAf/Hj/+qP+5TI09xenVc5W8/ElcmftfLB132TaBhOHXcv7rnDnahtKCvlJC+FTPabY2BvuKpS8vKzX9H3jwrQfNRlvKWmy0T1b/Z5xbHRvlkp15e+md4Q9fnZVQOIryg/ZEUzioh6BiYxWbmpv3z6iYG3Hftc8MmN7z1Fs3tfYdvb5lK9O9JhbUPRz41216fclkbx6LHs2nX39b24f19+G8Bl84izjwO1mT03Td9THa0edz+z5w+u6q3PoZEPkUMFPqLEvHPEr5cG+x/8+MVGWCQXT74YcmK1ww8j17VQdpc9tteNnJhyX3h7XVYre93FhZ9Zvjy3/V/kjg3ftGbq8T99fOiRv3lscHKu6R5GIPMSUfFvmn2csc24J71diTlxi6wTkg3xbcerG9x0MOJyCr58sr42yPuL8tcRPJ32GvcermxtPFm8Ji3Dkaz6fFX98lxc1DTLp2sZJ/Va5JK/dzBK/PHF3uG+ZNNNlXt1vxd9ZSrcP1AvF2uNlNefSixWa8FxBUDeL3dP6/USHJDViBcE0XwmmezWQ5MCv5vu3Ir1cDDVCObz6WRNGKHqEnX7YXeYaAxNJP3CZxtRuZ2w4JEAeRB+9Pl407WL3uRlwDWgL3Lj3QPRs9rxDzoJGcL7EUB//jsFrJ/med+p08iBORZXcasd5uJxSP2p6RJMQL9ZqTFfYl0FAM764L1KI7hHi2Qro0gkbq6vy5XyWVn/BE7g/FVBKrmj2JXDJZS9B+1ztWejvf4flXi/soaon49MVc7V2pXnmUIF7UsdeHcxpqkrifGDhjeu0pjXcPEFmQgZxdpiVR80q1TgSxrXT6eCRtoPwxs1lm+Qu0CA3+Uj9P0baxl/vJZJPSz57nF/+nfnPLZWeZ6tI3jvmKY7IDIWRqw1eN9TD+oNsdm05FBaMfkYCdIhLlaR8MpTyM1IIt6h71i2sigXhaVHsrJI+lorPJrMFrL6LEjSpeJ0YbMswxR7JxqQhcGYl2iu9enf2AjS/vQ9xhNr0zuUIAPol/RdgP7tg5um8/3r5hZlmRAqdVeK6b7ZY72fPfLEupdVF9NvYEXyLA+zHOJ2ymQuNelPr9Fa57ieH3UNFZtBw0WenMx2V9bo/KCeWdUn63/KzhiCsGDdAVnGmMNKmvUK9VxLPpLHYd1n7m/NvSnP5n2F8tApfrX4URYs3XIFpXquWkuIFd67sx13UM+yF3Ru60igI4GOBJ7HEugQFs/jxusUvSOBjgSePxJos4JYdVnO5oi1e6xWTWD1NETIeVc+ur2pVQWQCfBmQYcB39iEsJnqdfs/fMTt+C+A67gbYONvLgjM/BuSwUzVAfNt4xWvk+2ujIShrGxwyANwi3qhUc5Gh2cbiMIGHDCdsrERYvPNRomNO98pI0ATGyfAXTZfaIFzH5sqrmlqACttUUJ7FNN18jCywwAV0xqjftzHJosyIiMsIXBTRV78hksSc6MVJxAMHI/XF+CQv9GGBFaFSCCmBKAzeuP8xrvXTPUNiI7vSOP5xuUat5Iw2VI3ykR+yMxcV5lFSfx+IyWQI8ceVz58mZu4FfIAuXMeOSFf5EK+bK4fp+94r21ueJ/TESMvyMf6+urb1NaTWuPifHbsK/I7j/GjsRamREzIX4h/stQobFDo50MC6mfWZI8WZG2BVjBuEnBhcsYyn6OQkDF9lw05WuTImk0+4wrNRrTXaU/AKLPEou8wBhnDEBZY5sQPwCsj755tGbmPtr5DCQCHPvweLA7kEssNp8fdO0f+LPfNuVcLDF/nH66A+575gKxYmzmkgjWaxMdIMFvsDktbN9Qm09uC41szfv3HfEI2n+FAb7UhSUQqWWQzgm5JqutfvPj04C/t+333yqlvuJ+++k9OyeXPNr3v8tdMfPXyhWSX6wpK7nBug7u//wb3qY23uOnUqR4qPvb4L8xsKh8sX7qw8zd6grn12QbDbPn4tr4xr3Aw7zjFrXDpqT0uNXdkIT25ewWI2boOd0JYgTUDaidlaiDQ82QUVnvHq/dk5uq73OXdH5AVBFi66tRz2brKSz/8p09d8ca3dO2/Y9cNP/RHkYgKDmtbxjrAEYmx8U6RFWsqYd6N19a5o9UtbiYYcurLfP+62q13TfroAzr39Zlg+MpamKH8gECQFjMQEWcUfutHXcvzm273Ttac2IUmqdskLH5gyLvy/nnvE0kvU/PDeqlYri0odsCMn/CK+j4rIqJLDJcryzV8KHdgGpcJPwySizVRGop+rAoteNX6XC1oTEblaD6fSzcybvNsFN6ni5vkXbsWPFZiEHu8q5i76LPt9aC8JBoZRg2SiXcHRN9qrkmoCu+fv1BiDNLTVsv3XMT1T3UN9cPtEu+032orBJZEvDf/viWzsqwAmooHIgSYjxjvXzu8aSQxPDH3tUTQeIsCdv/z6YEep0+nuBVuoTun4PCLTSuDci6Tk9VFc26GjBOAf0qdRVJBnjyk327rn16YHZ6YTW4aG29c+qGjzbZqWUbEieb2tQTvobh1nhH/fLIeYA1hxIUpYEBY8B4H3Ad8Zl7lPfxjSr8bK+TZHM/ZpV/UF4irrKyknk5XgwMavzOhnzglTo+uYXywhjoiq5/ic3hXIAdbp+FOhzmf9wAKEPRNxjDzPWsg1nVMoLy7ec+f03iOyeH7/itg+LU33YLsmE/oT+8woVSL8wLV665raG0+CsPXi3yd0gR2gcD5qXo1+aRiP7h0vrZFf9P/GE9YwbDeo9/Rxw4rMZe8s5Un7cQ1TUUgcYGhXDAllMSMuCDbU7kp31u+p3d0/luP/sNl/yuoJf+ZrmMMnM2CabV2ZI42ZRSbD7lO84On+GXRXDpXq8vKo680lwvk1mpe821WtEtCIYVYb9CXcFHFmp31LWsSCA/mGVO6OFSvJL89e7x3raxNWDuvZkmxKlmh9V3N8/0rZMmSeUava7kan9E35jKzpF2tfp1zHQl0JNCRQEcCL2AJdAiLF3DjdqrWkUBHAs8vCZyna6dnUznmfNNGZRPFBuKQEmA1G5mSKz6x6Ga+dqfrf3VBcSzYdLDhYlMFOMAGjA0T6B0bZdOSpyxsasjDNsoGQJgLDQB08mGTw2YHZA5AhXvQIDRXSQC4XMt5NubcAyBhlhc8mzwABc1SANDCNGwtyCBlxdUUpAUWApTbwHyuNQsR6gVgDDhMnvuUyI8y8Rw2lQDVaJ2SnwHCRhgYQmNoazMQbisvgGWABeqDrOIWGvHNm+VlsrNPIyh4BvkbyRF/Nr8hOwN14mQH15v2KfeYlibf75Kj5PXOz5xw07cB9vEsI4noE8jM3GEBbv2TrRdahMN3A4BpjKSO78snFi/rSc4erYZZb7Y+VHti8brwyq5vPT2QnDjovHDuObqCkiiXD4At+hvthNaxufSxCwDDtiiZpQtjCeCBvsrnErq98gB0pD0B156rzBhrWB39lRJEzUcSXsPlfeG3yci9UiTErZMoYZ/5uGX0v7kt2d0qjO+yftm9bvEh1x2WC4moURhoLBRzYfWMZFRUdPeFx9xjChNd1/daVHUfaMIXMX5D1hNuoD7tRqon3cumv+nuHcCw6ZmjmCi491z7l+5N41903cGCfHmAC/luJtXXck8FHbN0DNUm3Y7i7v4XzT3SBLRTYbDswqp1iZEVyw9Izh9xuSMPuihd6Hay04l8YexygtQ6AKfMcoZTOwV4jXth9ET3Qik331N4XyWc8B9b+F13SeFnXV8KvkrP9Xsu6O9+1V+4q27+oYcP/4fxO6d/kjHK/EbbM3cCym5RegdkRRCl3HzQ13TLhSWLAqMrkqlChAf9KREUlcPVbd2Lje5rRMZpTvXeqvuYVyFSHhMRQRltDl0hO/sjpqHNXPBUpeEu/8ZsdPKdI15THiNpd9GbhrzEhr3jwclqutrbnT3Zlc8AZ4vs8yu5fFIxLJyXaoS5mhdV1HxDdWkO4yBM7Vmbbrh1MtJQgG6vogDJ9XrQqPh+f9Xzs8cEqt2vR6zmtucndR4yGcIPYi9uxSbyZn1SMVN6037t7cIEX6ffIfkOKJ2OrKAqMF7MgQDt5H1mJm1Vaf2TnqS8vLOYC+JWW1aoX2jVa48A9SMA6sT2+OPY+7uwWO6V37fF9YdP/ndFSH9MLp9+S4TEULGQcVODvS5blpscrC6kb26ZrkZW9MwXpy958uCeTQfH761mUnflytW8LIzWp2v1LhEVzFGmYGAUJH3Q1hVmtWmWMawF6P+8Y7metqFNAVI/rwRJgHIB5BbriF9RwgLhlufQGvQv5l/IZEDnJ0Q4luRWi/GMbCEUsBxtkpE6WDP9aOs8Y4u+9lysLJAH7TimhBx4Dn2XNQXf+TSrEsqJVRCEqrkdfQ5V/768lXcefYe1G/1zIGxoSlE3TyiGRaNRd+lsF/K3+aNfVhW+gP6Tx3ePPJnpqjb61s6PKGoP/cVckTLPmotK2oz+YG6ObE3NnMqcPqERUdLbKJkp1N4gq4U7uwZL++dOdB8lzpJ+P991GO8M6sR6k/zpF7w/WuM2KqUyQSPXU1lIpoOs3FCtr5bS9Vx3pe4nI/o1+wSuJ84Wz2dsmrIPLtYgd47pzXF/UE32yZ2VxKWX/BKBhsIOz6YPM0ZXPeR2q6LYFcWwvkIpwK7lWVta+T3f5uHTVblzviOBjgQ6EuhI4DwkcL4vvvPIunNpRwIdCXQk0JHA95IEpCE/I015Nk+AMWy+2ZSZxixAAJuZPlfZl3JRIE2xBGQFoA0afLwvzFUTwD4bFwBwQFfTwrINRdwtRDsYCaCEFhrgAxshs3ywe8kTIIL7KBMbLTZAaHjxG/ezcSdZHUzrjHO2OTNXQ2j/Ul4D/fm08rHZZzMFQninEuQErkDQZuM6ysizAcIAPtjwWX3i5ALn4snKe63OQ4aggm6BtK0cOrWsLRcvm5ER/B7/zsYtbt1h9aMulCtOGJGfkRWcN7dXlIs602aSS7DP7ft1/mZzTX7Im9+WyKsl0Iu+MkjfoUAv8MOTRnpvsdF95UR99KUS4ojc64wpbsOu+aA/KoeF8a7E3HMBn9rFR9sAMrGxJ1/Ai7iLGtoAvXr68B+02ogxiGY5bUbbxQ/yArgFKFvyu/TcDsoHeMPYgFghZsAXfXn4yngVgfK+25rd5Y5UtypQdXtRlh48mj7i+pOT6lChK4ht2Fg/7gKpbYqkcF1h2WXD+pn9SEXuNi/r/kAxLRbFSQyq1ruiwyJdA/eLyp5xjQY1x34REWu3l/blfnPXh91vXPLb7oG+62VNsegWZVXBURLG+DfrlhRc11TH3XjmGeXq+CR1zdy3Xd3LuKRMAqAxks0QLGc+EtVFlz/ygGSScJkJYYbLHgCb9zHn/q0S44lx9AWBvworXSxlKvX+ZL4xHyQT762F80NPLv6RG83c5Lbn39O80fdS14VR7RMTtW/hEIfxebMScxH9YNm3OS5D1G+b1ityZeaKYZdbCPqeUrDtlFw/JUVmzNajVEUEhlmbMa8yXwK8AUZByDIvN60nzlBb5hrSSU0Yh249GRVEWDQv35BxV7912HM/cMP10e986oH65nV9i4pLMRmG0d5UMpGVMBVQ1uXqQZhw9brikqe8soK+FqsNubEK0+lUUi7BUmtG0tHTUT04Wq+Hesf0KjDt2ppLj+GLnfp/ZJWyvVnn6IAWXwaQeFqEY1oB4neImHpjPUy/TC6xrpaVFG1xmdoVUo/84gfupSDnkAUEIprJq6JoZ5BPPA6BXWbdy8jk+O3Lsn6uLnvigb9FQDBuqQOa+UbGx5+LzO5RKupa5hn6Au8/3hvTcvO0qZLLDE6M9PFeWCurgp2ylMglwrBf7bh9347VuNKVUrn0yTEnd2YDIiteWlisXCGLhF8W2I+M0ZqGaOBZyBq5MDZ4vzMHUm7GthEVgJ8QAYC9NyltVkIRgP7KexVy/WeVGBMczJntbbuycKf/6zb9BDlG/+D5lJd1Ec8ZUwJ4rj59yeaa3D/x99da5yi7gbvkzhqCeyECz/nd2eY20EpJHwHgZi1Gu1IGLIWQCXJgruc7fRvShvKyNuJaA4wtr87nGSTQsrKgX3Esk8yQFvVa2YWKryNfhk0Co3Usrb/kCmn6cH+hVkoXr3zjU/tlHYGlEvORjXn6Bv2WubPpDk3JCAgjL8iSNTcH4+JKuZlK5nrKD8+Nd8/rGVx/vgfKLIwp5kdTmGG8s+6mH82msvWpbHc1J9KiR+TFdpEtE3IFdVKJdQfk4Fir3DyfepAoM2OW90i3CPNLq8XMfeN7h4m58W6dQ3aMW57D8049ouiwfEiVZFmRK81Oano4hY9gj8HzsVae6biDOt+m71zfkUBHAh0JvDAk0CEsXhjt2KlFRwIdCXQkcK4SQGuMTe6jSmg94WYAYIaNB5uMjBv/Pwtu6IdH3egtO/U3oBgbB9O+NzCeDTybIQPVQfXYvMUBfdus2TlACDZsbGDYsFEWNoeAZmxs2OBwDUEK2ezxjjINTMAINNbYZHEdYIJZDBiQT1kMOTVrDzaAnGc3ZFYVBvbrVLMOADVoCVMHNvicY0PGvXwHVAUEQEYAIUZOcD+HaSYDwJgPacqJnB9onYvLwgiTuMWFkRb2W5ys4Blx65X/n733ANPkOut8T1V9qXP3dE8eST0KlmTJChYOkoMcMMkBTFxYm7CwcEney+UuGBazd7G5l4VngWV5YC8YDCY4ADYGBzlIVjCWbdmWZMkKo9FMT06dw5cq3f+v+ntbNT3d092aEXc9U/U8p7+v66s6dc573vOeOv//ed/Db9xLWyA/JpJGUhh5ZGXkGqsPQLaFeWq4g79ddnNfRY5MaKk319Iu6AT1QEfIh3a64I/ndT8SiJi4VsSEiIpSovBFsciKfm02XdaEfFor1ad+7YV/ca5eC8vliJwNXATUpn0I8zSmBDBAe4Kys3klYUm4lj4JeEefyR+f0D/EaKd/rY2yr69FqS+6T3kgr/5QYO/Plf224kXE7iXaz6K/NKONquVVIBV9cO5WfS+5b970Ea32H3Cs+u/R/glb0kl3WXjcbYsmnLwqXH9SdxV5LkBkLDsA3kBDIV6elvbtU8YPSIMTERfl5LBuaGU6/xklbAJgBl4g/yCPjS3bm8fetbV54jW/8cSvu+990d8vkRXLH5InK/jNGvWKhafdy+Sh8byFJ9UQsfYgXXNRJ/K+yYnU6D7wL66x42Z5VrS0tbRHPQBbIFoBD/+8U0762SIpkLr2Qk/tmAKBdPaIUSwQkTpHW3e5rmCr21Fd5GJ8r/K6/tJVX6j5m++QJwZx+LEtAJPZId2U60lVoZ8ucwLp3Vw8GB5sXn7PdDTiS38TeVo8rXZoyLMCjzVAT1bGUmWeC7CGbcFuYids9exykQHEo5vo5KgStiI41nZj2qT8ZOAtbka8uZzp5YFfe8siaXHp9oFZeUsc7K6VkyDwtcGrm41d0ut7aSDCa3K6lWzVAzc1S9V2IwhOtpy/UE/8qcvK/v6Ki4/VG2F4ct+ro94X3E8/wVuOsYG+kD/Q959WeqXS+xVsC9JRWdc2KRTWWxQG63p9vwpdGyhNOnlcoLt5Ut3yguhARkZYmC0/QxYrnchtmMzPRowzZphs6a/0JZSKhB6gI+aFeM62BU8J2kWJ+rH6mfF0tPNpHnqUj3jy7CfxJ0roJzKknOgV3xsK9dSjxHh9gzws6GsDir7KWbsAACAASURBVJkH6LrqQaio7ccm3dDkrBs5NaM07bRB9xahkVs6+7rwzpF3ywLM5xnmJWh558vKOfPCXO3ZRlbw+7MhKyBv/o9OWVhowPN5/4EEps14H0DnEzbS/v2f70NGjIvoI7+/VIm+kX/2r+r/z6tNGiKTKP+6jlWIK/aO4TnYOsgUEuM29gUbiJ4RHg4do1yQF3jFASpjL4pj/RIwz1IIesIboZuZxWw35rWPRaBUGQ/K1ba8P2lvxuTXydOi1Vqo/GXYLDfT/uYtAvyN1VseIpD+SdsZBrNSCMFukdAfkceCwPyuqp49puvpm/aOnefY16pZ3ruPPm7vyBW8NhTKaVLJ12ha9cuxJ9JiXNaLd35sOuMb78e8A6NT2Cr6Ae+SkMjYe0Vy8iYXJrs97b/x4kpXWJEc7u7su2Gh2ZaXcSFJ4jltZt5YmDxxddQ6Y30Fz2eRBgt+qDv9sTgKCRQSKCRQSOAilEBBWFyEjV5UuZBAIYGLWgJMAAAJmPyygoqJLgApoQQA2Jn8zrjpewdFWDBRYwXhdysBKmSrC5WYXXAf/wN4G4COYFdaRWrnuI58yIOJD5MSJkOsqCQ/EkAA5ch7DgDssFLRVgVDXOQBoeXEiBEIFlLCwH7zOrDrzTOD/KkHE7mfUgLEQ0YQKYBkTNy4hvIyQTVvBupr5Iflxb2AGExIARW+XYkJo000l4NSy//P18V+y5MXVhdkT/swIeRApkZW8L/FO+YaZMp9tDefyPsP3NO/DviJTMaUAJIApFm5CclCff9MieXpAFoX9AHQ1zf/u71/O/8j6ZF45wmtxN4rkPO6/mB6TkDv8T2N6w/eOfWmuPah/5zJ4dmuhl5lBS1tgH4Tax2yiNjZEIJ5UML2K1itHdC1v1JCL+ifp+nVesqbX6G97CHk1ZCM0J0/VNor0uLHtWL9BX0iK67veUCr+sFcUi3FPqjNnjcr9FPdlctt7QJ9uP3m+qcqiWoCUdEjr4qywH32JX0mCNPS0yBkPqAEUMgzsRHaKUEODyXtb3CF/L4eWOr379VvgJQG9tI3p0Va/GIrqO7c1J78kR87+J4X/dmlP74z9Mtp5JWwO2c9tA+G+5n9f5QRFsPtyRxZcZooaacDnTLSr1iNDbNwTVAfn9AG3KeC5qxuSOlL9CM8U+hL9DmALTtShcdJ6z012urTStiVLLa+oiG5ffUPCjE+KU8LQu7LMPlD23d3f++P7Vl4jwihDPvEfi+6jvAAEUOTIfyqgo/7jaMiMCrtpNLUp8id9A7J+pSIDQB59APQGUIYwvdVSgCbAKHoIfYE24c8sWlWeXQR+4ItQ+78vr8eu+NKv9xXcu+hHCIkfuLBQ7P33nxJP89JDx6baW4f6Z2I5UJRrfgzge8mgyAYSVzaDLWnxYyAv3Ip2Vkql/rmw/TE0YabrnteNOsl09tc2BrSBiWQH9I9QFhk/bNKv6OELWPs4MjIEh14iryTLyKbxifDLfepCG+UB1BJJE62AfluhSYreZGTp1QZwq1zoHPYf8ZGCB1s+IbICsuo80k/we4yTjGW0TkoK4Afuk0DMtZkxIASJMmEAGl75oos2Vp9uENW0E6A1thxA0w/qu8/p7R8zgcwDxnKeIWuMmZQZj7RA/QEu/ICERXkxfi76iFPCnfDQ3vdoHB1eQ6xR4sLtFfLahvQdzJaLTTX8rIugsbnfqCX2AJkTRipzynR9ox/1JFwSox3XAdZsYSkZkTFw29m03sO2ghSkn47qrQSqY9nJeRaU/cdevvT7zGFW5GYWqt9lQ/32YKNL+k7ADaA+quVjKjivYPnQlTQxzO72CnvORNiWc0v/APdoD/gbYXOQ+6Ju9a4pb13SpUuERZl5GwHoRw5HhBZ8YaDD+588ppX7T0ozwXGcxbCMJbnD+xD3kXJ3h3z1+CpMKoT/UElnhT4zxiBJzB277xiN2Gzcv3k4aGjXf2ttNIdNpNYbG7gDcgKYLduU2JgwWYxpqF39Fn0Hm9Q7AV6/ZLBnTOvbS5Uy+16eWHi4KZ6c66KHlJXxhM+GW+yQ/uAnGrX5x6dP3Xk9jgMYTyWiSjz/qL/MWbZ+/zya4r/CwkUEigkUEjgIpDAeR30LgJ5FVUsJFBIoJDAN7oEbMLLJAOg4hVKgGqMBwBqTILn3OQ997skGtLMjIkJAB2gEBMVJihMPJggAyIwIQY4W05UGMhu4H4GeioB3nG/ERZMpgFImAwxuWdyw2pG8mQWA6jD74A9RmhQVvO+4Fwe2LfnWXnyK9I4ZzMjIzwoh+XHb9SRzzEl9vtg1SSTf1YjG/FgK2TzzzIiAaDHwqow8eUe5JT3kMgD0fadcpjHBfcDSFqsequLXcP/FioL4Iv/+czLwa414odPyCjq+oR79Ifu1SehQgCtmJjS9vyGLiB7gX1ZOyD/C36F5nfMfsmvpFHfQG1h/K9bbxlr+eX+/e0rWwoNdVJeF/5cPLBWqByJaX3HCsBUBs4LsGSCTp+0PVVWypCVjXi+ADRyMLGnzWh/QBTuP4OwWF/Jzn4Ve3cIeMMWQCygS28XEH5Dd7DQ3yWCQmo4M1SaqGxLDz/s2pX3amPt6d3p4cZINKN1/62XKbTS8wVeXh24hFWZgDnoKH3kfyqxUtj0HICHOkAWooOAJWn7/UvABf2P/kGyfox+o6dPdsf1p7e0Tz30U2N/csMLp79a+eSWb9t8z8gr/+Px6jYAvBWPl0594YlbJ++/o+XX7tjcPrmzlBKqKsUW0RYAyvYsiEGAcfqIgZ+E3bmztHBqX3n64NGkXFN/8mlLgG9rC9o4W519WgHe/eGYfQR0DlAZcOsH+B1S4kjzM4SEcru7Fpt6S+WlujlxkBYKE7VEVkD84D1Q9Vvjh1q7H1EIqMnxcGsqLwN09kH9/rUoLeGVRtmxMfR9wCTkzDW2wn1U3yFfKDdALp4s+b6PrLGFPJt78NRo/8re9PgfXrNoxvSX8sPqPdnxsnDHxudbozsHJ/RbW8Cb9rFIZ8QVjFfjSCvv/UsPK+Z5I/QuX0j8NIyT/ceFdc95Xnyzi1r/2xufl9lr6V4oOfFs9AVPordnD1w8jLjIvE2Qh+o7ov0rXqTwWKWKwpeVvVYmJU/hzAhhtrl8bGq4fGJBpMWdup+V1By0wZjShsNA5cqCHi56Ki7aU4Bw5Ig+QCIgKOwtZADPgtBAL9F1dAzZmxdGLtszvwKe5w7ytXY00BpiiXZH5wAaAR+XH4RmggxlnOPZ6AerqUmEnmO8X/VQfz5W1SbU249OjFz/tX07RFYMd9Wb2QbcHGuQFWfL2jytziqDDfxIP0bGjGvUDYMFKE3b0B7oO+8l1B85YHPyhN1Kj6Jv0FbYqL9Xes3yi6SPH9S5X2/EPX+u8GQz6pPoR96Tk2c0NSas6crVyduIXBsreDY6Rjlob97fGMtpTwuhiSzH8dDQc+jvxXF2CRg5iwwZq+Q+KMursFB4AuBlUe7qSYJShbbMH9vV054XtsrbtY/DHaXUe1heFo/oAmwqOmfkHO+DJMYGyLLl+ZBntyzFq/R5rHuwMTB7ov+pqB1kY4iSvVvbYhmuh3RGJ3hnpM8aIcL7+XJPzNMKLYLimLwjHhwf2zSoalbkbbGgfTj2aQNwxgfuRV8ZC7EhjFX0lzd16kTZ9+m+sjbuHt48OvH4+Njwl7UfRr/nVZSfDO+iDbL3/uzZSRx2L0yduDEKW1uR7bIDG//flZDRmNIF//65XADF/4UECgkUEigk8IwECsKi0IZCAoUECglcXBJggtvSngQt7WcB6AhYwYSA1VusAoY0mHCNPVe7I//zbnfJz0FUsMKMiRUTJCZFkBi2nwMT/PzBNXbOAH0D+Jn4MAGy/5nsMJkBfGdyyEQboIfJEc9l4shEHBLA8uUexi4me0zMbALH+fwEzlatGVFgkzz730Kf8D91YkLFhN9WxtrKMVa8M0FjEmUkCuUyQoC6W9585zcmi5Y/9bE9Jowc4br8YRNXy4v68UyTE3kaSWHABs807xbus/NMEI3EyE9sqR/lp40/4U68j5WZeNbQ9gBsrLAG+GOFMeVFNwAIyastXXHSmQvyUN081zpSmSj1+0NaBB7GtWisdcXoXNofzie9scLpoIMrx2E+vxKhje5Rot3YN+YXlAwwNH0GQCGxCpjVlrcqQVgAyNFeAHBLS8fPZ/E6ACn6BbmITN6hpB0MtP7a0yYKIjYVRqumfRTKXm3e1Ssumo+Cp+tJJemN6sdFWACcATZTNwBzVswTcgLds1Xt1rctbNxSXQT25488OXca2KfNfD15WCzsHbpy8uGBG2tf73/+DgGHvy/vi3dm4H6azLX9yqhlpo26P/Dq8bs/9E3TX36ilEZHFETp67qGPmEx/WkX7IKtjIc0MgIWW2dt1koqPdHsC77P2/7PbzPPD7ecpFgGNFMMbAv97TeUeO6rlXoFu4u0+LQ8ArrdJbXvyIq7tXKbmw2fUtioz3aKQEH8R462L33Hsfaubz7auvTqhbhfO1p3HdO+DSBcj+l3vEIy0kcJWQE63a+E7mB/qSfoN2QXtpD+D3mCPkGOGciJLQBcZ4zgOytvgwPNVPnlOVh3o7ws9sjLIoW04LkKD9W+6rLh6ThJGtrDoqq9miva3+JAj5c8WU+D2p6W//K280bbsdeaib3eQ2nX5Xd5PccFsnoCWa2tkSnlQ28+pQSJDFi7dMgbKtvL43h7lxsPt+xqqhn7ghmROU2nUG/ZXivaKto9PP/iR17Uf2/SX1LwdJcQAoo0prQucGxZ+Ceeb4QBdhtyHZkRqo8+CnCMntO2L1MCHAe8ZNyj7QEzkSskHuMR/cvaK1+9074v84jKVv/roF0YT/Z3vuM5CcFGvivt28E9lBHimj74ylUfeOYPn/RSd2+12f5wVPKvPrF16NKehUaly5MvlEteot94rnlU0p9X86ZY6ZH5FehnK9K0+vZSGCbtf8y1+9R/eZ+4S/39vfrEViFfky0gMrLHK4JwmFZG8x7lcz0EgtkA9riinyD391AAiDMOQuLJU++HFCbvDvVH5AwIjCwyhrfznH3SJ9oG3VuLJDFZ8Gx0DNsJiWyhv5AF70u8G5Cf7QWS6ZuecyrXnyyv4vN0CSBb3kHppwDzS6Rdqz7nFApKxKfvBz3llr7Q3+zYRRik2RN9cwqJNK7QSlrvkzylsRHij/et5cdpRnP5jwqzNJtE/qPaGyMQAfLjnXJAQDBG0r7YQ96ZbY8XdB5d5J0e0pKyMW7Zu8Nq7bxdz7lt6uhAd1BK3I5rj28Th4Dtp3zYIXQMYhWPCmy/LRKg75Sk7JuTKJjUyUq5KxwOytF0qRpt7xmu3xM2yjvlcfEaySXzgpMnxXQax1Ot+dnZJAxvXIGs4DJIPmwgtp52OIPRWK0ixflCAoUECgkUErjwJFAQFhdemxY1KiRQSKCQwKoSEOicCqA1EJAYtIDWbMDJZBtghQkPE4Utbs/PeyIsAEAthBPgCpMimwQxkeAcEyKusdVinAcMgJzgfu4B2GPM4ZOJtHlVAEzwbEAzm4BTPib0PIeJFyC7TRoBfZjcL8agWXw+4IN5Uljd8qvWDBjQZdlki+cxmbMQF3wnfyaDfOdeADsmZORv8attVbMRMeRnKx4pu5EmlAEQhP+ppxEpeVLFJqvcz7Xcz7V2DbJaToRk4B8P7dSDT/LmWpuU2gSaMlA/QChkSN04d5cSK4l/tJMXYDdtBMjGsyGnPqb0IQgKdAWd6Tzzgv6oJuGx97bfGn21fcsVCmZysOK15wU4tQQ2AXbRL9CD5/JAzvQ90UMZgI3XwduUbHV/foX0mM4DKqA3gKGEjAC4elbhoDZQKcpIX0ev0BsL5ZYRW0rosBBmD+x4Zibomd8RTlBG6kI4HGwEpAXgHWU1TwRb0YyOrgcsPKPIBiKLdbR+Qv7km3l2CcQ8WE7D47W4KfzEe5UCfFwvsBrb8v5/3Padk0/3XD79pw/9JNdTJvoC8qQ+2AD6K/XgM98PM0ICkmTx8z5v06/dd9b+skLoLa5vC3BGPrT39ytBD26Xp8UlhxofD0RU9Fb8RVz2qp4fcRPhQwJCJ9HHe1WZykj5xCUDpanPzcf98/KwmJX+nlQbbFaiTbIyG1ApOWFb0RfsG+AWz+cc+VFXgKnLlADXaV/KhVwgdFlFjr3hOgiOo9q/4nA7ce/VeuMfzgr4jCfaEtnUIS64J/rAfftarXbkhVE8ezLxTj4ZlgdORO5J5THiPL9LKOCESgyhBXlKW3CfHZTjbiV0EHtMzKx/w4+AxKp3RkzgTaHQWNm5sr+4Ebk2HHfaz8JJRn8n74u+O6e+8+BNvfffNVI++RXtbQHoZyGZco9b/HqWcGn8jK6Y1wQkDvIBoGPcYwwkX0BL7DzAMeQA4w2EBrKdVwPRL7arIWyMhWigfyUbAJjNM48xEgKG8Ryvjld0ynO2vR24jpQ/6IeMGyvF2Ed//izRZiQzg73zSnddueeI3zvXKAdRTLsAcKJX1IGxFH2CmHm5EoQrB3Ukb+Sw1gFDB5HHQdimF2JjIr/0H1p+9dp60H3JeGXkEZ3bLZJitj+a3av+ffzBwZsf2dk43L52/omDvdG8ebqQh5F36Gh+LLbf1iqP/W6LOLATeGyMqQyj6Jr2jlFYt2507prJcOS2kh/OtOMqdg/5AMTimUX9kQdtR3+ETDTiYj1lMIKDfgKwnH8XQg+oG7/xLsVzAbjXvZ/GegpwoV2jzZ2TW17+FuwL+olHDu/I2aE9F1xzfkoeFtmrYJ6sWBJDFAYDIhlq3QPNQb8U0/8hVvMH71z0hVXDnImsONSYrY09+ulrtjVmarfKxmMfbM823n/Nqxm9Y2y1UH3YZ2yLlQ3bBPHCuwM6RkLnyAM9yMJVKf+hqFVyk4cHXd/mub6+LXNbk9ivawNu9Im8sVumP4yZvJ9w7Ja+b9J1W7TfRiyyZkibb1/TO7zABt7dIm4unzg4VGnXtQ2HelwaRa3m/PTh1sIcdmClAzKRMvI8FmU8q3eBVfIuThcSKCRQSKCQwDegBArC4huw0YoiFxIoJFBI4FwkIAA6A4D0GQuQBsQA3GDiA3gF0IDrN5OTq92+dzzoLn8nq52Y+DCxNqKA/5lYM+li8s+khgkQ55jkcB0TD4vfy8TDPAKMTGC1FtdbeBVAI0BYVmCTB/cAkjH5IjHRAzxm7DJiwbw5jBSwcc3+t5An9kwDKiBUAPItTArlMNd5Job8D+gEaMmkHyBq+QTVgEkjYwADkIN5V1AWIxMoh5EQ3AfgS54GhurrUmgAy9fKbJM2rs2P21zHs83bwwgcAFrKwQFoBmDB5JsJYMnd6TEBB5xC7oDhAJTkQVgBPgfRDW42XenkdUF+dAiZRvqZhv+F+iuachZoDnkzYVueFSIraKNsRewGgMNzlRP9CBACAOw/Kll/IuwIoCf9A8CAVb30GVb8mxfIvxa5hE6SDMTP1KVTccCQlBBS/N9BsbE1AOIAoKz4p362ShR9NeDtfJef/JDnU1p9vb/p1bqafo2+wSrOj2qD5rmT1S1TSvHjfddGH9zx/Ss+f6348uZFcUbIpw1oguTFKnn66IeV9ivdq3RNmM6/7eG5/9p3S/9/uV0bcNP+7qWDv+e+NPNLDzTiE/cp/NHQ1+ZfdPzhuZccExh/UjqLHTfvEOxpO6+7nfAzdREXkHDIZlQJoAgQFWCZ9gBYZSxgZS8EJ3qGLQZcpu04IDQ+Lzpqtp64T+YIi3fq/N/LywKddPK06Fy++PEDr7g8G3/kdRHt0U4S00FZeJn/L5EXTCmSUJ8aAMCNsYH7P6FyAtrngSvKjDcC9hp7SFi0lyq9PE4DXegP7KyOZc+aiobxsJgWifN0K+kqK1TWJsloj7yATjyxcOPQo/PfdImuf4jNytfbv1fwrsBOA7BB+iI7xkkIF77zm3lLAEgjYz7RfeqXEQKqs7byTbvVgW5RRRW4yrM+wfV5wiar1yoHMuI+xjRkg92gTzLWMI4xFtu4cLZ87DcjYvLX4k00psR4AtlCn6Y+rRt/8QDEHffQv9EXdJVyoNPYBBZI/JXSazvnGE/Rz1cq4cmIXjEu0f5/2LkGPaDs9Evambo9qr68c67UV5st9S8sBD1jd2z5tuaDAzf19UdzJ26Z/sqnRUju/6dtb+x6svfq4flSn9cTzc9tbp+a//YTnwh/5anfSpf103O1ObZYAFn/k9LbpId4VmQE2dcXbhFJ1ve9A8HU30gPGU9I2G9kwthLfRljeM9CZub5cZqn3FlsEOW3kIKQOWNKvJfR3rQPOsS7DkdF+ttar6537rkYP1YFygW5u9bCtPODwJVqPS25F572XiiyoXpq38gV2553Mg5KccsrJfgGvlHpJR1BLoWwW0GwszKGHzy5b2Sv0su0J8S36xre8ehvtCF9Gv3hoK9hk+lj2EP6Ie97lJ2FQNyHTmKb6JO8zxpJwnt/3muU34dFOrgjj20fEFlxlUiHx4YvnepVaCjIDvQSe0W/Jinam9cnxnA2apfa9amu3rnxnjRN/ZO1vla/wldpA25/RPdO1PqajzQVZFZF/1aVpi8olW8OymUvap3R7TjBO83dShmR26lLp7rFRyGBQgKFBAoJXIwSKAiLi7HVizoXEigkUEjgGQmwmv5nOpMZACwADSZATHS3u/3vmhBhcae+v0XJVhvb6lZbdcyKq1El8ygAoGFCZBNuwH8mI4A0HIw93EviOpuMWRgNABbKwfW28poJE2SFrYLlM78JNvkbOWEzIfLnPsphK6dtIso5gBQAHiZ5PIvv5gViYA+gnU3sbHU19xr5QH0MqAWZIw8Le2XXcL2Vz8gMwC1WU3I9xAHPZ2JpMsyTEyYrI3GsHDybfLnHyAp+Q3ZMXqkzk1zAT8LxAA4BkmSrt5VoY8rKSmbqiHyZjKITF+MR/F/Vd3l/0P659Lgiiky7AWSDjmWEgIAe83551ptur1OotCXkF/0Cks68iHbrO2AF5ygX/dU2e402EAd9ncU4/bI1NuXm4vUAf9b/+DS7kD3oXEOOrUEqZP2vs7FxBqTrwJ7hebBeQPhZyW0jN0nG7GkxpnvopwBhKlv6z83k1FNHW3fv2FF99Z9pX4tsxftV3T989LH5P7rvKws3H71r6o0vFSB/k1a7og8AoPR/iGfAytOATyuP6t2QPIjrzzXola2yx25AlpntRD7YJmtfbCK2E3tUj0DbvdM2Hd4VJ+lQ4Hsm59NEYID/u57xVLF9iigzNpzwKQBr2CNWOLchLZz7McuHcnAP5eT3XUoflUvPK/Y2nt/eU7/+uktr+35Q+wY0Hl144ee6/frIrtq+x+VN8+W5aPDFc3H//RPh1qMiLvAsfL4SMpjphOVZTVan1SH3jwGCECajSsiKvssiAFa8Y+dtDMHOkgAHGfewwVzXpUyGVakv6vObFGNlV3catdoiXkLFnnEK46NrljxkVitI53wGXishe+TDvTyP/gbZRBvjaWAA9hrZLf2s5sp0goPxHv1kTKG9bHzD28j694LIi7wHFbrMtWNK2FPaF5KC/9Ezyko5AfzRNcZO/v9jJUBZyo08U5EUc3dtfs2Jv9r1lk2z5YGgFjceEdk4Mxf0XaHN1uv/sOO7d4ZeeST0y3gYodvHZ0r9Vx6t7ag93H/j47911dtD9+6lMGNLFTzHL4nCsB3V896tMnx7K+26Sv+nTzeu9WaioVDERZeIMQUMSvbK+wedYNU94wvvDLQFsqG+ANuE98NrjnZa1etnhfLaOwZjOGMVbW9gutmTsCAr1m7pjpcF8vvTTvt8d06WTiGN5AwWuHIUHa329B3Xd3QUW8JRWZju+hZ5SNxf7WlD/KLL9BU7GHewX8vJw8wTUZ4Op448tm147mRfVd9LhJnSAQm90kHeEMfXKfFeQF/C/mODeAbvlST+z8Iy5Q6ejx3HDqGT2aFyu+NPbRnsn5nbrv0zGiIuMpJcB++Pf6B0vcrUH7eDXhETM7On+k61FypXV3rCHoV/GipV4l3lrnZan+p+3PPCA90DJ72pI9tm09gdjNqNm5sLM9oLpJntCbLsYJ5xtxKeR+jrirZ4+U3F/4UECgkUEigkcGFLoCAsLuz2LWpXSKCQQCGBtSTABIGVX4A3gKAcTL6YyLBS9DXus+UPuFeHBsRAVox2rjMPAgAjA5GYBNkqT661SbOFdDJwnyyYsDN5u1KJ1ZUk/gfIZBIPqMH/gC957wwm4XgDMNmnDBaqiYmVeVYY4M8kkHN4GZg3B/lRP0ASWxlLuYxQoWxMlpj0A8qRP8+xkDeUyZ7DtfmDMhvBQBm4lny4nwnkl5WQBasfWUXGb5SH+hK6w448IWLnkLHJLy9Hvhv5QLkpJ+AU31l5x+SP5z3hHvoOJqaEDTAgngk1suF/yvIVpbtz5bhovgowD//+E+HUiWTLv5xKR1oKLYJMAecAgOLnmhBYJmjamna0mProMYAdq42NsDIyz7wTzqmttCJ+pftNl/M6uCIxsXwl/fLMlhES6yE3zqk+K93cAevs2auuoj3vD15Hhrm9LbAbAK3YAOzn40kavmBf/QMuTGd+anfX9/0t2Q2Vr3/LLQO/eedHJ8K9Ws09I7AUIgN7RggQW72fPRmSYBVCB/0CTMNWQ9xiW7FP5v3CSl1C+hhJxrXYXVbCIr8MFBdpgY3JDoSrpba7PnbPnsOvv/3q9bRzdksnX8pBfwOsNUIaWeRJWnsUz+c6xptIAPGdh5u7dz5Vf0GPyJuPyouiPhMNN8KguiNoXRqeCrcdno6GN2sfC8IJYWux67ZKmTHPxrj1lJkycC95EO7JPLG4F8CZ8lI22sFCNGFnAaXpyxaahzwgAhhDy6rQgK+Y8PI5ubTmokN1F+y4PKm3etJ4QSge9616LCMUE+mTjX0sAGDfj3uUAP7XRVZIRg/LBj6pz70igz6srPf4vwAAIABJREFUNdPTkt18xW/Z/jJtvIJWK1COvEhEXuSBd4h6xkXINfQMOd2vhC5a+CLkYmEMLU5/Q14U7t/f9KcjR6s7bmgGNXS9L/aC7D1EZS2prLQj9eOTPNAndBewFiLs75Qe62xAveH+fxbSNnnDZ/+SEIKNwfL4vRWvdWV/aaYlmUVDpfEJeT0dPN7e2VQErc/FafbuQtnwwrFFH/Q5xmtIOvQZW09fZPyhDhs5jLSy9zBkTbL/N5LXxXwt+jim9P90ZHe7Pq9AIHHYcs3ZKcIc7S7Xuo75YizkabEkqzT2Ny9MdQ9p82psMoQA/Zv+SJ60P22EPtqBDTgq74y6wij1i6h4Ut4O6wmVZvdDgKI79h6LzvAcs0voFvnlSRL6He97vLPi9ZSFSFUZXGOmy/UM1bu1GXdVpMUBhXwiH/SHeYKuSwfjMFhoztcmfD/d1b9tbjhqlir16a6uWm8rEskxXaqESdhI+7WfxaZab23Pqf1RHIehi9stPSNWOq378a7FWMLiGuxVQVbklKP4WkigkEAhgYtZAgVhcTG3flH3QgKFBC56CQhErCtUCzMHQoIwqQIEACgAhAE4qipwb4/g2q+6oMYqrmzCpoOJkYV/AvwHELBwBkzSAB4AczhnE28jNpaD7kyYmNTxXCZR5AuwzsQFEI2xyjweeDb5sWoVwmN5iCQLo5QPAcXkjQkRkzWeTbnI3zwwyANAxVaB2gTfwFojD/J5Uo48gcD/HFY3IzWM2KBuXG+rR/9G3z+g9J865eJ689ywvPMhofLPWh4aimfYRJTfAIQoB5NRwBtk+LAWn5bdxCcsTj2ftDGTUGQBKIgOJOiEVeZi+gTUfUsj070xJfTXViqjexsFjTYsunV4CDyn7ZInHEReoD/on31a2BM+l8AENlbecEUv4BtWCBdktc0TjHZumexO8yCgH9vKdb4/rE24q8db97IB99tKXg8rXbVPw9B73j7q3vi56QTSAPKRvg7ww70Qotk+CKuJHAJHZQZIw9birUBYGsLUoP+QEBZC5DJ9N4+fW/WdFeLYxcwz7VDTaRuDjOh8VcdoQkJDzp4BsqPny+SEHLCPgFU8B7sFUGt7J2AzsU8rAfZ2r7t/5pvHH5h75W6B6tufalw/X/Ua+1pJVeSKRjiXfq03mN03Hm5rCtSGsLWxCAIGmfFc6ko5zlj6uwLhQzWpP/chd+pKPpSVumNXKRtjKMAhALSFhuI8382jb0onZpQhY2BX4nk9Tee/vuzSjytM1MKEV9k9mNaP/Pj7vr6wO65jh+LOniD6uvrRCTGGHiA7nsWYQzuPKv0bpQygtIP9Pkj6G2qD6Ie0BwPeDgfHmlc9urf+/Pkj7dF0Lhpoi7Bol70wffr1N66773f2eck/jnJBWOQJURvjIHny413WxgPfkXFijN3IGFkx5kFMoKs9Kjv1IV/eRXg3wF7y/oHe0A8Y5winx/0PqE2Ry0b2CFkq/0qbrj8wNxVsLh/rU9ixie3VQ1+diwe7eoOZo5dUnz7V355+9GS4/ZDKSLmoH5UZ7ZQJIBldJ/QOZCALSCyEj3Q305+zklUUbIXxw4iLAvxdarn1f5GXRay9LNAhvKDep4TNsPdfkRZtFzbnXZIMXym2whbN8IB5ERm9syf7XrL1ivF92oh6QhtvYyPQT2wLOoud2dtp74z4ldfCbNgsp9pge0phlvD6+rb1lzaz8eiWvTNCgLHgCLKPfkb56Cf0GXQPPUPneAfEdn1WCUIm88hJYs9NHRn4okI6pQPbZw9Wu9s3eX5Kv7ldPfOYNtl+Qp4Yuxtzte3ysijr+ljhodL+kXk/qEYH4iidipotvzmX1qJWtKkxc+oNrfn0kgR3PIgdNrR45sAGP6r0D0rY/hU98zYgi+LSQgKFBAoJFBK4gCRQEBYXUGMWVSkkUEigkMCzlADAxFuVWE0LAMXkB0CAyT4ToBvcod/9lBv9VSZbo0pMtpjYMBFmEsaEGwDcQBwjMiz2vsWi5fc82J4H8QDDyJOQGeTLqkhWc1EWVnflQTfAffLmk8OeZ6twbTbEZx7EALShLAAaJCZvlJvnkXhGFiamkyy/fMgl+93CY9k4mgdYzDvD8qOM1I3JL6sqP6LEymlWLgMg8Zz8vh0G4uS9OPLneKatqrfykDd5ct5WawI8HlBiopq44++FyGBlMfVm8g2AAzBo8dQBcNCFi/1AhgBGNvkHJNzwatz/lYXYCW9FEbMwV3nvEZEVRlQYcYfuUn/0hP5r5FuiazmfFMTFohfDssPIHiMj6ZdmW7h0sV92dGuVzbi5DnsyrRXz3s+84C/TBw/9j7/Q/7+kRB92vYH7ic0V9/vHWhmADrBJv6cwAFHYt7PqbsfrxGLgQ1oCpGGnsP/kYQQ2ILvpAjYEGw2Y1xgqZ2Ucs/r7vtezaaA7+Ng9T7JXRUa8rAGyU0bANew1ZDT/81w+CR104O1Pv4f8zyATyFsJWVMmxoo4jCuluusBJByXt8Xjc/HAYa1yRxaUF1KGEE7s5cMz+J86U18Lg3UGGJ9rX7PFlNXCpfCJneATcBDywjxl8BxkDxz6y9KYpz7D7xF7ClAO7VsxpR83qcLDofObCmGV9qXRpv40GiilSXeQpodanj9XTZM5yTSz/2sRFx0PiEi6Qz3xYsAzBjlBXgCMEzbsZoUpekM7qdQlJ0/Ezs3H27umBLy3j7RGpw81L1cYrcGF2WiwV4A7K8EZo7eq3BZ2EO+zNckLkRYrHfn+wO9ZPh1Z5/M0m4Rced9gvAP4BXRlnwsICfSfMZ7QNUbYU9dRJVag2/gI4Ub/oN0n9azmespvhV+tnyv0U1cj6R6Wd4V/MtzxcDOpbdX3o7uqY18W+fPEbDR0SJ4qgL5GKBLSjz60W+nVSoDIgMvUD1KNNubdxrzrzNvOilJ8PscS6JAW6B7vadiP3CEKuVl3zZmJsj+05UBQrkAQLHn8arPsSn2ma6ivHE8J+Edf0VXGUOw276HoLLYhlFfDnhNPbf6KNr2+cuZEP3tCsJhlXZ5QnQLZu4qVD/3HjtLf6Q94VqHz9Af0Cdtj74r0I+w8JMkvWAYiT950av/wEyIrHtp61ckH+jfPv0q9KhSxUgmbpa3yABnSZ7U5V2u165XpnsH6zsZ8de7UI9ue6N003pPEM7vaC8nljVlve2s+coF8oJLoDLKC0Gd/pQShixcYcikIttP0rPinkEAhgUICF7cECsLi4m7/ovaFBAoJFBIgdvyDWoP6oxIFK52YUAFcM3kGSAFsG3NH/niLu+ztVQXu5RomQhxMilhByljCd+4DGGBCDiEA4MDkiN+5h++2qtPACFu5bdcDJjB5wmsDcMxWri2fkNnEy8B7nskkjEkh4IztP2BeFUwYAQus3EwGuZ7y2kTUvEIsjJMRBgaI5Veccy5PVpCv1cWIFCM6jMihPhAIt3TKAoEAWEEZbPPyThGXyml5mrwoM/nmiRXOAXwAlvHdwBvb8+KElszNuyd+mv/HlGgLJoXICYCEvGnXAF3IF+Bi+r7CCtULiqSwthTghu6YNxH9BJ2ZB0ydmK4HC412EAR+sJB4pakw7ekr+cPVwGsfazsBcm7wZOgmBJLPbqt4s1Ki9pFm2upsjLwmaHkR6RN9nj5tNoe+BvDOCl1sEUQhIDn9Dzu75grqXPgdQB02YyXW94TvuVf9223efb9/MD2mBayAnUaQYAs3soLcwGPKxz4DfGKfqAdgL7YLm4WNoMwGvLaERWFbluK0KzzKzGBfNZicqXPvGSDUSqvBO54e+3U9oU2oH/cBaAHUQvYwvmSr4pWWH6bT2HDkgm1GFuwdMO1SH8CRVegQMwZqM9Zhe2kb2ol8Lea/eUis8KhsrOM6xhaIfZ4DSYTMsM3YYdoXsDADJJVENC15LWV5dkKwGfEc3fpAMq4G+GelQ23Pu0UQ342RvAa60vjuQ0FXSYTGoB+nYclLW9uSloV7Whe419GdUMQFpBDypGxP1eOetvZbGGvE3Q8fa1+SiqwY8F362icWbrryZLjtZQqpdVLEBeHGdsnzolufEEK0BWQ7dYXgOohMNwL6ryRUO7eMEEDWtC16RJ3RSWRP4j2B8xZaB0CWazlPPdEFFmFAcgDKGumKzTOvOSOanq3typfvcnn3vDx0lVFtrr2gbYkXRDptnok2QYxpr5cS+oG3hIHFPJPns7qcerHCnWsop+3nwnsQ1/R3PEJWbO81vPPOJu7it7UlYO9Xf6ZLWfCxtBcEYY2ac1NDXhDEPUNbpz3fH8GBQATFfFd/M1LYpOr8ZPfBga1z6CV6yIHOor+8d/6jCIBRgf4H9335sj55LVyWxt5bdW4jZAV55hfM5GtEX/9WJfos9hv9w6bbQh7qhg2z9wB738zyUPmvmRvvfceOa4+zoAhb2ZBzxOHp4wOfPb5ny8u0d8VV8q5I/SCdCxslOYbF5bidXJ9E4ZC8K66aO+W7+QmxHE2RFfLa6ByMG7yj3qPEOAJZgWeF7bWTL3/2XcTRGeeKE4UECgkUEigkcHFIoCAsLo52LmpZSKCQQCGBtSTwIV1AmAgAIgAAJlNMlJlcXePa4wfd9J1fdEOve1EnIws3wO9Meph4APKQ2C+BCTdjDBMzIy4AHGyfCbKxlap85xpAJSYyeBsAWtkeFgak5QkAqw+THJ4DOGHABvnyLLseQApvAib7gEzmTcF9efDWgD5bGW3PyBMWds7Kb+BZvi7kb3nwaR4clIeJKCveCK8FSIGsWHEHeAb5w+/ck8837zFi5JCVibqNKZmniJEZyIM2oW1OupPvY/Uak+1RJSanTBq5BwAKgId80YHiuIAlINAL3QJ4yGL219LEr7ik/eIPjoV7DoynSVDunptP+qNKeeBw2yv1Bdp5vJQoTE1QfaLhtm2veqXJyBs/0nLjiUsbisfujrfTU/0lV+/5yHR9Ic76v4W+OU2S5wqqrQBkUhezDfRdI+x4rvXxpTKc6/M3oBb0QewMINFlSgBcFgoOzwXIYEB/AH76P+DRUdXP9gZY8VFWfrxZBHazyv3FqvxvSQjf+YYR72cPNt3//eGTaRIu7idxhxLgPjKhTTZyIFPacEwJm4xtYvUt+WJPsC0AwmZfk22VzN4aUcuzWsoEG2Y2NpFXAOdXBIblKcBvBtQCgltIHwBbno/8kCPPXYmwQBcgtwnHRNmxi2yCa2MTBIKFVKMM5IPdA9DmPsBixiqeR50ZB1d7FvWmDwFEY6+RM3lwDzJC5rTt+P0v8q2sZrf5zUh2CzOXXaNrI7UtG8PvFznxGhVya8MLug/5Xdd2u/gLX9PG0fuC7sZrw3ELW+VJphkKuJanBddwdMJENR+Zf1H7RHtnMBmN+KfC7Uma+k/LQ2BE3gCHakF95mR7+/fIO6B3Pu67Qp4pNe0HwriMXCHd8E6BTMKGoM//qAT5ti7yxMqyzk8jBJA3zwJ0Rc60K32LvgTIT/loL3uPoHxcQ3tSrpcr4XFjXgzoKn2PfB/qkFhGHp1RtLPYDhvT0U1InOtE6gASP+alspGe/0IRPWOSIYAs4/vyZ9i+Ep/Ub9xn7wEsKuAdiIP3ILxIPqPE+84Zcj7LHjVn1KU48awkgH2D5Ltb6fvzOSRR27Xnp0dKldqBau9gl+e7et/m+c+LsLix0qWwUa0Stn502VPt/fBReVPc/+R9V/Q2Z2s/qb0vbj89WtK6y7rEBiy7Ax2in3Kge0bMmq5xnn4FmQJxhu3l/Ts7IF9KFcV6Sr2tSuJRU7bquLxUjp4a3DY7Iq+QmbmJ7rrvR5vazX7xNe1qYy7aeXJvsLNU9l1DvTBuQ1YQZmqpZOgzXhXIEwKc0IVZqFIRE8+WOFy3oIoLCwkUEigkUEjgG0sCBWHxjdVeRWkLCRQSKCTwnEhAK+vvkZcFYA+TbgP2mUyzAniL1unGbuy3Pdf/8sdd0MWkH4CGST8THwMKLYQHIBCAHeeZgHAdYEd+Q27zkGCCbisnAe4BEAByWInMdwMkbSKTB/N5nq30ZSJvq5cpH8+zSaF5W7Di2MqDHM2DwlZs8r95LtiKZwAJ8+4wgJR7rRz58E/56+y7EQu2opNysSkrAATnWPHGZJF8kIU9I/9pZbU8AWIoJ+0DUPMnnbqzcg5QhrYhL7wuyq559LD7+lt5Hr8BrNCmtA3XAOKR75fRAR5UHBe0BNAb+gF9tNGbRkcuSRrl673GpkOTaSBorDuoJH2nouBKhfXZMlDxeuVWFSuw9oKWWA9PNv1oQespr+v2xu6c0hYKnndFO3F4RR3S6v5DWmnf0CfgsG0u/FwI00g5+rXZFvQa8Jj+ZTYB0Nj66b+WtwzPw54AltO/sVHYI0ChjypB5BLuBVCId3AAJMBVCEXCFRlpsVLooyVZCtgmvNCeMHH/b8V331n13e6fu8T7jfHQ/fndU+ljSZrJgDZYDchaT7uYFxZlwmYYIZHto6C0VEZ5B8QC3AFU397J+MqdW/or+w9PcR31B5BirFgLkOJ6QGnaEvvEeITMWAWMPJEVXgt50NbqSBn3K2HrIIU/pzSmhIyNrMDLgn07yIP6kLgHxgQwHiKZ3ygrq4qXe3QYMWJgOTKGwCF/fjOvNYgLG18ot+0xZIQFz7VY7TwrkyleF5Ilz/yEBEXddwkl3B6k/mzoeeOTXvmKT5c3T4yU2vH3tI4l6yUqlM/SAWlR+9B7KKuRaIwbr1Pqf6J+w1O+FxOOqtkTzE9pE+lh38XsA3I08KKn0rQMIA/JTVsD+FPGNyl9RDKlvzEmrdjXniVhiJwsTCUgPu8o5I/sIASR7V2dc7QF8jc9s+vu1Dna9LuU0Fnsxrd0rqUutCUkCMTHRsMuIUfKwbsKbc7/s5KRzKBWyS+Sh4zxALP2LqOvpx2Uk3GcBQP0FXQdEJe60DboIXIlb/RnRUJ4eabF/+dHAoDo2svCiFraCNtNiKXsSMUwhM2GWxg/dlnq0s9Wu2raPDuZFGHhdQ00dvWWEmwLfcMIKNobr4JjIgH65KlwYvrYwKu1dwUE6Pk+jKwgX8Yk3muxk9SHccr6FnpPXzjNkxnypN2oOHl+jGvj7S9qA+5v1l4WWzbtmv4hkTGHT+3vORK1FMKu2aq1FrTrThL2Ru3ZkfY85sxzEWRFIq+MxHUp2UG4K/osBAl9IrOVhRfF+W76Ir9CAoUECglcGBIoCIsLox2LWhQSKCRQSOB8SOA+ZQLY81WlFytZmCWAjcBNfuZat/DQpOu/NQsh05nw2CSa5wOIG2jAKiom6QA1i/c/AyYwm2GiwmTKwEVAdu5lEsXYZAAP+edBNyMADDADmAIwsNBPtkLRQHumSQBKFqoKsCJPWlBuA944z7MBjABCbKU019hz86QFeVP+vCcI13LkATWbBCIDJoVspmhED6CPkR75ehrZYiuXuZfnUVbKyKQTgOXjSkygLYwX5UYm5El7POYmPw4hQnvSZrZvh5EztDXX0vbFcQFLoONdge5s02a+Vyg2/pM3xLOBFO2yGb88X0/C7i1xu9znl4cG/Pbl1ZI/0OV55fG21zcXp8cHAm/6RNv3K0Fwyam2n8xEfqil2emlXW6uy/fmldHc/kbaFmiOvtMnzU6sB6her+TpB9gTbAegNuAeK5cBjNFtQCHO0S9Z0g/oRx86bKuoz1fomhUKTJ8124WdMTAbMBL7Q3/kPDYK+0S/ZQU4crJQN8RBp2+Pdcq9KsAPafHhp2a/eGnVnVBYqK1lz23/zSu8//TvHkv/6+MLme3GDgDOe+up8yqAch5kPfsK+kOzEA2Unbb/9d6eKvskUA7ay2LxryC2M06xUp68AAWRGTbzGiVsnBHctlqdm01GPIP7AOZofwhYI5Dm8zLohIYCRAQgJm/u4WDMok2sPQCIyddCpfB87CmEH/cxXuGRgR2HMMces0o5FIFj+gBBSPtjm9Vj0gEtU6ZOjEv0FQg+QLsMbMfTQqQFHi1lVexKAd+bFryAMQPd6j3lV46ccpW5d3VfRXirTrFX3HR56Tf70rEB9CHKwx4WfNJvAMYrelZJ3gBtNXSPPC4Oyzvga1pVPaC9F9SXvJP63bwuIQ/QYQP8kQNePQa0n/HstU6ssDcE5aSfI1f6CH2bBPmFbkPwoRPoAnpmQH6eMEE30AXAUXST1fGQh1xLe9ieAvwGMUZeZxyr7FthYzREF7pwtxK2BplQPogwdOMgz8vvE7TCI+in1JH6oG+0Cx5Ao0rI9t7Oecpr708rFbU49xxIoENaoDOQX+jKG5V+3h6VCo0P2w03d/xAtd1Tndh5XTw9MjrTp9BQ2+WRAJmOTUG/0OeMqBYZ8Ghzrto1dXQgSmKfdkd3aPv7lfCGHVNCl7Af5+tA5/E2xiOKsYY+hg2iL9MveL69m4qA8BQWyp+IWqVSq17ZIgKGMUAh4lwlKEe1Wu9MPWykvXE72tJuzA/jbcK+HkkUyyireyxaZnTWjn/RF2yrESWrhfg7X/Ut8ikkUEigkEAhgW9wCRSExTd4AxbFLyRQSKCQwPmSgFbY75GXBRNsPB2Y9I8pARYApDChmXN7f7XqbvzUuIL0MvFiOsIk21YxA3xwX55EABBiQsR5Jjvkw3VMisiX38y7AOCfySCAI9eQ/1LYEX23Fb5GLDCBZOUhIBPgIGUywsO8Owyw4jrAQg57phEJTJ4AyQAruJ7VmEwUTQ4GTBhpQV0ov4W8yoNbtqrWiI28pwWTRe7jOUwaLd687V8B+sQ1Fj7EPFj43cBC5M3El1WXY0pMOgHpICQ4n/cumXStw19we37h1ToPyGP7eyAjvC+u7cjiKG2fSaY4LmQJoE8VrYOMpKQDDRdc/njQV70pnr1CG/qGE5Hr7U3afVEQDMelZPvEbKO3r+zXXbVc0grvkTj1p4e9OPbFdkw4/5Kra/GeU20Xv6DHLx9tu117G+5ahYgCnAcItlXn6Bp6Sr9ea3X9WrKnLwF+A1oCEGJLAF4s/BsEAOdtBSnkK/2FvkM50PGgs8nuWT0Y1irI8t87QDD9lDJRvhs6ZcU2QApynn5o3mTYJyvXqL7T7+mjclJR9HutsL8sbhw+EHSddUPjH3wkmfmlUe8Nb96cbYacHb8y6r/u559MnpjRJgg8Yz1kxUbru8r1RlTxc0/ge8gcG0+9rI3W4xVA26BD2GuAW8Yk27AcgIvzi+PRM2MEv5P4jWuwiwC+2EPaYCXdQ/7oD2QDIbYgIoxc+oHOb7YJuZG92GzsM2QxZaPNsb+2xwbjUEukgz6WQhRyHQB/NZHriw7afreIi4aIC41haY8+GTMpJ3Vd+ImdXvTuI+pmi6A3Ywn1Mm8/nmVeRquGMeJB+SOno4yTJPoH+QCQMh5Rf74DXA4JcNSeGhnoqDIGjBWMh9SV31/ZKZf1I8hDxiDaBblTl3PxaqJcRkryXNraQk7yG4SR7cWRhaNcgxBgc3PeEwhfRV7oJW3KqnbGQvIjn893PtdjqyzsG6QaeoHOoefmmcQ7Be2KLq/X3tg7Bu8k6Bn6QDtBWGDbKCdtNKZ0LvLV7cWxEQl0NuDGtiB/+uMSYZHlIwYiiePbWvXG1af2Re/Z8fx036DeZL0gazfalfvYvwxdqTdmuj619/7drdkTfVeIGOB9k/bENtzeKRf97Lk40CvKlD94rnnvoLfZHhoiK+U9Uh5OEq9LNWhoT4tP+IpyF7XTG/wgfLrW194btxu3J4k/DFERR6FLwlVV/ZeVJbaBfoZdY5w+Own+XNS+yLOQQCGBQgKFBL6hJFAQFt9QzVUUtpBAIYFCAs+5BN6nJ/y0EqsCAScsRjcTnK+4qbsvc/XHA9dzXcv5AYCUgelM3gHMMzBGCUAAwAEwYFQJsJzfADIA0riP68mDST6/MybxPEAkgAQmeUYAGMlgXgjMigAguR5QivP5/SmMMLDZE3nz/DyhoH+zg+cDsAISAETZqtds1amSkTIGJliYCltBTp2437xJmITZyjXziMiv0gV0QD62lwQTOMCTvEu+haaiHuRv5acM5I+8ADkBQe9WYiLIZBiZLsYpTqIxd/yvb3XxPHVAVkyECU/B77Qtz+e5tHlxXAQS6EnjLu1ZcVAb6/r6XpOSAVReq5j59WrJm1ec6ZH5RvsyV0m2uiiptqNothYLrdCmopWa39+tINU6t6+RxFO3ld3059qlTU/Oe327ujxIPvYt6FPneZ46GeAiIDA6Par0SQGG6PyKQODy1f2rrGimX0IGvKyj+4CLFtoHUJMV+fQ3QELbaBeQEsCYVdAQnFw3rfxZCZ6tyD5PgD79lH4FYAvJC+hDfVldSx+DYMTmAZYC1GBb8G7BdtEP1RbpMQnnSClNt5dc+gotbr1TGy577kPT868MJ+ZeGU6mK4QAKv3ugTTsD9yfvnaT9++Vj7uq273wFYPeDZ+dSj+nPUXWA7xy2/k+eC52y9rcwHazy2d7HvdyH7YY22iEB+GAaNs8sYs9x+4id4huwpNxP2MIz8L2cf8ZBwB3x+uGEH20z/cpoScQTNxHO0I0YDu/oIQuEwKJ/QgoH/+jQ9hqnkVYIfQN+4y9zjwiRExsVoFGhWf2CtQc0XffS9NB/V9NvVQuTh7gncaedEHEBfVNvnXYa4qwwPOC5xp4ja5DrlymZETdinsanFnb7AxjLaA6cqSMyAldZIymX2ALKAvyYnxADhwW3o1ymP4SBgodZuw0sBNgHXmhz4Tjsj0lVinOqqetL9GfSQC8tkKdvoRe0daUFZmvixzptDfvNdxjHjt4hXAQCgw7gX6hdxYScqVCUj76MmVj/LWQjhAXANrkg75TPnRnox5m9j7xKt3L+w3tji5ByBJeiHZ6jxKy+P+rf68klwv+XIe0YGyj//2l0o8sr3Qap8Mn9/o/9dhnyr90y5vb3bW+dJe8LMqyENgMdOKwQkGdmji46WsLU91XyrsCbw36NWPFagd9ieeVGo+/AAAgAElEQVTaxt3PhayxCeg9usb7bFvl3Nycr87NHO/d079lpqRQV1tdkJZkp3rClhvc+/nkrQoHtSWOIu1V0crCY+nAhmFr7LhHX7DT9CvsWWbjlArdfS5ascizkEAhgUICF5gECsLiAmvQojqFBAoJFBI4Fwlopf0BeVkAOABC3KbEhJnJB0AFYTN63In31d3udzK5AVABTLDQCkzSmZQBGpIHQBArM/mfSTu/c55JEQmAj4mRrTbmO7+TJ/cYEGQEAECBJfIDPGJyT/x3gEyAFSZ0AFpGgFBuIzP0dSm0h5EPTJ54PitrKTvgF+UEdKAMRnDwu21YSH7mNs915m3BNdwPiMV95spPGakDckJmttkn9yFbztsKWpvE2cQRUMLyol6cp04WiooyAsIAFJEP+UFKlFz7+DG3/7eQBxNh8uc+nm1tSrl6aHN9FseFLwF0KxVZMTqQRLuH03Zz3iu9MPT8y6pe1KwlAsddGpSiuKdc8nrK5aDLSxI5ZMStUpwklajc9pJQm3T73Tf1BJWS720aqCYHv9hIgicXvMaOihcEztu9v5lOT4dul5T2NR09pR+ge3crWZ86Tdr5TWPPEn7FSEDAG4B+dP1blCDp6HP0DcA9QCELdcN7Ls8HpAXoRedJ9AHsE332bODkmlqRW7kOkEj/B0wFYMUeAQjb6tmP6TuAJn13S9klAxI4JM/lfuquqLnkCZEWAO/X1tJYe2d7L1C6Tg2w79FS/12UW5ssx8tIC4Ll7/idA+mxS2vefpEVgMhOK/RfPxm5939+Oh1bswLn7wJWg9uBjbxheLD7ronpOu1GQs7rBamM8MBe8p22Ro7Uj/8htPF+wHYhdyOzsHfmTcY96MaqgHFnPwvaCTCecCXfStsoQTywwhn7e7PSNymhY7QtuvX3SthjgH4IDEBwCLpmJxQU9UUXdsipYlSeFZcrQNRuz/e6Zc1DhZCJIrksCeAb9krBJq1kVjm9Pb6fkRalXVU3/RfX+dM/+vUEMgGbzfhG37F66msGhqNLGTGwQr/hGjssvBJlpy+Ytx/5Ma5baEL6CM8khBLtad6E5IPucgCc/q0SfQ+5IF9+g/RBjuRP21if3IgnAHpDHhArEPt8JxkZAInCewJ5oxsWBqpTtDU/0EHqhm5wL2M+pAO6RX7YCtrtbGQLv+NNgg6iK/RZiA7uwf5QX+pPWK/1elbkC867AnmZ94+Rmrzn0E70AeTDpsUF8Ltmk5+/C7SXBZnRPoDvf6fEOPL6/BPA7MOm13fwodIPKlJU79WvjGa7BtJGUE4ngpI2Y/fdVnkkqL9EfYSEEinA+y5k3/KD59C3LIRgngTYaKXIxzx2LUSTvQOTF3pE32Ds5Ln9Iiem9OZciVvhif1f8qYXJrqevvLW9vGw6ZL5SW9I9bt1+lhrKGor69N3CrdyYnt/W4mxkHHWCOjCq2KjrVdcX0igkEAhgYtYAgVhcRE3flH1QgKFBAoJrCKBX9T531cCkAF8AAxnwsPEvOFm7/dcc/+467p8m7wsAHQ4z8Scyfv7lQAXmFQzYeE7nhZMlgy4AJQAHOA+C5kEgAKYApgIWMRkCvCAlYxcz2HX8h2SgWv4BKQi8Z1rKLNNwMjXQkcB2lMO/mdSZUCYAVpMpGx1GMAAXgtMJvluz7ey2MpS/gf0AFQgVAfn+U5eJABLwIcsHE+nnLY/Rp6A6TxiiZCx55AXZeIeZIxMAZKQNYAO4BwrgZEbbQF5cbW8Ku52X//BUy6egTDiYGJtZd6n74AhyJu2Lo6LRAKKSZ+2nQ9A+dI5r9Tf8IJy3SuND7lmUkuSK1PP6w1c0p22wpori6wQeKf49Yl6VaPZisJYKIYIDE9kRbf+VIeCuPWttejwft8fHxns8scjb/7Lc97Jj46num9pw2T6AeQiQKiRY+sFMW2VPGVBhzPSRYk+DojLeVZwAhRiU6wvAsrQ57ALgJG2OhzQhGsAHDNSVUAv/clWaa8IqK+xYTA2BztFP8ReYPsAsrFjdyphb3g+YBBga3plvHCk7fmb1AY7+l18QHuBHO1N421b0jA95lc8eVh0V1zaNedK17ZT7+pIwTn2BT2PN72APLAHdiCfksI/ee94Ovnj97/AByByWyvuee+83PvN/Q3vTYLYng1omnvEur/SztTPNnodqZQD5Ml5ynlWoAoZLwPdDSwHRAegRYbYPeQJmUCbQzawFwNtSQIYw25j022z7bV0DfnQ/hC9lJfV9tlKaCWAeDwvOGehxigP+sfqfEh97of8YrzkyHQoihO/FMiRCQ+LNK3Ii0nbxiRVbcw7p140L8ZC3IQb9GIvG+O0yb3GB0+frqIfgpGyW3hhn9f66lxKPdEp6g5hYuSDkdnmfdh5/Gkf/IbsIXXQT/6nnNgAiBbKjTyRHf/TP6gn8luN6GEcQc6fUaKtKRd9kz6O5xKyw/uA68ib562XqKJ8jKOMz3zy/oC+kxf91kI7IpNVN/jWbyseHYKKtoZcwlMLTwvak3pjT3geMr5PCd3KHyZLxmQAZmSKzuCVg4yxM5QLQgRbt5berVZMzlPnLykxVhNejncwxn5k/r1K/1YJuT/YOX8uzzpbOYrfVpYA7QPBCY5CW78tfxn4fRK5Vx5+pOTGxwLXtzn5kIiKR+fHvfaWK5JUG2yXWgvtJA7Dk15QsgU2Kz3JFvPQ58+FsLD3ZbMVfOYJi2wMS+IImyIjFIzEYXM8ardkz712c6559VOfT/oPPFjrTpP0OjbQlg2TVwW5nNG1IVKZPyAbSEz0mCub8lAp9LToUYUECgkUEigksCEJFITFhsRVXFxIoJBAIYELXwJacd+WlwWTse9XApAA1ACAW5w8NY9UXTTRcg1Bkl1X+iItbAUtAAKTeSY9rDi0kEcGHtrKLiYtjD+A7fYbEybADT45BwjETAiwnzJwTz5MEgABQA+/mwcHkyILrcRvrOwC1DcAjfzMo4L7+Z97+A45YqQLdQAcAbACeAG4IB+upxyU0+4H/GDFpa0M5XfqYOQA+Zq3hJU5P2mzSaMRFBaqg7IAHHEv5YeIoP7IGHCIZyI/ykIZAG4XQ2Ml0Wfcod+7TQF7Pt45Rx0N/KNOADNMfj9IW+uzOC5QCeQAYHSyP3beFoHhc0p1Kd72WprM+C6Z1Sr+zWngSjrXrxWf2n7AE3fhRbopaodRv1/yWwLVFaUo9cPYddWipF2q+jta7fhkV82bvq7Hm0nb9QObenqqYy2PfRhsxTH6BpFAKJPRjv4CatO/TjvyXha5H+gX6DqkIfoPgEefAHzFvpA3yTw4ADkBU9knBkIOG2Cr4gF9WU3N/dgH7icfAFZAFWLNrwiqr1I2AHbKRz48lz5IGclvtPNc/gfQwnYSZz+UlwT3+CIrWnG5PFHxEjZXTse9yo5qmgwNJeFMK/UvlcdF0O0n5QmfPUTS0Xrq7ZJHzOff9P6nHntxNN3seFoYSVA91HTeB0+kf/f9Wz0AdtcduG++tsfd/uCh2U9qg+71Asbc+mwPs612/4ljp+awO9isPPG83vwps4VRYTzCFiNH5Ey9yZdPbLN5/CFvSCN7JuNDnuA549mdkGDscQBwyAp+8+oAvIYYYayiLNhggO2XK2Fr0S/AOSORzYOEvubHsXg+zxtU6lHwL7g+eVZkY0xvFCXqX/Q3L8B5qeT7XXpANU7TcYVlOy4Pp77hsuuWp0z7Z55IIZepNwQ/BArfGY9Z2Y3nDSvtV9JbZIHczRsQ/Uc2lI862f4ejJmEauG6LBSM0lrAIr9T7492ykHZAPCREyA+IDt9lusoG/1zLR20MZR2hhCiX9HW5M1BW/I/OrGuMFCd+0776JAWtDXkKW2MNwT2Ck8a6g7JCQl2b+45WZ/tlAmiADnhYcFYarqBnhkxiv6tVd+VimfnTPeRHfaMtqZs2D/Kgmy/XQmylbLw7HN53tnKUvy2sgTQR3RkTAkb9D35y8DxtQe1W5hULKjJ4Lv124t0bmpu3D+hlhoMKt6uge1pVznIPJWWH/RJ9I2x77Rs9Y+9Y9LejFn0cWyCveeu1l7oTZ70wBbZwhqFqUq7o3azK9Hu4eWunsdEVoy0F+a8sLlQSZL4cm2kfXmTGi+tH1qJq8iIQEg7ysUnNiIjLguyYrVmKc4XEigkUEigkMDZJFAQFoV+FBIoJFBIoJDAShL4kE4ygQfsY3WrhfSIXdBVdq2jI6400OUSzZPTqrZ3DWzy8wpdC1gIIMBECrABUJ3JlIV5YqLFhBtAndWNRhxYHHJ+A5DgAFThd1sRxjmbmNvKYYAY854AbGBCx/MBUCgLz6YsTOptM28jCgBAIAZGlVjFyKQOgIiVYYAuTATJO+8dQh4W+ooyMJYywbRNrS1kEysuzTMCoMjGXGS5/LDyWF3N4wTgg8mf1WlM31+pBHiB7ABaaCPqNqJdHwM395Wb3NO/Tnle06kPk9IsnroSbUl+gHK0cXFcPBJIu9N4WkD50VmvNNaXRj3ytjgiduGwQj91+UnSUkiiZrmkdeHSNwEYPVJuRbHx0lJQKpUDjz5ZU2ibpFIptZWGBGT0tqO40ddTqdUbYbK96pqvGfLivzqWPqZeagCkgW/0J1YjA2gCtJ5Blq0Q1oZ+i34Teob8AEDoe8TIByyEEIGUALgDTuEa66vcC0AD4AfIDNGHLcA2AKzQT8mLe25XYoU5oDTn1gv+AVBSJ/IGRMZ2UR5WmgN2m12iHxtZkYULGi6lw4EfDQm4vkyrVuf7XbsU+d4l8nTZ1ND+QAtecOkurz2/zYX7J73S1pNeeUuY+jufKvf99bhfeVLER/SuRYAU2zimSh8XYXGH9j/YNVDK9nIQYO4+0SlTPlwTPz0XB+Uw0Jb8G6+//Wr3sXueNNB6pT041ioH7WD7oWDT0CFkjX3Eu4Fzn+983tKRBYDymBI6Yl4Paz2H33kW9hybyjOwr3jiYO85x7PMuwBAnfGFUFAAc9HSXiiHZg3c7lUn2qb+s1NEXyh6v1teF/0iKLp0rttz3oRIQXlTOD/1FJov1c4xaXq5ro20ejn25bV0c1+mi4yfjEmMT9Qb+w/Rhl1H/wHc84cR43gPcECycB/XcpAnnj/IFU8LgHv0nuesh6ywZ/F8xpJ/UsKbhXKh7xaOjbxpe8bQverbAOurESFmK2g75E1ZWShA/6XvAgijW5STcp8T0a62gqDCDpmHKDaG8vEugBcDxCbPhSjjefRZ6kV6lRJjO32dMZ97kC99Hj0Z69yjj/Uf5sW1zAZST0gxI+DYx4L25hl8x/MHnXxS99kijzMeuoaH2PoLWVyZlwC6jM7Q7r+sxHhzWngoLs45IECOXYJ3AkcSJ19S39cYJOufauxK07rcq9Bz9oKACZ+Tr8O1+mdan+i+EYK2yKau6x6SDRnUNdtlvBr6znhAn1FZUumNxzPRzZXwHq1TSEPlHYpMfSqO2tOtuenbRFBc5qbH98Rh63lyAVHpKLCtzzmrAnxEv0LW8+6MXaRfYFNsEU6hPYUECgkUEigkUEhgwxIoCIsNi6y4oZBAIYFCAhe+BLTyviEvC+J0v1kJoBvwgMlx5OYfCV3j6cMuaVzmSpt6XVDShCSwDa8BNZlQM3kbVQIEYsJkQAiAhq1YBeD4rJLtM0FICYC1DNBTAlhh8sX/5oGQBxKZSZlnBPkDRjKxJz/KDMgzpgQYyXkmc1zHBMpCQjHZB2xh5SL3cw3kAvUAiAJAMQ8Pns311MdWE3OOSSv38FzqZuCGkQwGNOmn7FipLlYvI2YoJ+Asz+H5tAUAHUCkPRv5UEbKT/0eUqguzz36ZsoOmMvKbspPeZAHMbWZ9AIGfZg2tgIVnxeFBBQgPxgVKbG14fnDfalr6P++ibS8WQo5oxBEcwI8hqWAgVZ694i2SNPYhbGnOEVxXE79YLDZjkVguL6FRrrNecmUYkdsLvvejiAIJocHy/2K1d/c3eWi33uef/TXnk4mJsMMaESn0T/6BoCebVBPPzjb6nd+h7B8qRIhWOgH6DtAyCc7em0hZ1h5vnyVuYWRAbQGvOZZ9AXASfoW/RiyAZITe0VfAaAEbCHfsx4d7wqAbfoaXmjUk7wgLigL/d+8yhYB7b9+IAsr01UrVwUWDQi43q1QQKOlst8oJ2mXkKstFd/vaWt703qSNGfSYEczSbds85PHU5eE5SSeFOG0NayUTz0e907JQ8ZretoBYxHMnjzScs9/+97k479zlb9Tsb04x/Hb8rL4D/Ky2Ah4v1b1V/qd9qJ9AXU5kC0r95GDeR88m3ypH+0xpoStQ8YQrgDhPIO2hZimbRk/aEvqyjWrgrirFISyYnvJ59NK6Bs6zDnyZ0zBzgN0QwSgy8ufgRzYmFaEHvHUnDbYToeTJBkRNEk4tUqlXNqk0FCT2sdCq5fTQDvZq9n9UIRGb1e1pOd587pnXHlMaU+M9usfUsMLO1S+AIKQKJQBosE8hWyFva3KhiwD0LY+xjg5pgS5T19k7OAaDkgAC9u0KlG3CqBO3ZEz8qANzOuAciE36/cmU/rd8n5KmWlL2pY+SBhDxihIGd4D+A0yku+U87x4E6g+TfVhyEVIfMZF6oJcqQPn+ETX6NvoNCQF+m0g7Ji+Q2pRHt6PkANgLXVFjuslPXXpqgf6iL2jvZAPtoUyI1/OISNbLEIZIGfPIIVW8xA724OL39YlAbNttAnh+JA/epp5uZ21YaPwZ6eP7nfdgyNRudaTBpXaJrWc1gCETfX9TSIKTpa0DiBN4lIchXNBudLy/UB8dtzWuCv7lAbaCWdX2Kqf4Nokah+u9g4pmlPABt8iROJD2A+RIJcqwlyfPs1TaalYPEzjUNKcm7ytMTupra0i3QdJkco25NX3DFWG7IMQxQYyZnJAXPIejR1AF8/F5q8lvuL3QgKFBAoJFBK4SCRQEBYXSUMX1SwkUEigkMBGJSBA+wsiLVhJyoQY4M1WGva6qfsE+701dtFkmoWEinoPu1KNST+gIgAjIAiTOYAGgAsADSMemIAz+WZiA4DCb4Dp/M9vgIA8b1TJJv6AHHa/zZ6MCGEsAzQA+ACs5zr+v18Jjw8AD64BLKGMFsKJ8hkJQT25h3Ncx+pJwAGu5yBvykk+ABKAFtzL6l5WsVFeQA2IEMrK9Ryco5zkS7n4tO+dS7IP8jKihUkvgAQTPhLlQTZ8J19kDFgFgEJdmIjOuMahGTemNdfNY0a4sMJ1cd+RxWQg3uO0bf7hxfeLQgI1Rc2/WmGHtBrTe7EwjcrOpHlMqzxntMrymHwptisWVKhYNV0CLLqjKC1Xy8G4tHlGoAYxhUrasDsVsKqANs5vt4Ww10rVStkfETByqlTyu7VSlH7R0srw5GM3+fVbH0jG9D+gKWDeqBJ9B1CSfs9v6PRqq66NaKNfsMoY0sIAWvoBOkxfW4mssAa1/kZ/wbbQX75NCZtEv6Tf0afpH/R/yoY3B7HhsSUrgo4CAA1kxW6wsp/6AGZTT9trg/8BdMh7qY79PZWKTGZFIYN6Ja9+5KaQQJcI0B6Ut8tWbbxc0Y9TXc6bFrg9OOm82hYtsN3iRaciLcN/JAluk7dFV9o9+EXtuI1tA0TFPhCW6tpHZKXefST9o//9Uu+3OkL4YX1uF2nxfSItANifq4O2/Vul3+g84LX6fHen7hmBI6+QFZ+t8FbZ+bOsBGdTafIn/JHt4UN7QmhhL6k77QfQbYD4RskKK5t5WpAvZAg6wTiA/ad98c5Bp1cDptN2GEfqV/w+K0JiQUzEUBD4zXLFn1G7D7ZCEYAKr9ZohJEIK/rWdLXiL6h7ZV5BcZJW9YChUsljPGmO1rzWZJhSN1tlDVjNuABhQzk1IGdjrRHuLAxAPoQ2Yizjfzwa0XmIDMYlvCMg5+Yl99X6oMnkbJ/Im2ez+IB2QP8hSMiT34yUpKwQLoCa1q/oe9wDQUBd6cv0d8qLNw39jBXsjF0Q8Cvai3PwIKCNIKUAXy3UGJ8c2ArISGTNmEub06eRG2UkjByLIWgTQok9F+WjHMiKctJ3eQYyoc8jK2TNIgaIE/TjHzvl7VSh+DifElBYo5Wyy9pHG3Jj3LA5vNvy7vm7az07bjddc3ZKhES0qVxVE2M06vPdrAqIw/YLu/qH2dyGTSXacbulIIFBoJBNXX65EmkjjKn69Pjudn32ShEWx3XRTpEOR/xS+SMav48kUesWkSBbu/o3eaVKV6tU6+7WOJ29l4qjyFw/5FHRLcLDNeemRFKoq+qcyBLzOlqt+Izx1PVuJSP68K5gPOa3wqtirYYvfi8kUEigkEAhgXVLoCAs1i2q4sJCAoUECglclBIAuAO4B3RjsgzYUXPVrQ1X6qm4eC50YdJUNG6tRKwxGQKkAIAAwGC1IWGlbBKTxXFXAphgwm9x35ngAQ4ARjHhIw9Wf3Id+QC68918060heB7gAiAP4KKFJAFcANgAlOHTVlZbKBHLx0gOxkLAHa4HGADgIS+L9wvoYpMwng1oxT2AkQAFrNgmbw4LB8IzyIOycQC+GkjDNfm62HcLHwP4CIBD+bgfgOxHlJADiXxHO78DVgEAfUWboX+PO/aXTCSNoLH7qReypY7IlzYtjotLAuhMSRv/NkRWPN1y3i7Fghi4MmnulWLu9b2kJ0mTRitOw0olwNMC5GJAIGs91KrLME42+ZGnyFB+VKuW1Bc87c2d9kiRg6m5xvjEXHNmU19tqqe7Ml0pd9HnnMgKA9osvBn9ir6EPaHPf7Gj2wBxy4kB+ojZC/QfYMRCrAFS8xuALfdlYOsaoGXcCUkDGPMpJby56FvcT58iD8oEGE5/5n/6yRleSB2yAnuFDcA+UV/ywLOM86x65jf6IitvTwODq2KB5FnhK85WWeGByuWyX1bUjU3ainVIREa39qsAdNbPXjziJwtdYjOqXrAz9Esj43Gppo0vZkNtkbDglSfEHmkT9AwEBkTNQunEqQvvmEg/95M7vV/UPhb/DdnoeJ3Sd4m0eO9zuJ8FsmTlrR3YHV9hoWI9c/mq+txl6/5K/thhyCfzZgMY57yF6DPyelWyad1PeyZEFPYeXcu3o5HdK2WXarPxSCQFes2G6k/q+6xGhh2+528TmBjWm2EibHILLhUKrVaqlYMuEYHyx5BTU5JWoiQekIsGet4rQmv2hfr21bmsnpDj6Bt5W4iz1+i7AfqQ1fQVPAMAtCk7YxQy4zv6CvnHggLy4P8Ntc0q/SxRv2BV9R1KEOWMnZCClIX+AClA2zCum6cPeo5NuFTpaiXGK1ZpZ5HyO+VkLKf/o+Nn9KXOdc/6I7efxb3KBF1CNoynjNeUf1Tpu5R4l/lYp5zYJgtVxZgNOJ3ZPB0rEpwbKeBZ5Ist4p0Dzw8IFvY+oHzm9YNseW+gD5pH60YeXVx7DhIQmdEQafFlZYHO8g73a0qEFYMgX/EQOeDazQUHaQCXIC8KbUGmkVkkhQhs+dQpaKPOaSzmXVlrg0q4YMixLr5e+01MJGGo/qWhGt1VXrr3Ktdq/J/2MG2ineUnzwxXGxh2Ii50WSxShEhUi+oaNuadPCgXc1mMX3WGJ0YnP94d6Z9GmtEf6LPoPn2U70X4p3PQoeLWQgKFBAoJFBI4UwIFYVFoRSGBQgKFBAoJrCoBrcT/urwsAPB+QgngA+DmK27m88Nu8OW+K28RaRH1ubJXce0Zbdvbd0qzI8AjJmxcDyABuGikA5MbgA1mRoBOXAeYDsjBhJuJNtcQT95CMXE/IIGtgAR8JZEH5/nkOYBIBmYyqeKZ3AsICcDApI9JPyAD5znH88gLsJK8SAApFtJFX5c26eU5JIAMJmeAMIAcPNPKwX1GWnAv+ZuHBf/zGxM/88DgnH03Dw8AHluVDcDKCkryoMwcgJPIaNGLJU18N/ZfvsPt+w2ACurB5BEQiAPwhe/Il3q/mzbt/FZ8XDwSyMgDbbp9RJ2kLlikGnr+8wbT8OiWpB2XnMJO+PKycN5lXuJFwk4i3VCO47grjBIt+FcAqLJrVjxtFZq6mgiMCYEt1XqrHcRRmlRqpVJ3rZwM9Xehy+ZJZNJF3wGasR30ecBJ+hCeWLb3xHKgzzwYAGCxC/Rt814CVASMXSIr1tOMuc2V6T8A2uSNbaMv8R0g1UhOyggZCBho/d422Ybo4Hr6MjYFO0DfzJeJ+wBZzRNrqYhaPOsLhO5rtKJdvqfY46k3GCdxjx4Sa/flGclVq2jjQWFW/dpbpNlbVqig1A0Lzu5SpKiZwVJ6bCZOb2w6f6DiuYNll4zPCenWA8yzrH9GONX7T6R/8mM7vLYK+T86D2fFLyAT9XouDsoAqWSHEcJORIkTaXE+nmltgayZw6BP2FwDyoxI2DBwfDbvDuVvgPSadVA9E9U30h4VC+IjZpM4nRdJ0ZAWVRaaYU8sNkIkRlDSMupyOQgrbKnuvO4wjEJ5W2j/isybSTFivJo0LCPNf3yHl8hrxhYNQDwwtkH8QVpATrAwANuPRwBjIeMGYyB6bqGCOIc+0v6QApluLu29sWbN1rwAmbPKn7Zh7IaQZLNhQHTKxHn6PYse8Eyi/0Ca4AVCXXgXYDw1shJ7Qb/ifcL67Gnteg6eFUuVwbukQ7bQNxivsQHICrlyUB7GUMpI+fD8YAzlvYU+Tp25/jRPKm48H+VbKugzxBz2D89R21uLcmJHH1XCLnGe7/SNc/GcyT26+LpOCaA/9C/z2KMd2CsMLzzaCaLc3s0Ws1z0anApawRamAkdjL462iIbXFOWJPtv8RVzkWfI/pr376pFY/+JzDNDg0lj+pQIESIR8sq46GEh8gNPjkWPi9UPvIjpf7+jhL5Tfm6AxOPTxp1EpM2G7e7ZHlz8VkigkEAhgUIChQQKwqLQgUIChQQKCRQSOKsEBHB/RqQF+1dYnOndbuGxOdc+2XQ9Vyv0fTrgWscmXGlwi3DPbm3C3aN9LQAcASNsBRYAC0H+g34AACAASURBVJM58mAlMKQAgAmftymxetL2wWAiBrpl8ZmNQCDPxbnbM2QF3zkHoET+HLim2wpcAEkADyaL9nxAIAO+zIvC8rVV15avgSfmzQFxwGQUgAzgxUAVI0+YvPEcxle7h7zMw8KIFyM4rC58mqcFYCcgCHkS+gFgl/yM9AE0YVVnt4um2m5hT8Ud+j2AUwgLwrB8IpPCojypN2UG5Lqftuz8VnxcXBIw3UoUFqohbIRNnUcO+V1HFSJq0EvTpkiMBSll2BZJIUqtRyvAA3ld9CnOfiC8oylEpSWoo9kKE0JLtASy1Nth1OrpKrf6usuTWtkft0SJVCvB8lWW6DHePQBp2BEOADYAPwtzthwxoe+gu4SBAtykD3M/egw4uJGNsU9r6c6qasBTQFs+6U98B/ClH1mole/U97s7/88I1OSZZr/M2wk7ZQTkqL5TbvouYPFKsfZTea2URAL1yc1CK2WzPq19zv243fb6oiipycOFsFtZeCC/7HcLu/K8OKoOurge+pWuIIivqntBayJKa1EQUNagGbkgTDN5Qbog24k/FcD973Z479V3CM8f6tTtPwtMf8dzuJ8FJKod2HHb7+e0Nng2/ywDf42ksHBDzybL5/Ie8UupfCf83nLZ6w4Cb1j4YHel5NqhNtqWkrTCMJ5WaCjFpdehxtYKaxEW8nWK5bHoubruMfAP289YSV8BDEXP0FkDCjnHb4x1FlaJz8VQgYv9BSJpN3rRSc1zDAO1muxoFwPKGePuUkIP8AiArOB3vDDw+CD0GnUh5BYH4xdlpS4QHGNKhF0CoCfPJeJwtYc/2/OSBR5Y1u8hLHgP4H/AWuRqIa4Y26kDRBEgLmVE/hA//xrkADLgeX+jhLfFG5R4P2KfDfo/hBU2EhvEe4q9Ez1b0RT3bVwCtBFjBaQWuktfJFQXxNwHOp+0G+MaB223ubNx9plPg8zIzj47LiAjKOJscwwXtXCOXHwEJIl5WSx7KOHlsC2Mh5DdhGRD/7FB3M3/6Lot6kHH0lXCZZ1Zn+JMIYFCAoUECgkUEtiABArCYgPCKi4tJFBIoJDAxSoBAd3/XaQF4AckAgDDdjd9Z811X9Pvqls87dSnhb7z8j2vKFQM4LomQ0HZ9k0wsN08CSysEZN+QHUAP4BCA/gBoZjkMTkCOADE4DoDLIxcsNW0/M8Ey4gIVkKywpODa7iXSRWAJwf5mIeGNanlbSvG8r9byAwDYm0FOfUC3DDygXutDnliJe9NQR5GXhjJwbXUEbARQJSJIeUn/AfhH5AXz0JOgCiAETtcrFgCM/cHbuy3j7pwjgny/8fem0BZclxl/pGZb629q/d9kdRaWrKEF9nGliXvC2AMGGzP+A+MwSwezP73DIMZYzDMYTHDMoxhjMGMDcYYkC28yatkSba8SrJ2tVq9b9XVtdfbX+Z8v6x3S6+qX/Vare5WR5wT572XLzMy4saNyIzvi3uvubxiBygLTIANdsSxc3WH+vCD1lj/edFJAB1Dn14tJxOJYiGsawgHfzjqmexP6ke6ms26dl2uSgI3GcUC4UKnuNuJcPJkOhI7gR8J+d4/VKk1igoQ7fLZzKTwjl0C3YfrdTcuFzeTIjYa5UqttmH1AC6A5qMrdQGC6CEEBOMQsI9x8SJlgB1zKUHHGKmHPlNnxgPgnIFvgJeMl9NDcCiQANgaT6oT1hG3t+4BccocB7lC4F/GIrvDGUP432eMmSs7xhdWYIDAEIxYMgHAMob5zjg9Zlf+ZRuXBgKq5VtL8UCEUtdqTRmrJF2SPXOUAqrGPa6pPwRoi/Mta2d+b9xoysOQq+WjsFomiqrGdk0zjbwHNYRpb9QhBXBO5zjmH4gXwGl21vOb+r5LGcKC9AvKVZEW71QfIdfFTsjTEruKL9Z1Riy3XzzHRtTfB2Q1sUXxKHKKiFuW1UVeWRY0QaaQy4zI9VdFG54zIihG9b1eqic1jb1GNiuiUE/W9Gnx5DPG4nSgX+zWBjxETxkbAP7M/YD9jB12QDPOGG/0C3rMdfFZBtcZW+ifWTcybjYqQ1wAplsMEJ5tWE+Z6zezVOS9gXoz5hmPzBuLaQmSCrRDYrxyL8b/LmU2PmCxwPsEpAAALv/h9ocNFsgeAsjeQxYqd7GPcz/68zZl5iFIYCxskDFu6NAF5iJIU2TtSYvF7oETl8cYMFLVNspAvkHgEksGIgASj/N4b31jq0g2nJh70RPf5VTOSIkPIynSccWzgffX/9OqB/pi76LUi3kDchEdJzE+eAclt2+4OZVa+HO9BLwEvAS8BLwETkkCF+tC4pSE5E/2EvAS8BLwEkglwOLlfyizU3LYDd/6mMuurLsVr+922UERC711V9oRuq4NsjUvTrpoKcAJix1APRZqFp8CgMKIBEBLAA0WToAc5rKJ/8kANIAFLJAA2IyU4LeRC9TNdpDbgsrAfcB+wH8LYg38027t0E4aUAb3MB++LNA414IQ2iKNZyfgCgtS6sa9aJ8BqEZQcNzIjfb62mLWSBF+c1/aigyw2mBXNP8jD+7HJ//ZjvR9rry96g59WMTR7Vh6sNgE3DW3UgAaLJSRPfL+S2WfLl4JoEOMR8BsdGNUhEV1KsiEh8L8xOZmuS6QdEjg94TcQU0pyoI2+8clgarNbBRNC+jYKNRcFIYojTipNhrNWk8xd0Asx4i2iitot+JaJEH5sd3DjR+8XuO/c0If2f0PIMNYgwSgXnwHCGR3vpGJzAcAcYwh9BcgHoKAHcRmvXDGvdlmbUG8CsY9Y8yCOpsLHnaDIzfGGSAwQCtzCmMeopU2cJw5hnpy/jGxL6js1k3Lkv2HJ6pyByXDiUQeP+JqUw47Gs0UeBQgGhSqjTRgczObzdSbMrzQLv1pkRrajJ8oJndjPGgGo7kws3wq1Pb9KCiONwNAX2QFkUx9mHOZd4KWeyLkxY7eT7YE9mv6/EdlAgUvdmqPh0C/tf9e7Hudz+U11W+K/xJX1c+Km+52qw+XyGJJRIYUPghWiKDIBiKrRGh0ZURN6HcPf0WROyQXbM3UjZQCWaiR7eOJ7+gWuoqe8txAZwEXGVeQ1DwHbExBnmGll7otWkT3TyeSvT27Gb/sKseXP4A/CeKCdgH68+y/XtliPXEOY41nH22jjfMttk507zP5vx1ktrgovHMwd/LMh9Bg3CBn5qynsm7t7UKu1I/+fUFLpox7dOPNrfp9Xp/muifdBX8mgvHXnlgCC1gZpO+Vim9BH9h7oLlN5f0RCx4s4TgPMsPehYk7xH9fUWZev1EZIu8lrU+Ov6JVJu99EGskLBd5ttp76D/pO++UjDOut3dljqHDEJ18N5Ib8ptnGLrOuy+6Nt+CwutSS9j+w0vAS8BLwEvg7ErAExZnV76+dC8BLwEvgaeNBLRD/5CsLN6nBgF4sZAqual7l7j+5+MaSl7vx/Mu0zXtqiN5l1++1dWPitBYCvhgLpRYKAHysUhjgQRwAbDGs8iCZpuLJuTG4s7ICrO2sAUfC6aZvaczycB/7oFrBFwmbWqVzTXsKAMMab/GiAM7xm/qZ4l6AUgYUEHdaEu6O7t1T6sXi0wrh2Nm9WELO37bAtK+89sWj2nAXGXuwS5ZiAlATOoAOEL5tAGw+TFX2XWp2/HOXjd8C/Vjhzc7wdnxCagKgMkx5Mui83303Wyr/JeLUQLmqix1p6Tg22mg67riKQyF+fpYmBnqb9blOyIZ0O5vKXgwoA2Zykm+KT/a2u2fU0xgYevuiP7H0f60DDSy+r9eF+gu0LUyHlea73zzc44HZADY4CKDMcS8QB0A2hnj5u4MkNLcQQESAuyYdQifAJgGYs7245n4im/5sGecAPAx3hg31AFSAuAH4J2YFtSVHdcW7waLDIuhwFjdpQxYtKC7KixPPvmtfQpZEY9q4JeiXKYnisOaC5qjArazANZyC5RVP3S5QEHN8eSRaF4Qep1RyPNBBT6IGoq8HTUPPZRkV8q9V3M6CdapspGuVUD1dP4yIDvtC+4piwraBtn8Gy2hfVPH1uq/xZ4XAKGRCfIgIbuLLrVk3siKbBLpN6nx8ShjqVptrsRTvQgKQmhH6lzcf4UaS6WmbJoixd2V6c2kOnNIHMaYvjO/2/PE5Mgx9JVnKHoKUbFJGaICABLwkp32uJrhuYo+lp5CssLqac9JrCo+ocyO8te36gsgSjsA3NEXLAT4Tlv5pH1c18mt2lOhT+115/nLc9lIFJ7ZpHNFVlj7mUex9uDdgXmKuYlnP+8rzLX8/2pl2gKh6i0tngrNWeAeIjNikRb2L7rDuOR5h/5DGjB3o2c8dxjTzM38Z4Q57smIC8MmFJ7n9PttysyxjBWeXfbeyTsw443jzAXch88NyjwfeNfk+Ytuk/kfPbH3UT5TokLZJy8BLwEvAS8BL4FzJgFPWJwz0fsbewl4CXgJXHgSEPD9DZEWH1TNX6nc56YeXunqIigm7s26ri0ZAWuKYSGEs7Jn2hU3rnUN1szRDpfJsZhmQcZOUBZbgCt8snBjwWV+r7kAsIvMggng3nZhs5gzsMB2nrZbNfCdxfpOZRZqtgAEYLSYEtyv3UWTkQZ8WuYedo4tLNkByg5GFozsVON/SATzad++E9asNszCop1kab+ftYXFIotSsyYxn/qUTxkkFrQPyg3USld6qMdNfTcWWcFubuTKeQC+LFApk+MWzPhW+qxVhv+4uCWAbkAUQARAaD0sRV09FORzR4L8yEZXHtd+7pVyed3dSJoCTN3jcRJcKsC8IIdQE7K+KDXj+CDRQcMkGBdRMVxrNI80Go2pWi2sVesN09XjSdkC/wJskyArAGdwH4T+M3YZL4xXxpa5iWFM3KtMEFPKWNTU8mGPOyfGOfVh/AAMmfs6s8qiHoCpjGMAIxJzFOASZKIRGAvWL5sNG/l8ZlKyHpUbrVqt2pRnoGQiSBT6PI77tNO+r15PcpVqo0CAbt1oQP6CKoVsBnS7VIvC8XocjdUbwVJ16Jj+F2/h9nOe4ogAROHKZrodoBaAXhNBwS5eIyyo/4/r2J/y3yIKk7kMoJxd36RNyuZSZBFvc0EUxXhDHw6qX3GhFhD7No6DvMLoTtbjeJn4iiArQkN8VEAMmDjjKiKm9suCaQwSQ+PTLHWCrz0nxGLGnnfps0MuzfjgHLOosxgQ6AGAKGPKrO7OldB4hqIXgOb/rgxoalZAzBm4foJYQW9wWWX1PteAKbImIz8bI+0bEM4HMBe5EXOAefMmZdtxzxzFrnyIVv47QIyOs+wK7Fzp1wVz33kWGEaK2XOzJkID3WdQY23Ic5DEXA05yTsg/c2zk3dhnkm84zIXmCWEvcPyXIV4t+ct52KhyPk2R6Tlq04XqxXcBaM3vqJeAl4CXgIXswQ8YXEx975vu5eAl4CXwGlIQAD4Z0RaACa+WHu097uxr464gRcVXHnvRpdbnnVZeSZpDGdd6YmaK26VC5lqvwtWDmrvqAXCZvEPeAHADpAB8AeRYb6jAVU5jqUBCywAQVu8GRlgnxynPCM1OBcAh52GLNiMKOF8/jOXUraTrF0C5n6G/8z/POWzgOQeu5RZOHIewKW5sWARaQHDU1csyiwCzddvu1srIynsvtSL8gFGIVYsUCYLT3MPxTmPuMZkzlV2dLmRLybu8XdASkBUIEcAaICeLyjjSorFKv9/mb5qb6D/flFKwAgAdBRdAxQB/JdJRbCjEgS7hsJcajmkHd/Cw7GuEHraDJph5PQziIW0duk/Bdp2h3QslsuoMQGs43GzeUhExpDIivIJrCtM8IwJ6gCYBqiKbv+AMsTEc5QZnwAq1Jk6UVd2gjLeICsAa06GGDmdjjZwEvKBecfIC8oizgb3xe2SubWiHVhUACQx3sylxpx7z7f+0E76hnbY16u1xrQIi0MCrVdoB35GHp4OBUnEvNoTRsmE/q8rAHdBhhVNSaNeaxDnollZks8deGZX8sRUJd69tx4m13QHD4uwqO2ruB5NOoC/NkfNlwH//Sflv2v98Uv6/DeRFjs6xBw5HflxDXLD8sQS8y9A2cWaGE+KUxERpH6ZxtJe9VVejtVCWV9kRPjlZLdUC8RWyfJCvEZ8KIoy1TBS0HWXTOIpSoJrJ9jn6xbBohkf6B/jycBNs2o00P+sg+snsHJKVE/GB+Q5zyzqh67TPp71WArYrm7aeNbrO18hT1T/eeefs/q1SCqrDvVArlil8A5FXBN26PPOwfzFp5EYt6Ir58DS5mId+6fc7hahMf8dkXLaSWUjABcsX8QHY4p3wtmNNCo70XEjKZ5y/T1lYfgLvAS8BLwEvAS8BCQBT1h4NfAS8BLwEvASOGUJCAj/hEgLgLEfc0c/tc0te9UGl1/br3CedTf25dgVtxRcmMmJrCjJ2qLPRV1aPAmTj7LsBAVoB8jCCsLcvkBmYJqOSyNAF8AMA1tYdFtgTkBCFuYsyvmf/4zM4Dv/bVImzgakAwCaWXFwHgAoxyyOhl2LDNrdRbFA5HoWfoCru5QBUtkdatYgtIX7GEHBvakTmUWn7cC2T9uxaQAUoI3F7DAXDuZCxYIK094HXGNqyFV3XukOfSTrdv8hu+9epwwxgd9i6gM580OtOgOu/rP6CBcCPnkJGDjBmEHf0B/IQXM3NvKdTH/zNTU25bqqUFN2PxO/YlwEhc6V26das5sIwNJ0eYNKIu0In9ZnSVlWAjGA2ckm6kL5fKLzzCHUiXEFWYFOM16xOIIIAITlPMZZR5/xZ+IOqkOlGbeMOcYU90ZmCMYIUcY64CpjnXYT1JaxWsNK42SEMDldTXLZTEpG5jKBgMZwtRw69Yj4mZYrKJGWcU82E9XlJyifzYW4DCJuiLxDJdVslMnms0G+L5uUX9ebPHRvOYgHs25oqBGURhWsudZI58NGJ1BSpERT5MTH9f+fKEOOMgf/gTJ+SjrG3DiZ9sw7h/nyvcq/3joOcWyWdKdR3AV/SUo45HPRlILWPyprJayY1om46NIAyErZ6kkYlzKZTDFuJpGsaw5JwSZEaI3qHAtyy2eyEKnU6msIAYSF/gJUWjrfgEkbX0YOzlpKLvI4vuAVZ6EGdJATMq2p/+/X583KBG5mruSdACKL9xfIC95DyjqPuep804unbX+di4ZBTrTuO6ef246fi2r5e3oJeAl4CXgJeAmcsgQ8YXHKIvMXeAl4CXgJeAkgAQBxkRYAeo+4R9/+I27rn28QUdHlCpvzLsxVXH246cI9ORcVQ1fdHbvMqgkXrQKQB1QDkLxEGdc0uIcCxMeyAj+7AH8EtmWxBbBmfrj5n8W5XcsCnIU4JARgJ0QEC3SO285UyjDf0xznOwAQ96AeHGN3IsAaxwBMAUgpi0/KZQcr98BVDPfjHCMaAFUhYMx1Fc9VrgGIsZ3gneJmmIsq2mZ+89lFzu5urC0AGagX98648Ts3uMP/WHAHPwTYjLsVQFL+4160md/I9l+Vd3uyQlLwqV0CZvGDTjOO2IkLwomeQ7xVZCHB2Ep3Ob/nw9+Ux5p4WjvDD8sCIA+4qqjPWWHnwlED7QgPa7IUqIusYBw0WteerMSpC/e22DWMASwsGCfoPnWC1IAw4LjFwbFxdbL3Od3zzFUHoB/1ZM6gnRCAxOAAlKeuzB+MQSMoT+p+b7hhS/yJb+ypTk3XRjPZzCHJ+TFZrFwSKV6BCIoDIoyqsmjprVTqFQVtLmai9P6NfDaazuWzB+Wea1c+dMO9uXDihnwwsb0SlK7ucbWre4La/3puf6fdue31Yq54mbJZPfywvr9GmXljMRL69c/KRljg6stiAS1G+RdaGSmYTI5kVaMg2xBdcuGl4PZ6vuUzUUVc1G4Nqu4kCHsU8P6AyArOhzBDz8g8W07Ur64FZJ+3QHQb0N4Opp639b3QFK2lZ8TuYm66VJl3iNuUr1Q2l0HMp8xpZkF6ATbTV9lLwEvAS8BLwEvAS+BikcCCZsYXiwB8O70EvAS8BLwEzkgCLJAB5+90j/3it1196ICLy2XXnBxz+TXaGVwpuCAOXWV/5BpHiq42YQG3AecBZvC/bHElANOID/FsZYBBdgwC2EAWQBQAGhpIb26auHcKArXqAQFhFhR8WhwMwE6AUcoADOW+5hoHNy+cazuBuRfgP+WSqDP+7LEGIeGaxsqiftSB/7iGbLtGKbM9iLf5FzZ/+LQBAMHcOlBXAFtICzLubw66Ax+cdA+9ZUpkBW2jLhuVuXZ/65PzkMudrXvTJz5d5BJocx1iVkS7JBL8xOOW5faWLgFqmZ7PSkwEBOOpXqs3y41GPKnd4ezaPiKLimG+K77CpNgKxs+pkhV2DwAzxgH6zxihLOYDxiYZoNsCcVMX3Bmh43OsGJ6CXdnmpsZct0EiYhnGmDus+1dblhWnBLz+4PUb6lPl+sjUdHWnOudbhVwW4na4XK3vr1Tre+r1xrAsKiYk64Nd+cy+nmKulM9mRmWR8XAhnxvTTvwJWWHUBvNh8tz+IPwpTbVkWVAck9uHgXbp0x7cgf1u2/F/0XWQrouVsIaxZHPeYpV9wZTTsohIx5FyOgZF+I0p48IL11B7Mplwj0jBQyKopuhTWTFxPuPCnlvnKuj0BSNnX9E5EoDowsLyYWU2U9hvIzEgqtfp2eDX/15xvAS8BLwEvAS8BLwEznsJeAuL876LfAW9BLwEvATOXwloJ/+YrCw+ohq+XbnkHnrrV93lf/5yQfAl1z8YuGiJAnFXCy63YsrFdXnr3i/AvXyJyyzdL5dRgP03KbPDG0AH39YssgEmsbpYqQzASqwLdggCbuI6hnP4z0BPAE52YZMAPwEPjSwAAOK3uYfCQoH/AB5Z2BOUcmvr/maN0Q4+QhDgEgZLD77jRsViRgD2UiezqmhVYZawsB3rgAPmNirdLa3MJy4b2MUNYMy5EDb8hlQZcXGj4A797WXusXcccc1xAAh2nENW0H7ICgBdC6pq/vM/Qp9YRRbjU77XtSE40Ic8r8+NJTK/ve23M9Km3eWWucSaUy2VvRjV9GUsLAGTO7rFWGJMMF4gCXYqt7uQaS+F6zjXSAI6Cr3leLrj+yTjVixUM3SXsfgVZeqGlRMWVoxtdgUzNnG5tEvZCMJTIgZORSlO0od9R7dPp0OcDPYX41w2GpcVBYYr9/X0ZteVKrWVlVpcyeejw91BsEHWLYX+3sJwtdrINeJkMpfJHMjlw6FiLjcmR1HMn/SDWc+clGwgLURQ/F5Lvj/WktF1OgaJNVuGzjsV8TnOVxlcD6FjCQKXPl4sl1OnVKdzfTKkRUsmFtuIPqO/IOd4jlTV+WaFYf0IyMwcftLWFee6nf7+540E0CXecewdCmvMLyrz7sAYxIUk7x28P7THRThvGuAr4iXgJeAl4CXgJeAl4CVgEvCEhdcFLwEvAS+Bi1ACAp9nd9gJMD6hu4njiahFWvyxzvlvwmKybsdv7nBrf6rhamtrLuzpV7DoaddzVa+bfnTMBQ0FrL00dI3xxGW0JTjXAyoGqEUg222t7wA1WBhQLywjAHDYAcwzC5AT0JX6E/MC6wgsDwxoM0LA3DlZO7mWcyAnAGhvbJULAcH9uAcEQHsyCw3KN5dPLPohU6gPBAOgk/m351q7X/unyddAfHMRxfUcs0DIXM/O7SOuNnSJG7l12D38s7foN0AudQNkph644YJsoS4WYBNC54/VF4sGDLYIipRs0Xezgmm3GDGrFgOx2119WFtpkwHc7YC3nUvZ7TJvJzVSJgOyZF6/+J+nJgHkSL89TxnLBfNz/yl9hwgrC3A/Zg4QGWF9Z3ebJSpO7fYLno0uMwZIMyTdzLgHcLO4LOzWNzdMjOmnjS7gGuoDtz7S6OnKjRWLmSQKW+RD6LrVYWVZsDS0836ZCI2jkVwHNSr1Sbng2tOdyY3JbVAoF0OMP0gn+m7BGAcLSB9ZfkLZCIsP6DsdTh+caUKnLP2ovvxWWz+fadkX4vVG/KX91GoAzxzmbIg4xoGRd3xH9/mkj06nby9EGfk6L44ETNfQra8rv0r5lcr27sQ7E64ti7KyqPtYFosjdF+Kl4CXgJeAl4CXgJfA2ZGAJyzOjlx9qV4CXgJeAuelBNqICouhoDivSeqD/UyIixZQ/luytnila4wlbvd7+119ZJlb8rKay63sco1pAS9JxTXrS111T+Syy+QqSiBqfVCkxsAhF2WMFIBMsB2oLLoBWwnMC+CKhQNgPyAnbpv4TrZA3OZ6w6wrDGC1GBYWu4L2musoPslmDUG/te8ip/z2YMAQBEakYHVh7nQ4ZiRFJ1DVjtmOaHMfRTwOjgHKRq459V3FqniWO3JLzg1/ivsCIlIu/1NPCz4O8QK4yPHbJP9bqfhipJaOmFWIxQZBdmSTG8fND7a1ycgGADe+m1wB4+x9w/rEXGcZsWHWMvxv5fKfNpnPirMd8JttqrfQOKleR96QXFgFYaVjcRhwdYYOnVTA6JO60wInYYXQ5qbKzrJ4Fuzuh5xgbNvOX8Y4ukMaP9mg1mdSx6f62p965RXNj97xRNJoNkemSo1qtdbUnJd0xVFYlfstxTlIeqvV5rAsLoKuYrZaKGSPFPNZkRupWZK5q2I+OyUip7Xz/zNt7YUUvVoZV3lpWbiXOlUri7by2MFtrqGYBy7a1HINZTK1+S+Na6FMP/LJfMscafFQ7LxTJaIuWjn7hs+RADoFcchz+g3KzPtYq/J+xTsMGyCYe3nH8slLwEvAS8BLwEvAS8BL4LyUgCcszstu8ZXyEvAS8BJYXAm0gdAAIwD/ZBI7dFN3RTonBe3PkLi4VaQFLgeudgf+brvLrhh0hY2xK2w46oqbVrq42uPKO4ddblXoamO6X3bKRRW5KVhWdlHBQH+zdgC4BkxlcU0dscLgucWCGzAT6wx2ZuM2hnuy+KZdgJxGJJjFhQXspWzANFxLcR7l437G/jf/ROZLnDLN8sLK4j/u306IZIptswAAIABJREFU2HUG2rdbGCBn2sZuWnMNxXdcWWFRQXlHXOmRbnf0M9/ndrz7FrmAer6OQUgQ6wMXObTrO8r4oEYu1Aui5oHFIivadIT6cl8ShA1tJQN2GBmU7tJs1QE5GsFBOy2wJ1YoZiFjrqv4H6IHmaYBm1vl0B6LI8J3893eHrDcCKn5O/1PCaxtteti+kDn6BNALNyu0VdYMdA/jKUdT5UwFnCdRP+VRGbsbOkZ44E4LIxpC3p/RlZgT1X7Tuc+WFroOgJxT0+VqgcSF+SazXpGTN1EMZ/Ja1pWkPMo6unK4zuqLLKC841ArLcA8dO5NfMHMYOIaUJ6n/KLlJmXziRRvy8o/0SrEIiQ+2jjmRT6dLi25Y6LpqDzzH/trvOMqE2fIWfQr08HUfk2nLkEeLYSb4tnN1apn2t9Qk7yfhRqzq1oTuY8n7wEvAS8BLwEvAS8BLwEzjsJeMLivOsSXyEvAS8BL4GzJgEWrgbkAwSSAE0AjwGTUp/ZWFycCWmhMv5J+bXKV7rdf5Bxa95ytYv6sR447KoHK8LjelxuMOcaJd1P2EzUG7mwnLjs6rzLdAmvC9kNziIagBw3NjyrOAbAirUFJAtgPoAm4PclrbbQJtoDyE1bAGbbg5hSDu0HQIO0wJ0TIC7lWcBtwCLuxbVGgBjQxqe5f+I8c+MxHzA3SwvbBc1v7tEekJv63aVcckk87oY/sdLt/qPIjX+N83A5RT1xd2UWJMiDY9QJGQAys4MSl1GLmUzWyBVyh/tDmLBDc7Uy8TMgW2gL9eQYMT6oG5k+43/IB65D/rihQM6cb30LaAJA94Qy96IczjPLDPqR38gcUJ16mbsryuLaFOhtES1GFB1DXngLDEnpSf1GbmYZRF99qyXz9KRznNBxI/WMlGPs8P1pT0oRiPs9H/5mc8Pq/mo+l4nk/inI57OuvyefNGVuMT5VSVYv77WYPKk8zgTUbllZQPbeQ1HKVyn/ifJblM/E4oZ5EULM0mXnWK/Oi9tjsdJK7cSN6fX8z9TCpT2dgbXLedF+X4lzIgHeMyAkea/A/SXPXZ7LbHzg2VsRaXEUl4DVn07r124lOmfOzf/NOam/v6mXgJeAl4CXgJeAl8BFLAFPWFzEne+b7iXgJfD0ksC8WADWONuhDpjPrnjAX4BfQEADwDmXHdiAVGmshjMhLbTjP5aVBbv5KG+NO/C397mDf9/lNv3GUjf48i6XNI5ob98KV9vTcDm5hqofrLtmSQvqR47KGqPo8luyLsyPuSiLKxF2AZv1hNVvk46ZWyZri/nppy0s0rmO9prlA2QN5yIHFuWgQZSBn+dnt67hPsiL/wlayXcDyTkf0J6yLWYGZRlQzn1ttyyAHdcC2iNPyuA7ZXJPSIevuuq+e93kt1e5B3+CmB7mogdA3+qBP//trWs5DrHEMUBddk5+EVlz40VKtJt7oAvohrUTIBOLC/43AoVz+E1bqQ+B09nFCRnE8S8pA5BQDu8aXPdcZeJwIHNkRQBQCy7Ld7Ogsf6GMKF8iCXqQjBfI5Y4lzIom892Vyr6uahyobwLPZn+Ijd0lv6EtANYPp922Jo+t1s6Pe3JCpSrBVCnJJyy7bY3vTN58HtWHu2g9mkC2sxN/1n5q60b/bg+/1AZ92Gn6xaKeRpXd+2J+Ys57qJNHfrnotDri7bDT7Hhemdqt9K07/ZOga7w3TZBzCld7wFuAZd7nAfB/7gypCRzC0Q1BAbvIytfMHLX5Kd/etY9Ge9JFvzdyNFTbIk/3UvAS8BLwEvAS8BLwEtgcSTgCYvFkaMvxUvAS8BL4HyTgC1uAXiZ6wHMWYwCslsMB44DULOgBVjmf9yBABJjaVE5XUsLLaBLLdICcP56lzSLbud7lskdVN3133iFi8erLigErj66z1UPrUtdRJUfDURUTLq40i2ri6JIjbIrbsaSAqALdzHXtNpi7oMAyi2WhbkXMpdXtIsFOVYKLLxZqJvlBH11bUsOG/XJPXC3BMEBWA5YCJBOGexGByzgExdI7W48KIf/kDHl8537I2PAdXYuf68y9acu5urodnfvax6T+ydkTp2oH/7eaQ9l4aYKawTqTlkAy+a+ivuzY/KrkrH596ceZ5RaVgqQArQZvaAutMnIAwAPdmciBzJ12qRspAKEA9cChHMcPULncDlDNjdeyIdd/bgmov6QQNzvUmXuj3su5AGQzvVYWZBsx7f53kZnOR8gHvDF3mcM8G0Hdp5yYFC7Vrm/kV9WJ9rRTnC1mjbzsYC7pDnnnMEPC+LLzlrILupGXc5kJ/0ZVOfYS+e1/ynvs0VtzGkUdgLC4azIo+Wi6Juq7u8p/2ar2h/X5zOUU7LWYln86X0/NL9V7SRK+v32kZ9I63nj4N9jiWVpn77Yzu3TkMz5cYmeZwu1v92ibr4rQAOa7flAGR37EtDZp6evBNr0p33cMA/bswoLUp6f5oYSvTLykucpemOxo3inOJU5gTJ5x+E9am2YxGsySWPl0trRzCuHbg3HsgPjA/UxLDdNf+15ej6R2U9f5fAt8xLwEvAS8BLwEvAS6CgBT1h4xfAS8BLwEnj6SYBFp8UUsMDUZnVAawGZzb0R4DOLYRarAPYblAHrOYfFqgXAPWUptQD1L2uhDkD6K8pFd+gfDrlRbb5f/ZZB1/+8rS4sLnWZnryL8qHLr09cbXipm34s53qfmYi8OOQmvrXJ9WybcIUtl7owl5O7qI+qnDcrmwsiCAvAWIuvQD35j2OA7YBuEA0GHPF/u6smfgMCAJjvUsbVEi5M2NVvOw0BESiHe0EwALTz3UghykaeAOeA7IDtuEmiTGCuhoub0y4pF13p8TXu8IeuE1kBgYHFASQAoDwEB+A95UJe8InLp9TXtDJt4N5/KbnSV4uduAftANhAbtyL9kBMkKkHIObm1o3Zqc+5nAeRRFs4n3rSjm3KkBLoFru16Q92eBopRB8C0JhVB+2n7JcoI2t2aGOtgRyQJ8QEx6kbRA79BBCKbm1qlY/eUh5kC32UBra12Cz67kTAnQrIwyUnndpICogU2oYOUW8LJI2+ILOOYFPLJUen+6UAl1xypHVnJ25NTteiq12gnDaLw+R4rwvD9TPfmw8MpNZVr1/z0dyXw5v6qmEeXbtBGVkDKKPX6P55Q1qctLDPwoktQN5k2b7bOb3bL1978xndtQPg3d53VvZ8wHv2nmcL0BZp0RAp8Y+6kREWzFuvV/4H5XYLLpMJY8zGLUQkiXHPuEvdtU039w53R3Cu+GyrXVJqHuiTfE3vO47BM5Wvxo+RhGZVyFxMYi6wudossjhuVlnov11rc7mVYWR0sy6bwaBfRJ+iLQXLlQdcGCxzuSArd3aKyKQysH6z5y33ZG4kmzUac+HIUGYg/siSF6dAsNp81uajVtv9x/kjARs36JrF4OITXeAZwTOUDQ68D9j7BnM1Y4uA2Xzn2cJzlufpMWTCcUjvRM+naREU3XoO5OIgLG6ZfmLry498oZSPq2v1m2c8ZfOsZcwbWXL+SM/XxEvAS8BLwEvAS8BL4KKTQPsuj4uu8b7BXgJeAl4CTycJtLmEMtc9gCeAkixEOcYn4AkgCgtUiwMB2A/AgrUBLnsAiwHUU3c/p2tl0S5bgXX4TQYsZbc9QG7ierdtdstfX3C5NUuFJNdcZmC5LC4Ou66tebmIkoVFV0YwUuLG7yi5vudVXeESBeguTLv8GhbskAo8w8wCgIW/AWJ8Z9ENOM65gO22s92AKxb8FpwbcgYgGcAJOVEOQC4ujQC4kCHX8Z3zKM/iV1AO1wBYcc//rYz8CJr9LOX7XfXARld6dMiNfFHkUG2DO/D3u11tiOvoHwACSCPAZHxKcy/rFwAK7ku9sKq4Q6AlRMGiJ+kObUM/aBuECYn7IjfkCDQOmWVxQD6t77T5JmXk9QJlrDDQLdoACAixQF9A3vDfplZ5HIfQ4F6QDoCeBB/nflhq0GfEJYGAgPzAIgMdRS52HfJAXhAXyHnGzdYMUUDfAPpQDn1C/xooT1D5MwIJBfyouCctIlpEBeAo7YF0eaGykVv0IcQT/YauchyyAPByDlEwH2wSAItezVhG5V0crnZxoFGh7ymYlIy6/nCL5NOQZUtD5YWumFRcdyCtSqoCtOrqh9hVvrPuWdXfdO9efTBZld2d3XiTgslEPY2pu2ph7nBPY/rh99/31qEXHr2z3fKjo5uxp5MPc4HnRurSlWYZhazRX36j5wCCAIftrlEW1J2FAPeWqxebk83Ky4BxyjaXaUYamrVY+658d7YICwQgwoK2/y/ln0mVe2asbRGZwXPAteRlOs4Yo27EncFSjTEMmckYZ14rLM9d//Ure37uU4GLrmwmlUf2Vz7/IzvL/8KYhNQw663WrWY+TkRYdCD02vuQIgB2mauYx5iTmFeQKbvKmc+RPfXbpMyz7tvKzBucx7XMS8xpzBc9mnlpYzbodtMiJo5IC2KVtizocoVwrcjXGVuvQxqTG/XPdmnNdzRab9QnerNC1+Mir1tBmb6pzk4tmsaj7rumomJjOOrf/0Bx01gurkfjUU9UDnPUt90Sa0YobelE8jnmAn/gnEugNfaNoEAH7fm5Vd8ZP2Y1gS7eqIwZE886SP5NyjwrGIPoJIHreeYZWcFzLp2PmBuOQ3inp3DvB3u39Xxy1fcXD+VXblhZHdpy5eTD9cumt4+uqh56eLA2QlkWOIV5aQ6x/nSa/8+5YvgKeAl4CXgJeAl4CXgJnJQEvIXFSYnJn+Ql4CXgJXBBSYC53cAvgBJAUsAmFqF8AgoD0rBTn/8s+PTsblIdA3Qxv+NnHCcBoL3lIgrw9g3KG9zkg+OuNvYV133Nq0RCBK7rklEXZBSMe2SpAH0tnptlxbPI6f+C3ENlXCwSo7Kz6RoT/S63NqdjieJcEDsBgIpFPYty2mh+mFnQA0S1JxblnENbjXgASKCN7CymDGQECMe5nAdYwDEW8BA+fHIeMrJ7AiJ8ShkAb6lr1q928Zh24+7cpNN6RVpErj7ScIc+st81x6gvfQRRATkAmE39qQ/3IRAuxA73h/zAqmSvZDg3CqsOLmKi/bSVupnrKo5RP8gU2kcdAVqQL7KCSAB8tODYxALhO5ndougPssUCAyIMIoMEqI/OAeZzfFOrXHOFgTwguEicwz3pR0AdgFHIDGTPdT+ojBw/2zqfcwEdIUm4P7oOKUTZAMFhi9g7Y+KidT8+uA9A6eWtuqADyO2Vbecw1pAhBMu/KctGwh0RSZGSFunu8J9Oz07dSGknNy3sSupufRIG68Ji0qV/epIkcEEj6Y+bQSYoJs8XJbNGd+9r7g9uEbA6FeSSZ0pDI0lghzT6srgelK+MHz76i+FfNidGepKvhc/b/GBxW/elpe259eV9d68oHR66ZuJ+C5KOHJEdYDWyMlDdQPozInraZHFOvraRFLQDHaa96BnjChaKvgBEhKhkjCMXiF2OG4BHHxqRsKA82oBK5mHuZTuqIeBsPsEEgd+pL3ll9J7xj0s42+lsAcfNrd1ZkZ2IibpIi99V4a9ShpikXq/SsX9uBfamHQD6jC8+IdwYu4xvxvVPKaO7kIRjY41HRmvx2N58uFQu3pI1U83dU5mgq7uRlGgzYGx1vnXBAoCrbazis/05xPzJvamLudtjzFE+4w/XctznVmXIYyNbmD+YzwCFmaNmzEBm3OXwPa+R+A3lq9WaS4PQjQRL3WPKe4Oc+igSIQhREbnXybJiZVIW0VpQHUKVH7Q2A8zbCtYMwjdXdXJdTKJ2sh8QgfG11Y2RL3ZNV75xf3HzutDFvbmkLjA62F8LMuOSi7d4anVK+0cHl2T2N7ppz2GO2bsP32fH6FNJ+LTGvz3jea4zpmzjxIv0nbmHfobcRieZcxnz17Ua9Vp9QuKT0GOeX1zD3MQ8wdx0sslIklXbJh8MV1YPN+QSKr5z6QuHHum5ovzssW9tKDTLjAee/bxvMIYtdtfJ3sOf5yXgJeAl4CXgJeAl4CWw6BLwFhaLLlJfoJeAl4CXwFMrgRYAa7tNDSBj8Qn4uEnZ3AoByrE71uI+mPWBLfBZFLNwZbHKJ4lzaothZWFS0WKeOgDmfn96r6ywsajnErmHOuJiWSDk1wy6lW/odo2xxBXWR7K8yLhMb9ON3jnl+p4pfKcswC/OucyqIdd3tYCpgsCiwm4XZQyUYjFvJAQApMUSaCfp0+Diyraz3AJlm29/IyqQHd8B6JAfwCLAmYHrLPApZ1j8yuOuvONZLuoacPUjQy6O17nqniMuqRfk2ip0Rz97UJYW5qbEYokAxAOYAmQD4rMbmHM4/knlW0VUzGzpP8tJegQUh96QASyNpABQAUIHMCEAN4ArQCD1/gFlZIT1AEAg7TJwhXqjl+gS10DCID/Knp8giACJIUJOJpmFC7pLwuID0sJIkk/oO/0EcEk7dikTwJzvBn4mp2Nt0W5hoe/m8oW2AZgCOEE9cLxTAqTCCuczyg+uL+8d+qvv/nxDFg6puxDt1u4R3HZ50hNkw66kmFSDVaVcvjteHS3LDjaf0aiE12Xi5kCYTZaEtVgqL+RpMAzrw1HTTSZ78836yuzGeIaYzKovmq4+FfRUD06tfPyRytbVXwpfkn+8vmVo3dS+6ReXbju4LXjo/RsP7qrm69VlSU2WKbF28MazAL65QjMrA7NKarfGmG3jud6Bu0CMBfraQEt0E5AdcgldxioI/UAv0FVAw+cps/ue/7HYwa0Z+g14iPsxdB49TefFVuPT8gFE26wpkB3zAucwNrAI477mao15yUB+9JZzISr5H0sFAHR26FMOgDzELGPErD2OIZHP1AJD5AR1wFXb37XaNVWNj66/e+xXaS8yYH76SWXGMHMEdUHnkeOcFAX5b28ofP/WDcXX9mJwcM/Ee35zsrETn1qAtZDWyJV21SS3tC3zCAsjjm3ONhCfuRgZIVPmCuoBkckzjXmKZwp1Yp7imltax7HuY3c696I96PRz5te75Thqj8bhBnpEFksu5E7q4UDUSKgejGUHJmsnJ6uL4ybMMWphxk2GXe5QZkn6XWSFg7woaLDJNdSe0ah3Sr8n8kn9b5Y3xj53OLNk6mimj/pB6JzxRoHj1/DC+nfe+Lb3HT7RTTYSQG7znKL/eQaZNSLkdkr8nU0XXBr7zOHoK89u5hojz7AKZI7g2Q5Zz7MCfTxR4hn3Z8o8O3cpM/dgcQGJio7MElsdLCyQi2VkwnOJOYhx0t8Mor5S1FWRe6hDvY3JLXILhbwoF8tF5kOb82freK7n9xMJy//vJeAl4CXgJeAl4CXw9JOAt7B4+vWpb5GXgJfAxScBW5gCdJtbE2AWFtAGnLGAZmEPgAb4DmjMgphdfQD85q7GXGKwSOb6xmKSFXQNALwW9wR2pfylsjwgUxcAuW5ZUYy78bsAGNhNWBeBoeX/qjUus2xKvm4qchfV73qva7jqvctcPLlDFhhXKLbFCtfMd7uw/4jLKFj3jBwAs1iEIx/bBW/WJ0ZMACSw+AdkMHDT5GmuWsxqAwCC8wFA+ERGA6568A5X2fV8WX50uXha5SR7XW61AotPTbnmlOpYHnHDn6m78mPssjQ/57QdSwTqSXkAeICgHKN/yB9fzMDayP4Eib5HX8joByAtQClyeKkyQBCyMvdXHAdEQQ7mAol+4xp8bgMIonMEH+d6dAxSpFNCBkZWABxTjllZdDoffW5PuKxCXygHggRdogxza4H1A1YXgKTIHH1riqSBtDgpYNCICrupflMHwG3aiCsP2gggdbyE3r1d+W0KevrOd+36nX99Rnx/t6wjYu3WXiutGoyXRi+rrMj15PIN8XBu63StuHHn8tXZ5kBU7EtKQTZpiEFL3JLGpCs3cmE2K1ZiXSbSTu5NuemaW5EZl4P9eAatCpPseNyXPdK7/LptfY+4Dcl+99naKwaW1w+LMfz893R3lV4ThGp+4nYkY+7b8YisruqST+JuV6Yf6S/GkBFtEGvIjmSyNUuMEzT9Kf07JYCUzQ2LkW3oCMQaljdY5zDurW3zKwh50Z5wyfIPyhALAHyMV8YzwGijBVjaLmjK5Dj3wWXZm5QZDwCr8xOA5vwEWcK8g2UOMmeMfUQZ2dMmdJw6WByGM7Z+acWyYF5+tzJzVU8Y5H4wdJm7Y9fAeoox9uttFWXcGGE4p/5x0rh8qrk3qsRH5D9pOfn3ptyun0tcglyY44jtg+XYgwKiSy2rAnObxbzCfA2xnbqYUqbPGFsQToxhrKywBuEY/y+U/nPbH5Rhifl1buLuqp0sKTZATqQzvO4k64r0e4RtiUZvRA1OkOIkdOOZLifywU2HRbcvu8yNRj3p77aEjNMUuuSZyxrj76qEud1REmcyrvllyWVIcjntGFInquMF+r8RWegHcxOkHs8JnhlkYkD8hDIbCf6Psm1MYPyUJFM+z5i4mBePhjoZkQaNBXHG3Mj8Ye8iP6nv1NksV09G/Dw3aQcWVyQID4tvcaJnFtrMXMQYgrBAi5n7IC2Go6T5DLkFzHcFpbEgSXhWQoRQPnN+R5dtJ1Nhf46XgJeAl4CXgJeAl4CXwGJKwBMWiylNX5aXgJeAl8C5kUA7YcHiFJDDXCSY/2NqZjuLWTSziw6glWSAvAVbBgjj+XBcn9pn0tQWEA8Ax65kdv8B/ALo7VJmwW8g+BG5U6qnmQX1yOeoF+Azuyn5PgNU9F3f7Va9aZ0rXlJy+Y0lV9y0z4XdK10olGgGqAbks12ZAPIADEZQAKIhM+QAyUG7zQULO6/5n3txjGtqrtnQol7gW2W7rEKqN7rmtKIMlARI5COXG+iVdYg22HbJSc8DNTdy6y6RFQD7gGtWHuQHoAL3A9ynToB4uyWbe/V5LhJ6AViBziBv+oB2Uzf0hU9ANoAQs7igr2iDBQU30gNghPZyHJAV3TNQp71tWEbwf/tuZ4BeZN2JsAAkBjAGiDF9pjzqRaaeQIrsXgf0hQRBn0noO7vX+Q3ww+fUDGdxynEtaAs6y05ZPiEsGD/HJIVhoV+3aHd1O2AaFePyW3d3bbyi2cwM1OrZcj0MG41CJldeX/yeobVLtjRyUdQfTbv+eNpVCnk3oZ3aVRkWCWxyIwI+tSPbjUS9brA56dbWh9Od2zv6FP+3vNv1haX0t1x/SMmartrUdfpcGhx1azIHXGatxJuJRGyoVtLEeEgAcNNdEkq7E0k4KSmWgdFyMy1iF/tXlO9WBsoF/EKW7FoH5JrWDvnU8kI7cU8EpnUS02Ids13OZh2CngJiAm5z7C5ldBIC4VTfgXE1RLaEq5bbBTD/3431wztLYb67K64+U8derAzYiMu0n1P+UeVOVkXHazN1np/Qs88rf48yhAX9wVhgzNWlZWZ90bHck7TAYJ76VeV/oZDI5d+cCbv7avH4b+gnViHtqSNZwQmJi3vkEsplUv9JErQCP0g5zP0SlhqQH0OhaLru6fKhPe8cnHCHRugrxjV0gZFiEOo/poxlBlYTyGAxEvd6MjGrSxuobqAnRaiZJzAbM430hKcMI/4kUlMjTrrgJqMutze73O3OrXSKXXHcK0Uv5h4ubPgfqayS5uHBxsQvjEU9D7z/nlfvmQ4L5bNpGXASTXpKT1nA9VOrh9LnOHrIWEYfsNTkOcHc86/KWEz9SKvCkFrvVzYXkRB/kK88Q0y/Trpt80gKrrM6URfqBPHIu4y9z1C/+Yn6o9OzZFXbCTxvzW0izyYIBJ7HkBbU295RFiInqQ+Je6C9PJt5FlIuhOM7Wv+nLhz1XLpNzxKetbxvMK8w40PkHTN/e+uKDj3pD3kJeAl4CXgJeAl4CZx1CZzqYu2sV8jfwEvAS8BLwEugswTagmq3n2CLVHbvARwDxLCrb2b3/8wOX+AWc7djC37byU9ZoCkAQezm5TzKApSmnFj3XXQrizkNmAHo7xUgYLE2AAVvV7adttSLranspqRd7AY0CxEW11k38Q3cMRXd4Msrrv/6PlfZmHGFjVWX3zDpMoOjIi5YuBtZgDz4jey4J/eBlLBd++aj3lxlAVUhizG5eeoTMTHsyk+MuOyAAJFGn2JS1FzSyLrcioqrT0Ru+uFhd/TWSaedsu7IzQJ1EwA6AN6ZMmYsFdjVSBtxqfR15boARdwYnbOEpYH6GjDHrFsgHADhkRP6AkALqMFxZAYgA/gLyMIn13E98oI4oN8AJmm3WWCwIx15kJDF/a1y0FO+08+ATpbQx/Yd1GYBhK6jo/OT7ZgH4KQ/Aa2oP/VibHxRGXc7HEPvAYQ6ujjqULYd4lruDXAM8MTnQmTFgb6GgkSEXSvr4dyN/JNR75bf3fjOLRsO7Gk+J/x6dbIrt6+/MjVQ35Rdvqt3ZVAT4bC8Me6+mrtKu7QLacTf9rQ/O3PLPcJ37y3SzJm0vWut21AbcnIzk/5eWpt2O2rrXSauu23BI67QrLCjOyUyiGlPkn1SChMngqtjaWYMPCZID5c4aY/PWAmQLaELZAgAiCH0A7C7KeICWTcFcp3xrv+2+81+PQ6gid6hK6Dk9BHjGOAfP/GQRRAJgN+LlQAo10mG2YHm1GfVB9PXlx7dJ8CZ+etGZSyUXq2MNBcjQcKRSRBHjK3/2/oN0AjAyZg6bbnLyiK+Y+d3bylGq98ut05/KguLl3ZFa1aLsJhPVpywPbVkXEQFw5Fkj6k5l/2+qMI3Kb87DoN79HmVdnujtIxb+vEaZZT85094s5kT0METOGqaLWlm/WPV0tAKNIuFmoWwqAg0CwW4hNLMpWa4NKZMe5KEY1HmnJcSHaot7p6SeuDq+Yw7WpFlRSJPgDL6OxFZMb9tjSBaeTC79GOFuHaL4l58MJc0bpfOj15MpEWH/qa/mPPRCyzZsF5gjudZZOkV+sIcxIzF+VhQkS39ub5AIj4keUL0VU5TprZBBD3lWUZdGB9oCQQ2883xEs/ogbveAAAgAElEQVRFzp9v2fVXOgYBzPxF2RDBPEd5RjEumnpH6Di20xhIM21GI3k3oi5cx/PpF5WZ4S0xRnjWYk2FZae9ZzGHzMz2PnkJeAl4CXgJeAl4CXgJnAcS8ITFedAJvgpeAl4CXgKnKQEWqYB0LHwBjdlhCzhm7lDYpcc5LKoB6Vmks6BnB6D5WeZczgNINndJAD+QFrYIfkoWsVqMf1SkBXXAIgIwDp/xtjuSurAzEYDCrEhsJyBAxnWufvRhd/if+pTHXc81sVv3i8tdclfB9Vzb5zLLQxcV9yiHLrcKoJodyizikQOLfAACwD4jfgyUqLvayGOy1tgq5CrjKoeGheoWXWbpJjd5z5SLCkXF3gDaGnVTDyn+QCF2zcmGG7trzNUOIjfqSnsgJQAPuK/5wae/3qP8JbX9KZGx7nWihEzNzQx9AfiBfgByAJbQHyYbdI/dn+zkxCrDLDOwGAHQx+qANgLCIF98dwPi4lqHnbEQaq9rlU29ACjnJ/QTUAWrGhLlAva0kxrt10B8QJAYSAz4Q525Dh0HxOHTCAvGBURNeLKuoXQ+cmG3OPUAVAIoI1lMmPTHiurQ7ylGxdEbj37lwL6utWNfXPayZUezg6uvqj5Ufih/lSG57h2r/iB6V/dvFwu9w1vymelMOSdrCu3OJsnPfXvbTuq7AE/3RP5JfDmQj5uHG9e44XhZ2oFVbSHvCmS1ESqevYJ4Q15YAoCNRENJm10gWg2wFp/9KVw2d98tYD0ZAoB55beUAcEAmJHDkEA0xlPtbBEXbcKweYp7o2f0OZY1jO/vU24HLU9KhvNOgrZBb7Eamp/6Je+3Dkf91y1pKjBIWBjqiSsvxLJF8DVzGAmCcrETICn5zcp/oYweMj8SWwadJp0WcfHtiXfFV/W8/YHluWenNgXben7xqrvHfln+0xbclM49mR94rkCg1AIX/SyaZWkge7k7VP2KKjTrdn+mgoG7plLIve7eZ152+Pl3PvD4wNgUczEWHm84DYGdLFkxUzQkRespFyxx2xWXYrU+c3qa5pgBFWZCMZRcABkBmZEmjQN5ZGvZtOg7Gi6xNNXi2lJ5UqsGIgblok2Pmfs3bnaHC504VY0xWUkpjsBxm6jx+VqRX1eHSfI3Wdf4G4HsPJcX7NOnMqj0afTNmVyCIjERMmfynWcGz49OqZPLNTuPuYDnBhsePqickhanWDHub+8IPAN4FmDhQd+gJSciK7gd8yMWa4xfLEV3KbOBgZhVEPJoGPVKXc21zm8YWdEhOH3LmVn6nsccyHMYxcNqkfeLTok6UH/mDM7nHeWYQNvesmIB6fnDXgJeAl4CXgJeAl4CT4kEPGHxlIjZ38RLwEvAS2DRJdDu7xsAnsU8C08WukCLAHeAGyxE2d3Pd3ZE255Sg10A0wDVWRyzyKUcPikDYH1RA26fSAot4P5zIi7YCblJmbZRH4AIdlbarkSeXwDh7G5noc1ORKwvWLQnbur+yD3yVsGumaVu8CWPu6WvWK94Emtcfl3kCutqrvT4Y27FD9Vd2LtSMSgOK0bGVsWcqImYwEu5wAP59Kgd0Fb0/IBrjF6i+BQKSFwr6XfGlR7Ju8KlobbgAowqCHgzkOVF2dWOHnETd2Xd8CdB9qgbu7qRO3WmDwD2kCmkBYDBLrXXwMUTieYp+b9lZYFuAICCqKFn1NVioxAwl2MAKxAJm5SBtAFs6CcAE4BLwFrIA85DTpAUmAFwDJLDEsRCJ3c57CAH0AEcMrLCrkFfv6mMxY1BiW1FpjqMXrcDxVgB3KEM8MXud8YJ9aCd1PGE4G7lhwec4laYVQ7kCkAVPvJ7BU4/qB3Ws7EItkw/8YF3PP5H2bWVfVdsKe3cdrR/8BlLs0cPf7X3e3vvy1874yenlUbDJYrC/TPBC6LPZdbnd7iuEHEvTmLX91Sm4Gq5xG2P1rpS8nyXi0N3dfSAG87063vV9Uh15dZozg0zQF2SPPY28uaTkhaJRUw4VlJY2uCOBXAMAAyyALlCOB4UwAYYZ37RF7RmOU1wzMgKdOImZXSFvsWagj5i3J1sQkfRCQg3CAr0hF3c0DWdyIrZcvfkVjxHli7Pwaplc+2gLGMmUlD6BIl5C10F9mZcwVJJZxcK57ygihITBbdjlIUcCOjOHEOPnbAS7XUUKI48s0dr3y6KsEj/kjunoDfa7MYa4LyzCXCVMc+4+pQyRPJLlFHeQ2GQOaC4FczNgMsuJyYgCESNdZBJIxO9eeWh0TWFSo3xfDL9Nd/qqr1etN2s5ZiDeS7wbGMue4aGQ0Z6fbsMP7pUpS65frpBRw7pe0MGTT+qmW2prIpGdCwjC4txnT+z210chP4ryuJiQjNFWQTGGsWdSTgviYOkORQFR9f1u9KUHrvDifvsNrjZhdP6UXk67MlpbBYVlHuWuzzmApFhW1SH388362EmbH5Av4+04n0ct/wL8c8FLKd41vDsf64yQsU6od3S61SayoYBnkEvV+aZ82Hd82v6nDhJSwvqgj6go5QDIco71WuVmW9OlHgvQDf/RpnnG9aVvLMR6Jr3HNs4YhYVZumZzpkdiArbOMAzkucg9aJ8yvwDZcZfp8TcfJsy1/HsgzQpPQXE8onk4//3EvAS8BLwEvAS8BLwEpgjAU9YeIXwEvAS8BK48CTAQtV21bGotcCkLIgtWCnAlbkHYQELkA8YxyIbYAhQmmCOPAfYmcp1LHZZLEN2QHQY+fGUS6gF5M+C+a2AtriOAsSm/gAGgM/UF5CctuISBfSHYyQt9BtDintxqfKIC6JVsq4ouDAz6qKBa93+D0y6qEtQbLxERMVOt/Slg27q0SMuv6Tklr9xq6vu65OVRM1NauN4blnOFdbnXX0064rrym76AUU+7iq6/IqMG/tSyR3420+42jD1gqTg/tSNfsFvNkgfAMVDate59O9/Uv3YIi0AMgCHAPrQA8B5PtmVip7xn8WCMBcu6BR6ZIG2AaoBmyAy2M0JwLlJuX13LP/jnmt+op8XSgAzZOvnk2kXsQU4n3HzJWViDJAsLgnfT0hatK7v0w76zXEQvka/U8Kknay4avLhT3/v6F3uuul7n7elubMv31crrcoevvRnK3+d3VJ8ol5UTPi7k7nNe6y8zWXDisspbxBpEaZBs1vumuRbTL/m+oM6Tou1I7scB7O+eFxeZW4sbHf7q5vELA26fEbIcNysjgddvdXMKrdFAHu33ERF7apJLyoJlHWhYL5YzkICaTQWF6lWd5YU/Uo9DVD8mL4DxAOIAahzNUD6aVkTdQA0zZKM8c98gPsljkGg0N8nkwDcaQ36AKGIblMeVkPo9Rc12Up/kxH18SWC3EvqiwVB9W90XS4pir8E+RZpIXc+s/3Yqsw/65Oxc6cy48fi42ASM5gEkeaJ4FmCwCFnNydB6kesHCSxSCDjmjsK/2Wt8l+gT4gWCJZdyszjELnHnXdaRAVF8DzoP1L7xrZ8edBtLhJ+Q6ZEhZvc+NR2LCQgdehP5jRkxrxGOyCnIB+jMMg25E7q8yIsLm8k02Em6H5tb2bjUE+j/+bJ4MirZct0jP/+3ZtWvWTF4VG3bHjM5St1J9dQreZ0/MBiCmKCZxqgLGP4w8of5P7KgNHMN3LHlz7zIBYOylLi05qdBuT2qar4FM8UIXEFxIP+2ybRVpUj5aziWBiBesxufVkgPWnFIU2DEKxFmeDo+j73UH6D29+zzE2unbGOWigtGxt3l+zb77K5ppta0uWGB/pT0mK/AnMvlDTX/GquWj+sun6yZWnRPEmQ/bh1Oc//ROF5dkBUQBxisQcZSkLn5hC/reP090Zl9BI9ax+r7S6Y/mNLTywmEu6QZqINdU7oFXXhGc8YoaxfUYYUtRhJna6E+EQX/0SZMc/cxKYFnoUQ6DxnIdZQeL63kxQLVkZ/pMRiK9NOZMMmAbNAbI+1M78cSBrGKq4RuTfz8nn/XnI8Yfj/vAS8BLwEvAS8BLwEnp4S8ITF07Nffau8BLwELg4JAM4B/rFTFxCMBSyoB2AVC2KAF74DMbLzmfMBh1nEs1BnkczueK7nP8A6rqNMFuEnDZKebXG3gP4HBCgAQgFIkNnRDgAAMM6CG/CYNgA0Aqqxwx70iPZtcElT0Yf3A95JTrs5xwB2ALAjbvQLLNwhdDJu4t5hBfDuc93XZF3P5Ymr7G0oNkVBTsqnZJGhLeuHym70Sw+4+jDyphzK43oAPeoCsM/uSwAUAmmfquuJsy3S45bfFs/C/FsbKWZEDAArOsLOaogAdjGzm5nzcA2E/NlxzY53QBSA6s8pAwICsCA3wKeZbdwzACSA86mk4yODMyUBZgI2cS73+4ryLmX0Hv2gHtS/JLdQqZ/w+RWQLGYPycVTdji3bEBmNePTUTeg9py0ubTzA687fPO+jcGeQxv79zyn0FO7RA6nhif6uvviNXG0LbxvfLoYuYcntrrxxlzDkgenn+WKCpZdGCi7pZkhkRcKwdKs76yFmRXdceVIMwh760GmW0TGsGJlH20GQY8AU0C7UcBWfU+tAERW0AbIvsE4UQDgZo/Iio1uutmbkhcl1517MLd5eDzKPerC5gq5MRq4qrKnry8udbQK0O5zl1VPEtciFsWZaASlsS2OhbjQBcaipRm0e2ZcYImCfjD/MMcY9XG6QJkBdpBj5gZsl77/9/l90uE34Drk5m3KuGYBULQ5lNOZS7fLHU9TQbSrGdcsSu436felS5qTBQVDvlrBzrFBOSZ1xRX3ra6tbmdulXvh9INujYKhZ5Pmr6rPNulkxgFjAHIVKw6zgGD+KMRBsVjLbSYM+v4wLn8mE4/Jx1DzeeKqloXx9Hf1HVDyTTNE1oKGKtTp9lbZ79QnJC/zEIBsRxZAALi5uWFs04dXx67xjsPVr84SFityz3d7ok9Jh/ayc/vHlZlnKZf5lPrzm+9S93qi+BXB5szLH1UgoZRUjILiiit2TOzd1T+2faqnWCx1F+aQlIdWD7p/f90L3Cs+8w23fs9hl6styGkhN+QHEcyzgOca4/ujypAoEKvoGRZ6oyImpkW6Qd8F0TbNPVk9N6AvwjR4+gaNGwDnTlZaVPuESWPSSR/cE7nVKeFAoO2F0uqDR+uDRyfKcRT0du2tBBrTbkUwqkloyAVbRXyszLqb+1+QkiDzUz2MBuuF6P2yQnnr8qGxj8sqxcbPCet4gZ5glmy8qzBRQoK2xwlqJyssdgkEwIeUoVt5DkMM/JLyWxaQAc8bCNWMxgBWDqXg2puPGSN657ANIugJ+kInE1cFkpTUiTjh+C3KkAKQamwgYV7GMolnoZH/PHPSYEMLxaewurcsLKiLuQFl3tukjEUjbu+OZ9bD+PxrZcY3Y4d5Dxnhsu+0CGSrl//0EvAS8BLwEvAS8BLwEjhbEvCExdmSrC/XS8BLwEtg8SVgLgAoGXICAMwCGgP8sthmkQ4Az6IdUBkAB2CMzDEAdIApFtCcx29AJX4DOFFeumgXUDsTtfc8Si3gH1dEZFxHASKwu/hVygDIuDtANha3gN8s0mkbbTQ3Rym4pgSIwPlYZiBfnotNN/rlaWW1P1T52uA+cx4gEffj3gAplAUwj5y4N+DZp5W/oHpa+a3bXHgf9L9AfNoOoMFOUfQHYoaEjpgvb8gvQF6AJQtsTvBR5AM4ArCCNQ9AKuDOTcoWEwNw8eaWDNHVk90Zf7ICbXcUb5YhANQQJ5Be9LdZAdDHtsP1mPK//mvXZf9i9OvLH+25/PLxbP/66SJY+dy0pfTElS+Z+PLgNYMP9OaW1ZdM5ouZaiVb37V5dYK1wnQzLJYU5mRj7XH33alj8aV91c2uFosXE6LaX5++fUVt7OP7csvWi4R4QgDnzpyrl6I4OXgk19/VdAokHzgRGG6vdvWjb8gWkoi+4fNlzSSTrSV5N9kccN3RpBsUETLWWOpGkqUTPZnxSzNBbUDBonfWXOab11R3XrOkOb1iIVdGIfRO1e2PR0R2HnGTchH1rHn0Dn3aaZs44852wENsMSY/r2zu0U7Hkot+26QMeAjJyA7s/+8ESgF4yDUQauwsBuhkvsOygjqgH9GKxljQ15xOrqns6lLQ8yVyl9VTDnPdE2HXoADq54wqWPrh7ABEhHugQHFPpqrigpCOZvrcV7uv+vgzyk9UVzdGpgcbk18X0cA9mSO4J5lxZcxD6btbD8s24UC+u/zN0Sgei4qVe7O5+t7RMKlsippj1UZm+e9EzaPvz9eeeG+YlL9HVhhqT4LdC1Zd8xO6AFDKPMX892XNlfs0L3VyEYUs6V3KAcRl57j0cNwdqH7Rrclj7KGJL7OxVmoeFHvboA+Z52gPu8Lr2u0/h3giCPDB77+pMXbtm44mmYj/wtWHJ3qCowc2792wcnkchq5SbJnxtNV89+ZVsrJQsO5GSVYW8T1ib6gTJA9EGEDvZ5UBipmvAajpN+oOecHcQ5+mVlOR9psr0zbmbOYBnhPsrEcfmWt4fh5bibb6HO8rxALWNFNRQbFm+ksiKzqyFYV67bEVB0e3D4xMua5S5f5aLrMzP1Xb3TcydUMUx28t5sIVcRgpNFLgXnfZV923i5e5I4pdI5075vaK9/HXl+zdv2ekt3fPFz907c77n7Gl9jSztLB3HHu/MX9ZzGcLJd5hGFfoA9Zz6BvzO3oAqYbu8AzqlIiX8sPKv66Mbs3642sRFbxHzLgFm3m+/bYy883xEvPLB5SZC9HHv1KmjruU0VcIwgWfMxR8HPdP6BhkH+UQ54UxzoPoeGQFJN//VEam/6aMdQUEJvPd6RLGJxCB/9tLwEvAS8BLwEvAS8BL4Mwl4AmLM5ehL8FLwEvAS+CsSkCgMeXbzjoWzubGCeIBEJ3/WMSyq5+FKCAPvzmP/9l5yiIZkIb/WcQDDLP7nTIAzgB7bKcdAPwFsZBtEQM3C1wAdGT349ta7aD+AJQADgCkFrybhT5goREVCHeXMgAH3wEWALT4LpJHDv5nwDEW+8iFspAVO/QBMkxmv63v96s+p+KmSJec30mkRbNFWtAus+YB4AdNM9AVEAUdw4IBXUQ25rIDQoedsegiYBDgIjoH+AjYCRECoMjxXcqblM30gPvRj6cNKupa9N92twJq4saJPkQ36D++245X7qUmCyZtJQFHIVk/C/e4oHD15IPrRrNLXvRQ71VvtXP47G5OT98wdufOtx19X3Jt5ruXyb3SiuGu/u69m1bkonq8afeSlZnDGfBRl+tXROtn996hneihe6JyRWoBYWm4viq+8+irvrKt6579Swp3fCETjtwXZ8KuunzXN5NoOJs0KtPZgkU/TskYVRZdps7UE3kDlEEUfURkxRtlDRIKLJf1RXJJJe5ypbjbDWSOrgpdM3WRIr/4mw/nlvy1QORvbKke3LehPvQugfQdQblwi1sVrne3Cqv/RPNrrhgPyzqhmQLIaayCE6SfbP3PWGV+AvCmTyCzhiXn44J475u5GP1iDkTXsDhAl7j+vxzn3rhFercyVifMeQB4zJUcR5YpcPdLR+DNZuVIuc9vlT+Za9bf0NcsUecV64MjrlzNK2B04ERuOBE+ThYX6e2bbUZpRzL9rxNp8bhIj5tfNH3/p+QiirmnOX8n9T17hVS32lbPrCmM9f5goVZXXJzif5Q8gkYmKO/Jx4fDmuvK5pOJIytH/+d7e0p3XZJtDj0oyLwvSOrvULXlquaYzeFvVrHoCO1lfvsHzZPMXbHVoWVdQeUh8SA3UrJiRhBNBcq+c5awGMhcVRup3x+IyCBmBSAwcoOsmHNj9SNjvW/Fl35nS3ntsy+vrLomtdQruoH/evmj+13XdMWJtHCPbz0WQz68atDVs5ETMP/JfLX2SNSMcaHF3EK96T/0G8KY+Zz5hDkEAiUdA+aHv+XaB7ky6NAVnomQyujq8eJk2LPPiFkTx5xPs4IgwL0Crrt9uRUdA1GoAqO1TObb+9Ytf0hWVl9bt2fo0Po9Q4dlQTIZNbBXcqNhNX53eDDppjUrukfc9asfcQezS91d3bMhcdrvHQ6tX/Jfe4ZLX62F2Y89+xuPPCp5s0v+gnhedxTm3IPoCvqIcuDiiPgQbzrOdX+m/3if4VmBizL0IyUelQHy0VWeXbhJe7Ey70Dz0yYd+EPlKY0HYiONai6weQYLToguXEHxHDseWUEZ6CO6iiUFcwhEPvpZaxv3HePKdCAprJ7IxN5B0F8ISMbcTyqblUeHZqWHeL7+rTIywLKRZzNjN43b5ONWLCQ2f9xLwEvAS8BLwEvAS+B8kIAnLM6HXvB18BLwEvASOL4EWLCyAGfRymLedrczhwPumusmFqWAyCCgnA8gZ7tnAZUB6wAyWcSS+A8wFwDaQFvKOq4D8fO0s2g3YMV7lQFiASYAPFjcA9gBOABeIRMAKwBrjgGUcxwXCSRcvQD+QFwAlEHsAGoDVCAjjgHu4VIG1zKAEYBcgBTU4WmXAPCVADgAhQByAF4B9ABecDkDQE77DVhEdvQBbjzQNWSNPgIwArDwPy5b2GGPbDcpo4fscMUHv6XjvaOwS5S+O1HiHgDjnI+e85v63KaMbtB/9Ot80NUIQurQXY6KhbuXPDfOx9Vn1sPcdc1gru+X3nhy/6uCW7/1zIHvXJ9pNrv3LF+5u9KfazZyGbe3ezAj8Hq2nlHQcOsKOx2WD/Uk5x4tPelZqpFkwvsrz7xp2nV9uBGGD93Ue+sjxbgWV6PuZi0IlTPt9ZwDfLHL/Y++/DtHwsLQqEsyT2S7RrqG66vHdpQv3/ZE+Yp9q3N7D6wvPHFDjywt+jJjA228jBOZ8muq4827cysfeNnkd96zrjYslFm2FMcSAZF69jXC6h+Sq6jPBdNuXJYWxIH4oDIxLOjLE7n24jwyfW+WF8gZkgsdOZ6LEvSI+c1iNQBGz/Wt9aRGAMx9RJk57+vK7HZmBzYk1jE703/pC+k8ii6bi6St+k4Z7GLe1oopcjRKkqXd8omFOyDiVJBLQb5RCdXZ81I5zF+6L7d87YdzL01uHPz7tF332Ow791zalW804sFmHPeVKvWkXm9Oh2FYzGQzUSZc1x8o0E4pXHa4PvCrO5blrngiqu4+2sitj1eMv399tnn43bK4UBFz1Nisi1CwP1UGQAW8HBKgX/+z5WmAbZ4pkBnMaebCa7Zm0819TiSFG8xe41bmX4Dcp7aX/v72ZlIdkb7N6ScBruaqBoLxhqBRXRU0yrMWTnFxqeuaKruNuw67YrmWEj57Nq509TaxjQ30uC+97FlHr3h4z/jg0fGdimvxeYH7jE/GLfOykVroijU2/ZwXtN36kLaz+/w25dcrdyIreG4yhyMP5gjSc5U/pEw5EFe0g7niVpEVORGIq9TfkyKqXjCUHVipCixAgiSfV/yJx1TyXWrbN0XWVG64/T4jFwCzP6dWHHGVpClHbs8O7o1/uWe05C67vOJwGfW53mPjS+9bseKFxa7KdcsOj29dUpn80MjSvu3jv1DZL3dR7TKZ7UP7cppB7Y8p5ywfYAxBRvEs/T7lhcgKnvNYlf2jMu2GpGBc25zIJ88sdIf3At4BIDdw5YRLs/kJQuttGuN/uKo++pjc5CF/xgvPf94leC/oyCC1CmIO/Cdl5grqg76iLx1Jyg7373TI3vt4eECcMB+hy7QJXe5kWTW/HIuZwzMPMoY6VT1RcZI94E/zEvAS8BLwEvAS8BI4pxLwhMU5Fb+/uZeAl4CXwJMSaFlSzBcJi1ayuS1i1yCAhwVrNddO7P77XmUCKgK+s2Bn8cziH5KDxTvHd7V+AxpbnAuAp3Y3BRccYdHavYhbCDLBM5EPcREgI9rJC0AiZAMQSTsB2gEmcA9EAk7kGCAH4Ca7eQGr2F3dTlIAGmR03/PObVarHYv60SItUguEltwAlPiO7lj8FI4BiCAv9Inv/I/+IVPON5c46CX/82mEAe8k6Ch9gVwhlOhHQJ/5/pfu1DEAViPr2ttrfcoxgFgy98FPOaAS9QTkxoc3CZAawIsxYrFGqCv3BqRdWgtz+b7G5CVTme61Crh9jC+oG6p31jb37VoXZpL6cLN/6rHV65Y08tHgntwKYhK01y39TqyKTQqEPVZd/vD20tWXKUjznPex3dVLVw/V11S/M/299Yde/dwUGH7Ph8GbOiauzbznw/8tli+ZDJ3U35OPc9Xp+u6Se+T+eLBPdcgPu8wTy7Ij37q0ePcLFB/jehzatKXlqsPPTIWFxh3d13z+Bnf/Y2vqR+9X3AZkBCg4N2Xcr0fXuRsUF+Ct8ZDGTOxKjbsFCjZT4PYvlH9S+ceUAe8AhDvtTOZcWQe4/1/5z5UB/SC9LBaKAdR2b/oDggK9eIXySxeQB6QkZCKBbiFqmesoszzfdRHXt1y/QMAxD1AmEdHZ/c6O7Jcrz4Lu+p760Ye8kGycwE13Wbj/k1Nh8VC+Ue/ZlVv5xvl1ktsgwNWB20d+ArkA9M8hmmRh4cqVekaGdJlyte7qzbh/cqraL7MYBbAOXbXRONqVz67JRGFXlIm6q5n1+Yn8zw6H+UaYi8oTUWP47sHpW96Wax68JkgaAmQ7Tt8oIVYmAJ/0593fU3588p7ipbgN5BlC2wGI56RYPOXO8r9sL0Yrl4Que2hp7robm0nlg9932Q+lOonrp9YFjEPGFDvj6e/rRFb09ez4UqO8bsZbTbM4OGMeU6u7volpkRZmKDT3nkeX9S/9zrO2KtZDON49XR7e8viB8Re+9eH5FgQLPqNa/QkJw/MP8gzSAj//L5rfvtZvdATi9cvKX2nVHz0w6zt28AOGp6SXiKpNIiy3PJpfd9Xu3KpD+7NLuc+cJP2AfP2Yxt0X9AkJx7xS+rHX3NFe7ynJj7IPafysTKruaNCMXVeh8hbh5X2XbKi6Z8gq67vFubh0KZPPlgbyS6YLxR9dMTS6Zcflaz+89aG9XxNhgc5zH+5xIVpcoF2QDNgAACAASURBVEOML+YF9BILoU7pX3SQZweZa9C34wWWhzzA+gILA8hrSMxORAjWHLfJii0UYZEtJLUDsjRDN9Ah5pxOCcMvdIb4QcxNEF4QpDzTjrGmWqCMToeZ6xiT9CPuPnFbtUvZiIs5MWA6FMBzlmeduYDiGZ1aLHqy4hR6wZ/qJeAl4CXgJeAl4CVwTiXgCYtzKn5/cy8BLwEvgeNKAHzHCAsWzgClLIoBXwFQWKSzy5xFvrlAAJgBWGHBzPkAhoCFLH7Z0QxKBAjLjnOADdu5Cohm1hXa/PqkW5zzvY9E9BjZYuA1i3wAb36PqC3sFE93zgrMQk6XiWgAGP2SfkNmjFtQbP1Gtv36DRjC+QAV2xfw/X5RkBXW/y2dwNpi1oWN/uO7ucFCtpABfHIc+QCSQATQJxAX6K0RAYB1kGbIGlIBYBn/3+g0+vv9dIEyuso1XI8uAyLTb/i2J3bJ/PSkOcOT/wDg2N52LI0grABYN7XuydhIQb4WCMv7EaAQ94T0WiYuYs2DvVeX7hm4bo4vG1kiNF9avM1t7d7eWy9komY9OrAqGR3cEazpSFbQJgW4/mivK+/pDyY+uza/+/v2Vjf/WnsjFHvipVPNvnVT5T5cJqXg8DvfzCbfY5OIDIslUhLInZdTq544SXKNak90ZTPTn80UHiwFwX3j8epk9/SzM9PNvlueN/DZF2eD6n+fX5oA1lcezfR+Tju7qy+ceqB2RXUvO5MhFXB3Mj89V73yacW2+BXV8B7FC5hoPqw+rM0GZL5dF+CmzcDwhYIboyu/pIzFC/0A2Eu76bPpbz73Svet669ApyCWIGWvbZXbUR46CDj5v5Vxf4LsKKfUydd/az5gPkSfsP55oTKkA/PmQhY8Bjr/sfr+O6vqI8k1wc6phwobLhFQPSAZdtLJ32rV5xNyOzOkusyZOxpx0hXH8ZKpUn2Vwsasj+Nk+VS1vrrZiONao1kt5epru4rZZjaKqmEUTOay0SGRGU/I6uJAUHjjY3GjcnhV6SOHItfQfBWIaFkQz8fvfb9cV3Wtrx15YHt+bUNkC3IltkOn9Bsuie8WWfG2XNj3DN1vmywt6McjrXFCv0AOMOawRIBIYg59QxA3XXHv3bNl1vsQp0poNl2PLC1kPXGvyIn1B9csbQ+mnJ5f7sqzm313NZ+9YeT6vi//6X1XTJ1CrAbGLiQFVjiYKCxEVFjdYAIhqG9TBmxmPtulzLiymBgIdLoU5sP7ipfUFM9kx4786ssVjB1LoWOSdAASzshunkPVn/+Lm5Of/+ljTmXO4fnEs3wv40g2S19N9rqfc0PxS7at3+Wym5vu213g4XOT3Ga5O2649lkrxkZ7Q1nlXP7AnkTWKNtztXoaj+V8dhOlMTC/OegRRMUPKN+kDEBPol/QLyOJGdO4teSZAsHJb/rrRAQN7z08Rz6ujL4zDo4hu9VvfzKa6b1NcWr29MTlB7qSKs+ghcgKrJXIEApfVIbkhCw/E6Ki3aoC6w6eiS9Rhkzp5M6qJabZDyMq0GnmMOZTZJSSpJ6smC8u/9tLwEvAS8BLwEvAS+B8loAnLM7n3vF18xLwEriYJWAuaQBqbfcvwB/zNqAwu4gBVFggk1nwAwCzsGcxz25CSI5dyizo8cMMmQEgTNmUA0hi4POse40LkKxAT5CFLfYNDExBDCxX1Kb0e4t4gKxIkxETbb8Be2yXPf/PnmvnXOyfbfqR6ozkmwa5VTZyguNGXvCd/43EQBchDtA/9BpQhesAqNFbiAR0FwID8AUdBfjGvRegKOVAPqHbdyhDOlypbGA4VjAA0HyyS5dy0HnGBsAg94eAAIjc1LqO+9vO5HY3M+gTY2t0JDuY+8e1/6F6oLDmWeOZ/lU6lqbINWvK1UdyWzPPyn5z9WQ2O3Cwe8lqCSPsj6erE3FXRiAnYzjRzt3vShPjXFK/uRzk9jXCTN3lamNj40sA5Tqln9LBRwr/Nraz8sMDcwA5kRRGZPKZAu5RGDajKASY6ytXGt2ZTNhfjOPBYpyZLiXR1GiSi8fjDf1PlNfJ837tYzcO3nJEADtkBDKydInq+EfaYfyx23qvfXxjfWh3Ma5+VH8i8/coQxa0J8ib96k33xVd7u4MN7sd9Y+nsqR/blNmnqL/6St2NUMILJQA5UjsIuaeEK/75UbH3NxRT8Y5zM2xCO6TpQLWIRNkg65Bys5B8Fu78CkL/WFehCyBTGOeRM86kV52B4JdsHuZfjvSG5f3yxql65H8eulZQF8DqHYiAP6DjgOIPyrAlnrFchPldu0fzfXKhKJSb/TKDdRKRZsebDTjvnK5tiqW5UoYBFn1p6yOkkYhn6uHTY2XJF7SVSx0K7xJVyV3+dCugXdOTRWe/fCmyT/+/Wzj4N+GcVlmDfHbnxTJnG+vUr9P55N6VYHDc6FLtskKZFan285kvDTqyfRjIit2yuADi6bPZ+Io14pTwbMGayhIAUBlCAvIAcZdmsLakyF9Gv3rUjdQUOGZevPg5icOstt95/Cy/ivlFmo+KExZ9DHkE/MC5ORxLf/UpzYmmCOoF3rEvNEpMa8w7rHo+oQy8w9uc2z+NysYsypzcqHF/VOLK2X0A3Kmk4UX5CPnoq/o1ARWNb+8QEV0mHs1JVPG7mQy6T4V9LoHwr7k5flsrXrp/n2/2lgXbb1vnqWFFTc0sGTr2uyRdyvWzX8JaglkGXKlj9J4DucTSN2BqKAZPDvQJeYM3nEgJc2qaVaXWu3FCoa5hPGD1cAsWSEZLyxhDQbdG0sXSAXk/GllyKY0jk97mgyLN0nW0yIsXiUrqhW5JOWLuQ6XTJZ4L8AqjDKx9kPmFb0vHJc4OUGcCupisbS4D5Y7WHlBfp0ooc9YlDFW6HfmGYiKdAxz8QXiEuxE7fT/ewl4CXgJeAl4CXgJXEQS8ITFRdTZvqleAl4CF4wEWMAbYcFuVRbv+BoHHOSTxToLUwA3QF0WpSzyAUiwwGCxyi5CQBuAOM5jdx7lAMpQNgAVzwD+oyxAweYFSFYAGNEGC3qKvNJgsLSn1TZA9VhtO55vfJ3q0+lIQHLlMiwv0s+WfqUgXOs7J/Dd3EgZ8AjYQ98BAhqJxif6DKEA8MJ/fAIWodcAmLj6AojEBQpg0X9SZlc8egxqxb0AsgC/sJIwIBKdQOcZE+gLRIaRH+hN6gMegE/AErrCb+oz+YXlL5s+nF/Zm+CPvi01XZTbGm2/fXP3Yz27isv7hoo93ZNRMVrSnKoKBG60yAquCORKZjJx4SOVIATsUjnJxGh92Xgp7n1IvwkOO98lD9uQ/5tyKNIiEWkxH7ClLak1kbqgT/LPyWXQjmwURAK6l+h3NoljgWDNlUMu2zeVBKNqjKI5h+MjpUtL1f7uWwvRFDuIjbCwOQWgeFk1yK78VN/1h14/dgd9YYTFx9rb3/rOXPPngm7fGxTcv+fe6O6u/VMqO2S1S9ncQRGIFv827KQ+XgL0Jj/SyESf7p6uPCIXQv1TPV0rFD78dTq+EFmBDKnnba1PiIpjdl+3gG36f5My2/5x+QK49//Yew84ya7yzPumip3TTE9Uj0YoByQySEQbMNjG2GB/a7M2i71e1t5dnLMX+zPOsLbX3l2WYMMHOGHAgA0YyyCCQCgL5TDSxM65ct30Pf/bdUbV1dU9QSNpJN3z+52u6hvPec97zq37PG8ALMTLorPg7SMvIBsi7V7pgAgJNwjcsXsywTHkXx9Q0nV5zZBgBJ1CzwBfGT9D1nFNLP4hbRj/96lChsWlSiNaLdc1ZHbebwqa9txdmk2jmlejmYy9GIZRTR4ztqJFZWPLdzMuPj1RPooavcWct0fkRraQLx5Z6H1zye95zl07V/70toHSZ29wo1Xk/QOqP9nZISWL/gHp5muLUf3mup0t1Zwsz4rOgvwajWihruXz47bt/qi8Jnodv/obtV3P+f3CsVuYWxA8gKrGQ2XdNbzKnEiLihVle6z6toutKD845Vbnv6CsODd5QXCHPC0CkRgQRpArneQCemXCOpHzBj1MSiupdvu9DOgNwM26gqw3hOdqncB4sm4AEPOJpf5BVfrLeHXOM/M/axU6gOU7x28IBaVttBNZEgeLcFArJtfHFiHdaJb9x48aD9R+8brn3efuiBf6rPpLXT++c6I0fY5CUOWUN6O9z8e/T06MWRPLM8Weo/V/larcaPsxOkaYq49rLVs4i70tGDc6xbyDwGZObObZ9CXt+xdVyAGIbdaYE3lWHJdRy0OnJuKCcz+oCvnB7yXyWqwrU5nhnkey4z3kqdnhL1gi9trJCn5zQYqyXkCacD2Sap8qWWGMRYx3LGsSuVMghbnH21W7zcvO5uKRxjORdkCQ8ZxkrjAPtiT5Oi+U/p9KIJVAKoFUAqkEUgmkEjibJJASFmfTaKRtSSWQSiCVwBpoYTwFeJEHSAVIBATjOxXAD8tgXnSxLOdFH/AEAMbEPiYUAPt5qedcE1KBY3mZBcwF3OE7VqUA+k+Zl9tWGChDuNAn5GKsYgEp6S/bkR1yqOgc+hkYbwt9T8sZlECLuOCK7XpkiAz0uhPQYVwglyAH+G5yqQAcGktRdJ1zAeBMWA8AdsYXXUe3iTuT6LAqoBYkh/FGAvyC6API4TyOYz9zC+DLJHnuBjZhtZqfzW1zvzpyzfRcbixuuLmqPCqOyQthQJ9Wn10KXpf752qzGEaz2b7VnALR+5E7JitdW54UeHkkIKws2pVbxv4HCeZhnQuQCEAefW7hh5CVCW2yIYeA9qHD9LOTbGONML/h1Bfbtx27J+s5cqqIJvwgOtdx7EpTFvpWHMZl2+lTIyZcKzqUjezpZn17WKrtaeZ77xPBE5uwNu1oKPHj//5YZtS+oeei+gsr90IaIY9fVv1D+tRRGD+8NVhv7hRpwSehUaoCTAHfWGfoJ+MDaQEh8VNdrnN8k3IYXFjuK1w4PzZwq+95PSIrCOW1WSGhLjlKkBMEkInZvu74Vggo1k4s+gHKAfnQL4iQbl4GnC9rbOerGreXWkp8HtnFf7Gt4IFG9tzVSuH58dALTE6K2/w/vWMCi336TvgZCAtjKW7a8WOt/Yz/Z+8o/f5KGPyYrWTbXiMIXfmB7bWa0WWxFffEUTwkj5nhRhA1BfD3KgRU0GiGceCGsbxptlfqfq2a9ar9Pbmgt5ix5VFTDrwLmiX/FY3B0qdNSDN0nJBrx8PJKFeJFkFXrhv5nu3B0vM1xobsbZcV5CJEx5Gecq02euCvHli9+I0fCXP9bw7zAy+q7XnBvYXJ2w9Jt16nY7oB98m13NqiNXTT+63qxNXksFgOesb+ToQF4OotThSXZrcP5TTOzGsA/m7eEJAW5EJpCmgWpm/NATxLrzrHlTmC5xTeVpBFG0iathNYSz6rivcPnlfop9/Kg5QctknIItYUyDeuj7dMt0LOF9aSJMFxe2Ly9pBuIi8MWG3CGTJeZg20/vjlN0UvPvj++Rfk/+bafK68NL66uPKq3G3//q7CROZQdmNkoJnBIev2K59lXTL+SG78/oVrMjP+NVoZv01uDF33C61cGax1Z2MOA/SPuQ2RZLysOmXL+gMZeUgVncaLyTzvNxmKTTcjB8iKh7QuH9C8/k/6vsFThjBcpUbBUs4ia4fyvrtxSB4cdMW0g99YkOvo7+n8dkJn0QOeRxBhzFPWxZ87yQ7RFtY9ZIM8aBfPN+SYGmecpBDTw1IJpBJIJZBKIJVAKoGzVwIpYXH2jk3aslQCqQSeeRIwnhX0nBdgXqINMcF3QLjE4lsVAJawGQAoALEA9rzA8hLMfr4D+mLxCdBiQukc1HdeZrk+L9oJsKh60paKZ9Gw0CdAVtrP8wzAEbnQN8gYyBz6Rz+NbAHikEtaniAJdHhgtN8VPWRcIB0MgMd+xo+KTgIIAWgB/rON8QUw5H+AHvQeoMbkLIHsIHY8lrPoBcdwPPfCepfrARZzHPuYKwA86MRx0KkVRqUhoM//4N4f967fdnWj5hSajh1draPQK3fCOTh3aeaueHfm8LOyVu3hyHYOFqImoXZ2znqDF/p2pilADHCNOfg/ZUGPdwj3aJrEy/lP/pXxPoFUAXTqjOePlS35GO4VyNkO0BkCiP5D3lDH6s2A9eJiAeCDfhQpNYK7rRg1s/udytS0kx/KW+HAgJLKFoSGN2avPhxlp292MisfVKQqwk+1F2RG7PTpbxUvfFCEBfMGMOz9rTYCqnX7DflWbQfIg5zA0reJdbfkCEhIhbggLwbW559R/QNViIN1RbGtrHohW5sbGyx4QXiVQgZx7maF+zGOEJVcGzluAOxEVrA24hUAOE44Hzw1sJLmfwprRbciEiKajO38B0RYcJ8DTlSp9la/1i1WPTpGeCFImW5eM1wfvWP/85caD9/oNpfqVthblDdMXvkp5FAR5xXDruk4Vt2x44xo5JyICzeXVQ5uNUQeFUoiY2+XIsUa46zvy+/Cj5quG40Gll1eyL9mMTf83w5uW/iTkhPXDFFtQi69Vcy00HlPVYHB7Ew3skJhm+IfGVwqf/MFN9zjjc0u54vN60ebQ/vi8v7vAFiNGyPn/bA8Iy5U27qFRDouQzsKRFQMTTVHnjVo+9X52q6rbs3N3QthgBz9K295wL/hxZcc1HfCf/E8I4xTZ2Fd/wVVAOMPi0xg/qy5c117fF1nPqBbrAMbEiS0Lsj8Q4+5P54VeCrWNslP1NkGiEN0h3WC9gBydxbahDcXAPIjauOJnjM8v5i/xiOH7ybHj/WNif9YPZp9TvlNg790UyFeyeypzTVzkf+GCxpHdyjHzIabP6JIdXvdWWvMXrEyGWnCTHx5XFUuj1hW+rH1Xp3AfDybwGx0hz6jg4wLxBeeMZ0FIP+gKus6OsA4ny5ZYaE70qGScs8ccK24EFr2n05nhruSBD1R3Vp2e63hsGTl4+gvFD6NZw1EF88PniONdqKrS9u7bTJGKfwuY/1hXbpGFSKb/EwnUwiLxZypRbZbDu3MXdP9l8zuWb4FQuqp+FvuZPqcHpNKIJVAKoFUAqkEUgk8wySQEhbPsAFPu5tKIJXAWS8BQAwTIgCwiVjZvNjzgkwldAIvpKzfvLRDTLCdF//rVbEwBQwCuATMx2oVK3POYRugC4AewAXbEqD2qeB10Ao5ZAYQGQEiUQEA6Zt5+Tdxm038fMBLaiI3XSf1sjBSfAI/2zww2u9qSALjidG5DxDaeE8wD0zIKJPXgDnAfuYDABAWxXxHBwACAbPZzz6IBsIUcR0s4NEJc/0kfFXnPAD8yX/yl+P9zsO5c+2H/cl4Z64c9/Tn7Xppv3cg3u5ON8a9Y1Ep455Xd5xcyS5gsX2PQokUZLlLSJ7r9AkgZwjEsD15MGGeFO7JeJN8VMeRfLq9vF2N/fxY1ID4oK3oPTIw+s+5vfKm8D3HXpUF/pXauTeMrJEwtjwBcm4hDoM9UZ15T8nkrKi/bHujK40dB7dX9szaA9VP2Xajk7DgWMJRsf78juL3z75j7lPMH9YWYv4z1wBt24km1qEJ1Xervkf1/wpQXhKgF7TCbHFNEyqMdsvrRAm713JSYDMPibAYOc5wqb9gzY0NFe67+Bzr2O5RFigDvLe6cfyDEExfVUU+yP5YJ1Dclq8Cbx3CgUHy8r3DTj9ZR9oL6wfAIGvlfbGTn4vtbOAFs4Dcm4GCbIe0IEY+IcsgUH61s9H6/zdV32Lb4fZGUDnihIWsvGO2KaqaKz6iphwVo47nSra277p2wXHFL8RW2Q/jahCEA9LUfD7nOYEYi7rv52tNr6mJ5MV2EBdzPc70yK9wy5nx+d9D1z+mCikDQP/Wmp2zpr0hS6Sa9UAOnmx9UTyxj/StVOovve72PeNTC+PyhIC8+o7hG9/XX9/x7BVvdTLrD+y9WESERcinLcq/yhvj/fUdV/yEQkJdbXm5zOrF33do8PaPMSdDk1vhT/9rQhT9W0te6A3ERbfy09oI6H69AOdG2zxCB5nzeFj8iWp7+J726wA2c++vqDIfq51gcxfPCq4NoAxJgSdS1xBCrZtwXe6RhAjaTC4t7wrjHciaZAgL2m/mNfMkd7h5VfjRxffWv2/w178+7B58WGNzrzTvxwSgX7XobsxhL+DdGhlftbxRsVx3162IVa5s/ZiyDC3pvHdr9uVEHhoy+AlNwtwhW7OGsTayNtNfEm13zsGD2ga5RE/QkeMJpI18T5C7YsMwJOvB3KeQf27J7c3OewP/+DX3svm6nfkdrdsuHkim3FY4z7qq9qC1FPbdvy1erjlxgBdXEjqQeopkhTGaoM9UjCogTZmE/10VMuayzfQm2W67PFPykZv5ct3r+2QtO1Ja6jmneWz4ubUbx74vafi7Xn6c8F93qXYPny3vke5MJZBKIJVAKoFUAqkEUgmcJRJICYuzZCDSZqQSSCXwzJVAC4g3VncmvBFkA+AX4AcAG0AsZpW85ALAQjoYoA5ACStlQCmAPV76eXk9qGpeknnJZhshNgBgAG5MRtTTCWfwZA6YCZnFM4xK+7HChLTBEhsUDYC23YIegNsk434y257eexMJdCE0EitazQ8DijMf+I7e4jVjvGk4DOAa3aYAnGOFa8gswEN0A2AM0JbtAIPoA/U4adKtaW/MfFo5cMvjk/GOi2fjbUmb6nG+79vh5Sue6399IVe40HPrQ76dLYS2uxpYij5v2feoArBxbwBs6jqyou1exvujK/qrxvUvOhnQSfptPK+Y85B0yZyWw8S2ILaGozg6T+SFrPftITW0qdwHjiZIRp4ezawVFxuWcyywHP63anH+Zn/2JSu2W7vN6zvwP+Vl8d+69J9QSZ9UNV4LtBUrcuT4j6oQDiakFCQGBTkD0gPYf1UA4UoXK3b6AflB6ByIBgD+Nyrs0/Mbucy+uW1Dly4O91vl3kKSqHmTUs/4wV/IG+N2ncd6RgiedXO8RVYADiKrc1SfqwogTqz4zsIaaQDTT+g7/+MJQtz8ZTdcNl4bcZccChZhilogOuGLDCH8rzr3ZarkGOosz1Zmk0m798H5eHlUEZ9sxYRyFhWZbzGS5berpOlRGG93XIV68kNvtVnf6WW8iuM4deWwEKcRR3JEsYIwHqhUg+2VWjAnj4wgN9rnV2rNWKRFKMICfUU2EC+jAmQfWHWL5wuktQ5k1+czVnLhQOFvVvZPT87vvnvm+dtnFi8VWYG3CDH1t/U8ct0lxUPfKPj9O/KNbRfFje2Xhd7DX+p8jyAcF88qrOE/7tZX7aBnmx87bkbeKX5l38t9ERXrvF/wNpK8IBBYuwlxsxlhcbn2YQl/UHX6m9+8qGFV7mVe83zk2UgeDENWoAftCZUJ1WVCkk1qrLby2GkfJ/qHVwkW8Fi/dwtbxfHMETyp8K6gdg3J0yIrjEECugZJYfJmMMd5bhmiFTnWZ4Pzpt83/3fiNn/1wM6eb/6tE8er2/2l7xdh8T3tDeW78lxYU96w9bLyt63d58+J/VJ+djSxZv2MrtqvVv2/osOYy6wbgciL+pNkkY9cGTc8jTCyILcLxGVnMb9zkjWnfOevmWdAcpxA+FP67dLKX2MIqIxyDb1Q+We80WC172hm1P1a72WKjbm+CQ9nd4S5KDgqb4vJwbDMeh6dIlFhSc7ckz6jr5DAJiQnayYkG8V4em2Ugu3Mah38lIi/j0d2drBWGJv59rk/tjA7+ly75A55NSvj5fxQXK8d1eq+kVF8qvLpIv90UyqBVAKpBFIJpBJIJZBK4EmTQEpYPGmiT2+cSiCVQCqBDRIwpAUv4YCukA+AbYAYfAd04eUejwlADl6CX6HKSzQv/hxjrMY5B5AOK2HAXD45HgAAwgMAH0+D0w6t8CSOnwkZRBP4Tl8AqrCCpY/IDkAAcAA5EGYHy0yAIIAqJZGNm08Fr5InUcZnza1NbpU2Fwx01oSTMoQc4wspwO8aE1OcYwyAjd4DinIuYD96YkKhcQw5XDZYzcv7wem3PjK8zZlrfst/3pUiIcaH7KUHy1bveK+3fPiC3lv9nN2MbMU5V16AIe0n0S8hZ35LFYKBuYlVeNVYhOuanbJFh41HCKGu8AI4XhSG5M1ubJVu8IaufWGwZLyr6CcAJ7q9U7LZp4sArF5G7nNyIOj7uEL7KIyQE2QEb48rSXPJdgeFVNrFKFwZjP3zonDo3qi6p2L1PUxuCdpuEmSb+7PWEK//IXlZHKEPAv3oE4QQ8sR63xAW7c1GxlhMA+K6OifJS9IB9NHvisA85m+l0pP/UqW3EImkOHronO37Qs/tWR7qNLh+9BY7j83foWO22VFUnt4xsi5nRVuoIMaZPmHFDDj4NtXNcmFwM8gTPNX+UhX9oJ+MDeGfTrq0ws4k+TxU8UjpRlgozJHtOj0PLjfmrxIrlw3zeU/5Key63wwD5SKpycmi4Dnugu05g4Fi12Q9JfsOI6/WCFxRd0M9uaxSXEQNPwzPUy6LVQGWjaYfJnmLevTkaMmbMVtUkm2pkvXOpu09Txb6PyeCQvGQHk2xIRLLe1H1nhGBt2/KZRpT4onwDkGP3knH7aBpFY7dZJXP+1Urs3zIbg5NeD1KSizVapcL482cpA2HlLPinrA4zDPqHhEWy7GX233bkVX7yj3964Bmcj2ItGCOQqz8iCo5KHjWdeojOTNuUEc+nxWILAKm340jxhVwH1LBlHay4q9b4wmBZkKTbRjLTbwr0ImrVOkk68RGl5S1nC4kPma+4wlwfK5vuMkaUcAznfbCGDFPDJDNMwsyFdkxt1nHKBgvTH5y+fcrb3Hevrgj9+3PnNOceUiERbDk9b5GYb24xvEiQsq6J7/XUhJ4a+CyiqWQalY8oxVhwXpbdFQyakq/IxGFcWLRf7PmH8ThcY+XLm0+05uQAesW6wYkEGHAIKM6C94Ei3IS+1ZU3/aQv3gl8kdhje6cTugjfhMge3JlIN9x6dIvDGjKKAG9ZK+63QAAIABJREFUstr71hf61/MmCp925LbC/sn787tX5X0RvfWqL54SSSL5Mh8gKegnYa8YY9YFcrJcsoVw+Z32MZF9cMwK/lY8XBm/cmp+/IWPTI2/JFvvn+gLa3bR1cox6NjLy/Kv84MwzGZcT2sA92yKIEs8S1Pi4kyrcHq9VAKpBFIJpBJIJZBK4ImQQEpYPBFSTu+RSiCVQCqBk5MAL+CGQOBFk5dcQkABGgKcYNWM5Sov7nheYFGOZSkIKMAS5wMich6gJ8BAEupGFTCIl3UKx5sQSSfXsrPrKBNOgj4jgwS0VQXY4SWfMAuAEgADyARAi+3IwoTVObt6lLbmVCVgSKt2e1jG1hAY/L5h7DkuCf/RGn/jVQHonlg2b0Xa/XruD71qXNj3eu8L590ZXhbcHV1k7fUO3Rh68ZU7ckfOjzPBRUfd7XaPu8p98PgABMNbgPjieP0k86w9DFSXjhpvA5KHo7s/YY4BYVZYp8uKVjhYtV303eSS4LqArxOqI7rATse2d4u46NP3jMJBFdT5gjwqmPNKAB4FWXEySroN7p3PKWGCYqMxX1x/+aJqZvSGf7O9KuAhSYM7C14JVEjPOuGQBIAzn1iPAPMhJn5btTOcyb/XNtr8d6p4UhjCaN31sfAWWBzmGv5iodqo7JhaqD9y7k4vyHTmq147radSty6497A1vLCSObRvx61X3Xx/NLyQyF9m5MfzGgBYsyYAhBIXHwCY9m6VuJs4/4Da6AVW8uiTyfHTKZMT/t8C4Vlrldg8Aal/a8NJsfWzdnZh2S5MfTFq7olrtWCHPCq2RVHsREHcE4mxyHrRiEgKjWucr9aa6HFT+5uBH2dCEFbpnBJfrFbrzXkRGeV81mvuGOsz634il+bfWtHtrzx3JT/k3+lnvOfO5IaWMnE4hDKZ0rAzVskpWkMD5T09o409TjF+vmimo49mdlHylns/Yy28+B1JKCj5S1iRl9NnchXk9QFVyAG8Buj34cq+lzZjN6dxt9/QkkH7c2mdOFryYs6QEJvQbVBE5K5AEQDzTfmZXNS8Y1uwNCoAuSGdZkz/vLUT8N3ESoIoRC/RBa7LeFZO0jqeZyeyRn6Qoa9V3eDR0LqnIUXxZKmpH12BdIHHXDOjfCS9Gj/IxXEtVnmtP8o1I/aIdscxc5m5ZfTVeFyy/5jCQyHspR/Z+903KVfOn4h0OiyPix+uO1kT8i1p0oHcTuvK2gGr7BSsPq9qeTtFWmhU4kaS7+q1cUnERZx4nKAnkCwLAtbN74I2UT/6VfP0TBXWY/SAuYmudCMr8Av5qFZnNdxeDGvjvr/4bCPXLQH4bt5PuhbPBX5DQRAgK0g004bjce1Yb4tRQwnpEftaqTj5CX1MiM7gN8XbtVYd3Go9bxEUnMp4oz8QSniqfXdrG3oEWcRav1mBgH2HSL49sZevBv07D5f2XD03deV/aMxl9nrlejDSDO2imhnlI4X/ynjFZhg16w17VevCCuuH1gzzbGz3ItzilumuVAKpBFIJpBJIJZBKIJXA2SWBlLA4u8YjbU0qgVQCz1wJ8HIJuGjyMACu8MLLizuADcSFsSzHMhOgnhd4k78CkgIwg318B2T5cusYQArAVCrHPxW9Kto1w7yIIxdACGQE2AL4YWQIcAzIBWAA6GjkC1iBDJBdO17Xfv30+1kogRPkwCB0lNFrxprxZf4A1vBJZbsJv2LIjC17+rf+m+3Xel+85FC0d3zAXr4ntJyBY9HOFwsmHi64FcePcpPFuH5zf1SZFDh4VF4WgGCQFehmYJJrt99EsV2sLl4WtAvw/6A51ii5CIZ9IhdWymvW8Pwx3iEcAiHAmlFU//uV20DYp5WT0vfIZSTnaQMW8PKwEHOiDM5xrG2xJwJE2yI8sMZjf8CvPfyWamH/h8WJNAhh1Jn4lZBAWLt/1eQOAPQVMGhCVEFykBz8b1QBYtsLZAbtZD2a5ZwueQMgTrYpFNRLVN+8Mti7T0bDjyKGbVcbXly1Lr/9gDWwXI5G55afte/hqV93wxDAFbLhVrw1Ys12uzdZB+kfcx+iAuCbkFCblc9rB8QCgDfgMGsEhFDX0D5bXKdzF+N6SJWQQb+14TwlprDc+g/kRm/7djA9Xoqj7Kpr2wuO3Cr8ZpSVl0VWKbbBUYVL2zX9b2mfrx/vk1LgUq3hK5KUpWAwMSRGoLEPiwXRU2gB+PSadbezMDqQL9uFXQcKO98owuJVpWyRtXJd2d+Ysi6qH04s893tkRWdo4vdI48CrtSaWZnVKSs/dbtVH7/Mqu55oZWbuevG/Mzd79MRrMGAsGYtTkKIjf/nv4pvO/JnJBMGtGVtBjBGh7s+g1rhoRgzvDsgyBiPv+ho6nDNyX363vzezw1WKhd7cThBiLNWMWQF93yLKjrAXD8gvTvZ9R6ZQTDx3JxQJXxYtzwk3BIDAogRCJvEE6ejrcm/7WSF/h0SDwWxSNsKulm/o+QoYRx78tCSsby1qNGraj7zHKf/tJ85n4ylavyxw//UHL/kN++Sd8X+yLLx3llHWHDPz8tT4Krqg0nC6D3+vOWSXrpPuaNn5InI1QL9pggtSMU/UiXsGaQOusq8Ph3vhW5d79xmiAPky706c/aY48lvs6wl6w659ixmhm8LfvEV//2UPBtaFzIEtiG98MKEyCT80vGYaOiP9MjaFixbL6rcY/1bH44QGwprGLppdfHGIRwcoZ8YH+Mxg6EJkuaT+2JcYjx0ICvQnU4CFQ871jN0arcC+j0QZXsfWD7nFTOTz/7xXG1gYqxZ9ntqvj8sbwqvr0cplcRoy6Oiv14LLeW7Cfv6s43FlTAUYcG9+R3kSf9CeVk81X/3nYx+pcekEkglkEoglUAqgVQCTyMJpITF02gw066kEkgl8JSVgAEiAO54yQSETywwVXlB5gXW5GAAVODFE68CQBLAQt6uATcMWANAxwsvoAPbAFI4z3hwJJ8m1M5TTGoGgKDZxsqc/iErADG+AzQhI8AeiB3+B9Q1nijIlOTbMkrfGAbodOXRkRTcXMbgzp2XPQ6+bALEn24z0vPWSCrG34Buxtoc2bTLfUsAjLBCL6qU89NKI/D3wQ9M3B+ef4VrhWOL4fjujN1cyTvV27JetV9eFn2rdnFFYCMAHHPy4ZYebgr6QVp0FCX3XmaeA1itKyiQYre9UMa0Ny/amdpw7AOKGRDTkJhs61/zsLCLqoKxFEiEw4R+CpCT/Txhr4R4a63IxvFlui7957xGHBYndRC3IgdBJ2FBewBFCRuVhHZiQ8vTAnATII9thFPqJCw49I2qWAwzHx+UXI9buQv4Y81jLYOQZf5eLrJiYzZh7dg+vWjtf2gy8bAo1BqOQt30KceCCbV0hVbO77GLitlyvxW5l4qszGjtdJJ7klB8K7ICrwDGDvkDuLM+UB8zaNsKDWVyEhCrnpwf64qi8l0e54+8xitO/kNU3cf4C7tOQvUNabRyylkxbTvxtqgZyzrfbmrAlCbFERUVDwdBXJXFfljMOfmeQnakkPfmBrxmdvzadwZ7vv3BNQ+ajNezNNS3c2b70EXlYuEahdFaZ9mtvBXWjmDR2h4sKbO3KC6pBdXRSEYHdQWiPiVBgzTmkW8VD9/wQG3383aWLnh9EOYHP7X7E/+BcEj0MQkzaKpJqq3/IR4gy43XAiTbpkmp22SGXgGk84yDNFtXlDD8lTv9hfy+5kwSzqet4J0BgQU4zJrPfNz0fp3X1f/oIaA2Vvi8J3UL58VpXPM61a+27lPfzPJ+ZLDoCGAuiFgaUrCvnfKi2a7YXgoxZ7kK25a3HDtwIrsugF4Da/kakpqUD5nOaU4zPwj5yCggE0ogghSZXquxWlL9C43aunBV8gywvt57qTUh+RD+CzDe2y/SQj2KFOhMxIWQbl0hVO6POHlOov8QPRg6MA/OdGF9QSdp58tU/0uXG5iwWv+mfV9XNaToCdvSxbOC+/F7CnKE5/+rVPktQK6TdoIHvS3IU8fqD6sKr1T+tMiL54l8RgfaC3pwtSphy5D9unw5IitMmD7OI5TZK1WZa5Al9LeTVOr0sEBvkT3jfLPCp93UGL1gcfLFPx8vbntebsnu63Ma4W7pSF5LdY/0JFMqN3cFUVgVcRHntAY0/XhAOSzKWvIbGc+by2WdqXK1Sf9skRZpaKgTalF6QCqBVAKpBFIJpBJIJXA2SSAlLM6m0UjbkkoglcDTWgJbANrGAtwk6MUadUKVEBPEUAcEgoQAxCJ8AgAOL+C8+PMybsLf8ALNSz65LowlIy+rgG9JssiWgJ+qZAXNb/euwAo7idWvCkDAPsBOwBeTlBkkC/lQkRnAqQGwNyMTWmJ6zB+GiDLtNuNkrPvNeJyO5ehjbtzT7QJdiJ92uZ6yjD/hf5/zKvfL3tfCFwvqG7xwKh4/L28r/QluDJYT9nirh+txcUReF5qnMXMVYBHQCcvZreLYJ6Lv8LJAV9BVQhIlABrHsDAkyqO7jkbNvFwgKiIs2GTCn/EPer1TRvUCseyCOppRBPOc8l4k+QVEdug6tuvKA0VEhQKIQIjGzB3IBdr9UBwUM1FtfMrtOYQ1O9bN71dtJw6YUz+k+ohIBpJbJ/JseVrQXoBhQj+dp9ot1Ak5Cf5ZFcA1CSmlnBj0GaIVS2fWMgC+rmTF4FL5H/YemlnpLVd/vH+lYvWWqmIm2obUts4XEPsee8C6XiDsimL1zzgTSf9MQts1Qa4vrK0fUr1XFe8ASN0kObrqKetLtxuwrS2fxUdb/Xzz+mN1K6f6Cit/+ON+aediEGTHPc9tatAr4pmO1RXmSbqd11FDjrxnlLPCFnPRm8k6ddtyG7YVlQW2HstazWpvZaa5/94PWIP3/d0+3YN1Efn29JWqPbuOzi08vH9n1MxlWDOPl9G5Fev8+lFrYKBq9UY1XDmSffJSsVxF3Y8FzcpWe0lPkLfGpejcgTs+tqN6zouH6uNXWPUdV9zeHN4/n108QDLtzQge2Dnj6YRFOZ4FWwLibaQFZMf/laK8Rq0irNTxIkA5/2BuVwLG72tOK1GKfA3Whg1wn3BSzEPCSwEunwz5xHQDXEYHIbgAywkFRX4kvG3a5QZ5d6MqZAV6w/O1q86QaFtTMGfbTq/yqvdKuc6TC8wlAp2Zt57t2srTkMxJT+NeFsGoAE5RUd05pqFAh7k3ZAJAOM9ySEOb0FPMRa1Ht6jf7xbI/krJhNwMxwvU04w3ZK0ompySS4usUIg5+WQ40o5AaayhxTS+BdW3Set5Nn5YlXXoupbMGm3EU/ulT+m72mnICnSSEG1U9KC90Lf3tGTJ2D2Wecj9GEtkhncYnj0Ql6xjVAr9hJyiEh7r+RrA3yu7hUnJsq8LYcHa9j9Vf1eVtewoetryYjJrGcTrhCohoPgOQbI+u/2jPTbLO1vIafEHqhBG6NLC/NU/X1m+8kfdpajQXw0yu2qV5l4N2A6FfxupNf2MiIkBx3bG1Gbbc/0lKVk1m7EHewvZBdtxFprNQBPCrvT1ZhsiNrhXkJIWjwo//ZZKIJVAKoFUAqkEUgmc/RJICYuzf4zSFqYSSCXw9JeAsZhuD/0A+AEASuHFG9AFwOQaVcgLclgARj1bFdCRwvGQGwCIgAGs8Ybo4Hti/foU9awwWpDAsKq81APa0leToBygCVkBxiIvwFH+53gTDgHrRfabpM3mumfysz0MBXI3YA3fAZ8oWH4myZ5FZDHuJH0+k21Ir/UYJXBvdGH8T8HrdkzF2y7enTkyP2AvAUw6I85cvRr11JeD4aWiW1Ke4whdMjkd8DI4IVlB0zq8LOIWgYGHBha8r0ZpUYyWh0X+iFPYORCLO1nTGxNWh3nAvWexsIZNkYdCAt3KAj+xlae0kFTOCzCYVzXWwCaMmhssX1IWYcH8ACTtJA4IocL68kFV2nDcpL1FWqDXJJdmvXmX6ou6iJ8o+ISIukfW4TSJNgDoAa4TUgoQs1u5s1bMfWN2+9DknsOzUd9qZacbRq9PDmzZUNusBEXru+Oa9Z2CgT+n1u+RhLrFdUEGzL2Dqp9QJUE6hAXjRh8er7Ap6Ajr0UdUAU9JwLtWNE62E1wQFx8Zs/MT1ai6a1KcRBImS0tDLQxtgfuRIkE5jpcV5B0pE4Gie0k55rJu8yHPr9oDKwejkXix2lObahTv+/w+x6+SQP2KyLE9hdm6XLW8+8jc4Tuv2P/STgHvnJy3dk7NWeGFnuUp9UVbeCVLpE9SnLJyIDWs3eEj1tecaZls73rulWF+4JVWz+hzHvqvt31JSbS3IgTwejPAsAGJO5ux4f8WaVERIfH5QtSYaTjZXXU7Qy6V4+WQ0grgSaB8HNYufz7IxAEEB15CzKHrVHk2+ifKWyFA3RAVgNnoPs9Xsi+/UBViqyWJ5NaQisabik/IccK/begDZMVAX95rNMIeuc305TLOSDMId2ss+7M5b7rRCLYryTr7ehSqLed6IhwDhXez7TH5XngK7TUvL5s5qflDelDQLrwv2/OqoFd4d93eCke3oQ3kY1DoKKmLbUmGa94oLACSZKyRoYaiWTV3xvRU/HEtFiTDhnwERL9RgPycSIvTnhctsoJnrgmx9QP6jrdDZ0FPWF/IhQNhcSpeMeZaxkjAhCAzhgzMc8iy9oesyenFtg+pfkxfgpFg9f587H9IOSvIufPWjkZCuOApkR2bXfYkG/Q+IZ5UITQwKOE5AWm7Tldb1+kkvljv/14V/eM7+ro69/JftSoTVzur2TFnYbFs+816drXqi3OOilrZh+qNcDQM4mxkh4NhbEeeJzWQV4XOzalBo5mM21BIKE9ePAotZpWViFsZuUPzO3Oj5NMtqQRSCaQSSCWQSiCVQCqBs1ACKWFxFg5K2qRUAqkEnlESMC/YvLACUlHN2sxLLy/5gIAAFSasCkQFL/QACpeq8oIM4PZdqgAuAI4AgliI8uIOqGESap4xy+EncZSQFSUJddDqPxbaADq3qQIUYNWLfAAskCkhsiZUAWgBRpDD48UQGOtOZE/l/tyPcQAwZXyxoKcdbEvA5xZxYQiZVhfVyJTIOC6LJ/LL++Mf9epWz/hgZjG4oPe2hVsqLylVgr6R3flHlutxPr6y74aL+9wVQHzCl2BtDSBN0t2TmmNdPCwA0NALkm+/2vQVlKlpOa+ZdXLXxWEJUMroPWsCAPCCwMglQc013bih4xPnCgBKUlgk9IW4i7X/4kCfgIfEVUcPITYT/VRS2zC363MmqTckIEBce8FimJIjl8XLhjHGTnTXllmwImNNNkZWPnLr6PL7f98Nlz+joEJqAUDaWoghtQig738p7NBvz2QGjypp8Lam7Z2rvT+n7Vi0m3Iw6fKaVfnvcw8/48Y7j83forBQhPchpMsjuug+7q4MD2vMjlY7eQVMOaPWGx1mffcCWYGnA6A2niTkWuB+5ROB2pte8SR2tHIzAKZ/RfW3VQGEW6U1WrmZ/5wb+fb7onhs0g4z8h+xB0PlsPCcOPCDaCWw4qNWEOWUjFvocVR3msHMgDWzsxCslnbNXn/h6MLt+/sX7ytn/VKvxvwlAr0vVDiooaN7ttkPnb97dHLXyES3pgaea032jVjDkyXL3SNcOvHtWV8k1/NEl/+oN2CVIz//uTDX9zodAQCMvvA84tm0WQFgZ92DDGN9PunyjrlPRVOZ4ZoSgttHsmN33Vp41gYQeF6N0jFWX1QV31J7r/KQm+cja/66WFHdbixdRifQGIgkZASZBEEH6Qbx3Znvgz4AZmOV/5DqlnlOshnHqchtRrkpegUi79d03KWx3B42/F1hpGZHSmRvR4OaInllIZnSeu+JncJDalzM4oFAJvWEktJ+FIW5etwyv817h3ZAvP2l6ts6+3ld7+UidnKKIVayz/FnLRFAySG2Zj81YhbQ04Y1FFfV39i6UP/9mmqSQ0vAPLrbHmZvgyi7JeWWbGkrz0BCenFN5m83soLrAdbjjcBn4om14SZbb+C5y5rG/VgbWcMglzDqIAdJt+c9awwh4W5SnWedKkTNBZE85FBBjyBY29dBrv8zqu9zoijfzGYy2aaPTiJQCFeIQp4JneGkTMvRNQqyhAi7XvVzqpAV6FQJT6Xb3vmrtDWeOrpoV2t+VuHEcloDBmTeIP8YcZMKIyZyqx6G0p84HG4046CQ8UjYPu03g7piXQ4Xcpk5K+vV/DAMXd9ekF7NN5rBY83JY/qRfqYSSCWQSiCVQCqBVAKpBB53CaSExeMu4vQGqQRSCaQS2FICxpAasBIPCkgGE86IF3cTDoL1GlgBEJ4XcGAlrEC3qwLW8yLKeQBDgAu8sAP6JTHqVQkDdaoAwNk6dMYaFiAJEBRSBwAWmfBJYRtAAjI04T3YzjkAtiY01JnuoyGg1my+18AOADvgIArbIFYYT7Yx/masGB/GLPG8ONMNS6938hIQmaBxnMwK5S/0ZxbLQ7m5vaPN6eWlYLSvHhfKg978rnpU8AUqf1MgF9a7gE8n5VlhWtEl+TY6gYXucVAJqD+SijRtZ48y0EYiLgzohn6gJ9OiI8ZIp+vb5K6wMjqgyKQ3lvJrzJygULx4HiXqOASwmcq1TPgV1hvC6LDWfIwzk4BSSonhyDEh5wy/dyz7vA/vzL3ioPZDdpBIljWo6Xs7vemRX1pY6nvznYOlT/6CyIq391WuOy8THLVCd8jKNYWpRvXLA9v7SN3OvkuJGC5R/wCF28kKxAPgB9j8ZVXuU4kcx5KHBQAk4fDeqcYMKl/FswXf/rySbF8CL+NoxjvnWROK7r5VwQsEzwoFxEnGjL43Hk+yoq0x3Iu1i3WbdRxL8rWSjKr/MoWF+pSdm34oKJ/ju46jMELxSN6zt2UiH/IiXwjgNWM/9PK1waiUGV65Pzu2eMfubct3XlUoHRnJ+OUiBJXICkuhn6xKT95aGeyxBKpqDAzP+2iLSGJeLeSteM4u9y5W55Q9Adh+X1cB2ko+7Vo3ZzILdzhWczWy8qxf6Cpg/1aEBc8fSHfkDUB8UoSewoaho1lZvJM9w5HV+96xYNX6lz5UTkou0B3vAcqqWySxx7yIsMZQUP64QluhPxsSvJt+taz+kTrPXcht+szFflj1ZW39B7RuLxBd5NVg/PCuWJfHoIvc7LnFakZjWfA8Z0TeFNs0g4tMa82sAdeJBzU3Z/0wXgPalWhbYPOSPCv0LIuHJSkB+HZW55UU0Y2k6sxX5Hjc+6BFWgB4Q8R9sbUPj6V15abiBfZ5jUm5WLrWhY0jSZJpUzylFQ9FwygIWVJEWgCs/7HuDzlzsyoEGyC+yd1wwjFsyZgx5Hl3lSpEBYTdZgXwnjHgmb1lgvSOfBVmTeSZy+8B5pkh0sif82eqmxkn/LL2EUIzIX5VG32vrCnUlodwMAJh3ys6GjwssuJXlAvm05pfseYWZAw6Tn4aE25qsz6yphF+jvGGZLpOFV2tiKg4rkvyWIqvvXPaDoLIrTdFT4rZkitfVrlPvGYzzks/KvK2KPhhJHJSXhVa3WtW0Ced0qZoyXPdUjbrrrqOO6Cez+v/MKtAgSIsthB/uiuVQCqBVAKpBFIJpBJIJXB2SSAlLM6u8Uhbk0oglcAzUwIGMOQlGaCAt0peYgG2iMcN+A5YAPg9oQrAAjAPaPGIKi/pkBYAegBHgDBcB2CDF+kkvraKOAvZWj/1C33g5d4QMvTIEDOEbDBhmPgOQYHcANWQqfGsSOTcEsqZlIkhLGiTCXvDd9oKocLY4VkBekibICsYbwPkGVRx05joT/3he2r0wLFCr89bycz6O1500+pLranmHoFa8aFq2LM6mpl+pBHlr3dtYL4EjF09Wc+KLXrP2AOQQgAkxXhKOBb5KSyvueZuA6iXhIISUdFo2E5Z+xWkPG7ULLdfwV+UozkJCpWgdC2FVzwQLQBr64LJoZKEiFNljTDRpyKREoqLH9zp2sUv5+zBV2SdIavojivYfo+1M//KFytvwmZJiHUZhZ3JnmvNjvzsfXbU6CkVX9EYWv3bnBdK5UW3WOG0LL294niw9HvDYem2OW+A9Q0PMYA++o9FN20BDGZtA4SE8Fs4cN4u8iTE4V8ptv+i5n9Bx9rWZ+Nla9oZtl7lGP+PbgJuWPPRjPUhWZPfbeeUZyTSHMwlRMVph7o5DS2mX3gZ0C/AzWsfvYZGiaXZW/pJe9s/LReb33Xr0Io9aAe+q/AuQ3EUDAeZnrjXCetOdSmurTb8Syc/+5qB6uHzvbBh5cKylQmqusRadyAsavls8qnk5BZeFJ1l9+HZ+kX3HJpxo6g6tLD6qVzdr8iivx5NWXPODuv/69o/GzA//rQdVSctV4yIZeOV8LzbjqzeA8i6iUzYjo7xnILkgjTaUDpAaBrM2tivkFB4Ee4fDVauGQpK1hXeAeuOwv7jZAUXui+3x3oou7OvTzk4FDZqtRA3VxddcPL1YZpaFv88K1iLIcZ4VnIfaK43qbaTFZ1tBLRn7ACajTHBps8OwkHpOOZbn8DmEenquKJ69UoJFKnLXpbnRaAE3EV5T2Q0SUUVxZ6ICVe8UkMW80O2mI1cxh0QRVVV5pmCQOoDYRyhP4lXU3vjWvksMHbAk/JfVTcQFhz/UG6nVXcy1liwklSnjRd35M8ZQr3q6alcMMmIxXWFVYuT0GqJ0YMqz1C8H05E1HA72sj85WqQFd+pui4PSasPkCx4UuFdgbEFv2E2EPZdkmpzOmPJ854xNN6l3BeSAa+KbgXCiWMJG8Y6w/GsQawHyX0lz6Z0Ba85cvowxuTXOV5EoP6M54fnNvLZVQ3mW9bl09nkptpM6CeeF5A+yBFpm/wnG85aWK6KBQ4z9YbvatkfkA/msPQoE0oJ5HPTr9U8o+0z0g3CP+WU38YVs1yPIyeqNaM4JxZMoaD6dU6+oBW42iASYCKvJ3LN21wa6Z5UAqkEUgmkEkglkEoglcAJJJASFqmKpBLI3wkEAAAgAElEQVRIJZBK4MmXAACEsQrkhRIwwMT85n+AFcI8Ed4A62BengEnCGmCZSCAAJb7vHgDvABoQnYAbpiAKbAVZxKYf7Kk1m5hDmiLxSuymmjJAitJrGWxYgS8ARyA8CGEFjKCMEA2JhTT42FyaAgT7FUhJUxIEWPNy/gA1NI+jqVCYkA4AXBRGSvaBqeSyPppMn5Plt6c0n3fOPZhpad1hqcae17+UO3i54issPNOdXY8e+ThicKDt5+bv29GZMaDnu0bPTul629yMAMNIHpN536Ufijypdu28b5hU61uO/U5Jydr7bih/dNKyn1xj65C9BjFxE+CQCnRdk0Hs74YsArAirljPCz4jJ91zohz/vCHs1HsDy/4tz9L4fS3DWXAitdKoCD3IitOqp/ynGhiOR66g/L4UGz+cFkuXrGQWlnzS60VFopEwCbHxHGChm6qYhHN3MGbgnmRWHVDCAm0ZG5kRdcyh87TxS4Q/HaucHr61LVxAuBJLBzGq1bNrum8ivJ1CybMvueJBe7IcSAQ1HjGdA9aZUcX54Kl11xx9P9Uts3Yl/l2djjM9Ixbfn1nPTN4Z972+3pKB7/L8WuDRaUzgaTwlPQgWdqTVDgJGp4QFJXeglXqK1gPXLDHWh7amMu8XszdvzzU+4litfFQbzbzLbdUjnSZEIce1Z/WYP8vXQ4i1XitcflL7Tj4wfGFP7h1evQ3C5FTZJ4o/M1mBuxJkxibb6myzjFGPLs2K1yICsl8jirehL+kehFJtZXox3pe9YEkZ8VthfOkU8ejI+E5kCs5hby2vUjDzD0WJG/uk+RuUQXUZv2HAON5yrMS4PpHVV+qanJGdbYNHSQJPZ+QFTyHee6ejBec47qO5bh2TX5KsZDnph7EuMkMylkm1KiVRFj0kJ5EFvN1bctqnS9qCGUU72SzWafPD+JSMwqHc1n31nozroq46PrManla8EwhVNUfq/5iNyEfzYxZ1/deYr24crdIi1XFj1vDr0myTl4L5guzL4I6ZO4kq4P1X/QXo4h3qTL3ANqRcVfwu+VdgaxZQEgyT5gtnr/dCuTPd6iiIzy/T/aZbMgKxhEvB8LooTMQHy/vuJHJecXmT6pCuqAHeFEkhJohK8x5kmflz299A94ld4euAwGyTslX+4uvbmY9wkJZ+fqm6TYgRD7TahdeORieHFRlneekrciDZK0QiYVj1YjIixHHjoczntvjSu81UdEV8pfU1QE86/JqIWFEAyXfnlOeFAtvC+3bsVIJj/h+1BwbVqqUlLDoUI3031QCqQRSCaQSSCWQSuBslUBKWJytI5O2K5VAKoFnkgSMxbMJGULfjdWz0mHKIniNlDAgo8lpAQBjQkjxHUCAY3gZh6zgRTwJ9fI0BLsB/wFOAFGIFw3wBIABSEKfAf8BCAAlAL8APQ+qQmYYUOTk0NfT00TaB1BmvCz4DmpIm89XxdoY8ALwCzCHUECMGTpA+2g3HjIGvHHaclysa1Ga4+L0BmizswDbKuEtOXlVjFSj3gHBPjWREzVPAToEDO8f9uZWloKxmX5vCXCQcWqerndFR1goQFD0dx361fKyWBmM/QN7ohr6gI54x5y8fcDtwXOixL5lN/MSoZ5ChGNIiuSwBMdWegqBWSIQkjUF+NHMBciWw7L2buzfO5zZv3cEsuDVytN88Uj2yisUgqYdqLaa0bJQ1LUEB81oZdZzeuYdy0NH2UjbWXf4/0ZZ+t/kxPWhvsq1F/dWv/KajH/0+1dFVhzKjlgLXr+s4XepQRt/gqovX9D5N6vlyHVRoX2WX7N6s7/bn7ffcW2yvjHX92qmYw1Pzp5zkjwWXQZT1uFWJJoyCXPjW9vlifGqeNb6Xwp3c41Es09x+ckVwjqB58bJgM+PWdGwhP/kZ15cWh3oubvcW3i3iIVf6LxoX2n13J764T1DyysNO3JHZHP/HOV136eIQJdGtoe1dUJEZQIxLwKbJbPEs8JuhYKqFfPW1I4Ra35swJreMbIgsqIrEK9wNsEj5+6sFKr1rxzdMzb/6s/fyMWU0leEkJ2QRYC13RIH/8Tw6t+JjBo+tNT3g99uZnbfH9tZ48zTTUase5BSjB+5AjYL2mUs8lmXWT/JCQAAexEXJcQZYYwUUswaCVetgnKPl+31CTdEWvx2qwGsq3+uio6bfCiQH+TdINcDIPrLVXl+bFUAtP9ZFfj+q6oQFjxzT4n8l1U87k1ZUXaWwkOFittTJcyPyAemq9RAGUlCW3M7yunIIVwhdYuMwv9sE+iMJ+C8RnlMc7WqgF/GG2pDu1ukBR4Kf6PKc++7VdfNY046ItLi5sL58Usqd9tD8s5pLw5+iSq2ZkYk/4jooFrCE9W3vk9txVPi51WvU4W0oC3MfRNSDlLOjCPPWsYO0J551q3wWwavA9YlPBqMh9W6YyH7NP/bCzpiBh+9IufIhCo5JLoVPD0otNV4OfCdZy5l3XhqbUiIs6/f9cjq4kj/fUvDff9cLeaR5fFS7cnna4W1kGSErFOYqM770jfyUzCPvqIKSUGeimTN6bxn58kPHlqwBvvyjgitSPqjNVtedI5TU3IbEl7R9m1a3/Na36fU+obuPqRG9/pRLH7McZvNJo+BaqGYkYNWJBLMVqgo+WGkJZVAKoFUAqkEUgmkEkgl8BSRQEpYPEUGKm1mKoFUAk9rCZiQUFgP8+LP2gzMZjwkeLk1iSSNZaDxygCkB6w3SSY5FmDSWFPLKHVL69enomATwFYVzwngFUAOrDQhAXghh9zhOzIAVAYs41gsOI0sjZXvVkDb6cjGCJv20Q5AI+MxA4ADwmGIJIA8ADTCqjC+xMtmXAGlAeoAN+gXesB5XMcAHSnwcDqjc3LnZBf8bRf7cfZq5akYrkfFFVfZTf04o9wQUXiX/dyjw5nZh0RkPHhRz+0nnWR7s1tDWqATypsBCEXFA2hdkcIPPOIWn5WLo6Xvbc6gA+E9Xl/PYScvENTekY/DK3JWdOl2xfW3hWj1aBlxpEoiMspRbDddKwIkQ+c5F0KMObOkteHI9tHe7N4dg78oX55fEYaa5Om2hKPiTbGW51eTyL/fmve/JRmUBJY1FTdoNqucFu/eV3zT54YzV7BWGc+BRLefvXckVpgge3j+t26v2plDBwrnfEVg8i/em9u7m3wD3UomDpqX1Q9+/OHs+K0C4YfPbUz5L6jeNySQGt1nDlyt+npVAFCAUKypNxY5cAS3yAjfZKkBqiS8TcN6MVyO/iMJwtdV/1SVOXZYAOX8mSYtDOiJNFWRKv0oWJ/5Rraez44qJ8eD37j6sr8WGPrDCttUF2oNSA/R8IJKr7fXi8r/pPj4UAj74oTcUfIBIcexm8HbSgCpcPiEmIKwwPtAqKXCQEFWTO0aqa/298xP7RzpCsgLXH2vEnJ/S6TFl3S/WQHCQVvIHcBjyFSSLv+U6vd1CtmOatvyjbudYvbW+9S2y4r1W5AnAHa3AokFaUK+EtZE8oesK7o3HWStxDqeMWLdPk/137cfCDmjpNpWT1S39jWnZ+/M79ssvTqW/S9ThWBgfUX2yJdwZj+piofbicoHdABhoHjGQHJQebae7NqbeACIbOiVt0QkpgmXClsOF3jNKat63BR5UZIFPTktePY3Nf80sLZvh7Yfh1FBW22F9KlqLtY1yMpR4yj/cpTM/87Gt7xJ2MxcxMjhb1WR/a936+jB7PicgscdenHlnnAwLL/weE6L1hOMsFAufgtqWcSKtBYiqk93xiMF15XPqwLGs6488vX3X1R+8II9GSHrxkNwQtshBzh2LfHIxkLeDUKEGaL+ROGKaB3jyG8eCFbuwfhCXm7wTGu7Hb+b8Nzimcs1WANZt8LO/DWat4wbfRh/0TfuPmdqx3CmkcsWv/LKK5uNXMYQH8ml777sXKt/tWINrFSsQlVrb8sbUrv+oXUP7sNcQoLczxiidBVGx0a71giSsJWsyvpYEd8wb9vOoDwtUAxFhoq3aSmAwUTPuH2UeOAo07YEOixdC4s5LygO5IZcW0mZskrlnpZUAqkEUgmkEkglkEoglcBTRAIpYfEUGai0makEUgk89SWwCXGQpFFQ70zoJhO+wngJmLAVvCgT/xtAE0AbQAfLUUN2mJBCCCoJJdSqT33Bre+BAfvpOzIAiAAEAPgHFMOaFFAMgBPSAtkCPkBaIEvkBHgFwQMwZ4ifMyEnQ37QNqzYaRdgDu2ZaP2P5S8AC23FqwLzVgNmAi7SfvoEGMP/AKoPq6IPidW5KuN7pomWM9H/p8U1KmHf8GIw9pyZ5q7zZKw6XnQrOaU8zfS4ZUekxdGcU7tlLDN1IIgzjdP1rNhEUOiN0Y8NIY58y3mDSIpDzw+WjzygqCD3uz0DSsK9U24fb3LizPf3CaeKFUumLHB7QN+Ho2Z5IPZnpShcC+AM8BIdQu+niX+OZffQQGGvQFCRFeolQLiuIUteYavBN2eaX56cD278wUo4aUVCKw2BoeUFluXf3Vn6H1jMA8TV8R5o79dXFn/Mu374NeQgGJU3xXeINGk2bKbixtIXVq3RcDU70Zz+o0tqB98mlvXocFDeKYKIucJcwuIf625AScBPE06q82JN5bf4fdVnC9Z8AytkEtLmUXtm4zHAdbgmgDbr6u0CKo1suoJ6IjS2LC2CgvXE5CFivQEgNd5V3Bug/KCIiO295dpzt08v9oqwwMQ+IStMUb6OsbHZ5f07j80/7AVMdw1hYnSPy4xIC9ueEkmxLGN71rJtftb74sz24fvlKXHO5K7RSxWmJq/r4snVrdwui/BS5Fhf1X1Za7p5l7B+kgTZhLVbl7fEEWmVCSZHi7Vvvcl3t903UP7nGZEOH9HxJLruvB4dAGA2JDHPsKS0EmvDYEEKEJaJdfl2VZI0/0y3xhMaaru//I+DYeXaKW9kaN7r/50ux9H+16ripdGd2NpEOK3NhMICZIYcw0tjXvq9VSirbldLSDwByMtBEPZarrskY/lRTYFJzbOc4GVYwaas5QfFAvaKjppXavuqsGhPSWgU58upKofFIR0zr2TLC8rcPVeuNPxGI2j+xluet5VHEPpLW5EjtB3t/1BnAxU6a9sj2fFtvu0eEGlhDSs/CKG22vNacI4r/z9boycPpTVvixURh2u0AiQBHgTXKmTSwd5S7SbN21zGD2yRYcgf0uhXVLt56XD+X6riVYE+MMe7khV4V7QKv5GMlxVUCoVn6G909q3jf+b5H6qSuwIPLYi15H6GrNDcZd5SuQfE2YWqr3ODcGLb7HKPvCteuW1m0Tqytz16nS40PmTd8twL4svvOGDvOjpvidiGuPuY6kFV9J5nN0YH/BagnAphECtJtpZiG7mEmv4rcpzol6fRrjCyt8VR5KjBea3h4yK/wmSZUDQ4HdcU7xVlXLtPeVB8Je6u+n5QUdqbYHahcrLhtk4g0nR3KoFUAqkEUgmkEkglkErg8ZdASlg8/jJO75BKIJVAKoETScBYJwNC852Xfb6beMMA8+ZFN7HEVDWEBUCXsXA25MVaPJinb6F/JoEk/QdcMF4UgIS84EMSANoASAKG8aIOeEiySwASY21+JuVkLKkN8ALJZCx7GSPAL9pBlHBANMYSQAkgGYtxQkPRbsAU2gVwwjGkE+bagGiMfWIZ2qr6SMuZlICsmPPz/vaVUjhwdHfukUIYT/cfqF2YjEXG9q8vONUDeac+e0Hx22dSd+gCYwxoDrgFUYVHzvGinZcLxez/bHY7epVZtb2LtEhcKXDq+8lhUNJyQYOUx8IKIvuecatxvRJyjxfiiGsCvuJlwZqi3N0JaDor/LsoW9wxsHCFHUkgu0Yj/CWBYIu65mI5mDq06h/4tEyHAeE6C0l0Cc0E6Pg1WXiXWyFpzNw8X14VLxcwClg9G1ju93Qbp6K8Qvb6c1a/SIt85I8MhJVPi9yAmCP2+2Wtc76kT87fCnyelQT/2B5UyoALrY+GD1o3KhzU724RJZ64/Kb8ib58VhUvJ+Ys87Sd6ogFanaCjYZoNrH0OQ8iElAUgghw9XmqrDuQp5CRhLFZVpLeh3rKtV17D888S14QyyuDvYmbjSkLowOevC9e8h1fvDk3tLi64IbRiMgKwhNNiLCY13ATIKfQzGW+vDDSf8+hfTuG50cH9shr44WKq79HhIbJm9MpctZDwlDRPtaTJDdI50Gt/+k/FvKAzsinzUpeoY2iqkiL6YIXznl23GCNYp2dEwlhvPySkHt3xP648gOjs1qz4hURHcstjwrWMORBOB/0CHKKcyEZyNPUtQiw/Q154zTEr91ec+RgtHY8ADbeGaaYpB2QUaZsmuekdQB6TGUcQcnxUkiSMaueDtBr9EPYctwTO/GK5tXDyi0wJE5Rs420FdE+kYWeCImq6znHlEC5HETRbowblH2b3ARxU6B1oZCpeZ5bymW9+o6xjflIuggKuTDfWRIYBwB7SLp1xBPnKafF/tsL+2/a25yd2B4sjw2FpbpM9fN4s5jiyI8Fs4oYeotGmeCFkfU66doxhUay64Xs0PDiqh+67tHJXSPPESn2W13axSbaBMmAxyNkCt5e/jvmuuuhQkExv5AlOsT84hnPNjxoNtWT1r3x0MELhzHlGo+o1gyp1iIZecaa+cc9CB1G5/EEekumGezyMoF1+R0PW8MLpSQnTK24FgqKMr9tsF7qLx6t9OaXRNo8IO8l5ha6w7M9MTAR2XkqRMXxa3OudGdeHjoQH4QQ61Uv5MphrSgnChnal8hr4fuxq1zcUwoF1Svd8aVH8zpWfJd7rFprzpYqzWV58vjKU2TL8826ck//6banvW3p91QCqQRSCaQSSCWQSiCVwOMqgZSweFzFm148lUAqgVQCJy0B4zlgQjkBdrWCmSTAAxABoCkF8HEtFeaj4aP4bkJF8El5Or6UmnANIAaAUcjEAF8GRYAQYB8EAQAFYBbHAUQAIAAmcExik4iHyxnM8WFkbmJs84nVMPcFtARIZOwAMyAnAKUBxAASDeGERSZjCMBJu2knoIoJCQXAAwhtEr8+HcdZ3Xvii8Iy2beUPl55qHrJUDPOXiXioqjE2lPypvhSOex/qW1FCwfr50/tyB4JzrB3heksuox+EP8ccM7MefYTJmzPjJObUWygfhEVO4TAvZLBV4CQJElFKCQ0kAW6Z0cHD7jF2WeFlYODlr+iXbM6DMAOolMGuZbyuEZzst6t+0F0WEDq1zKefY3mwoHlUv0zQ32FTDbrTezNvDZYLN3wgBJuExrnh7qMyDu1DWIBPf60SAuub+YlYdheqrYB4BPOaUPZ05yzhsNSkpNgV3PeGhAILrKC47jGW9tO2CykTPs136QezugCQ4IzH5Il+Le0MkD8/LAq1uBblZ/VTgDz96myXjA/TdR85puJO29AaLPmsE4zj7H0Zh/kDJX7MoYcB+jPukVIJAgX+vYieVnsGJ9cGNz38FT8yLk7GiItHkVBdYA8JHL3XnzOSyYemSqNTy3eLMv1g9rM2uVoxToigPihb77k0iOyZr9IOTGqCu9UU8iaV5ygn3+g/eTuoK0nyr2CaqGLeNH8nCpjbQDiaSeqzPnenr5c84DG3v5pNUsDF92nY5AJQDTeQl5P7YahSuGFkmFUc6PV6bGl90IyIzOIV0ha9ASPmReeoO3sfi/tFmnxoPTkAMnmVd8jHWOu/KDq929xDU0buk3vW0sm/69tuhOyS/88IuN0SDJAZyoh304UpmirZjPurN9cazmXc4uBH11azGZ7Fb1noFEXWG9bFQHLo0qw7WpikvKcMEBKomz7rmuXC7a8ujxvur+YqRSyLiGhTna9ZyLxnEBnCLsE+bKBsKDxD+R2P+9Qdvtdryrd9q2eqHaeQkVdiKcF3izMxyTU0ZhIlDH5WIlejx5S65dlzh+6enh5/1GAPV4/pR2TCzcc3De+KLKi21ph5ERbmBs886BAzO8Vs781SMnI8Pw0ZALeSegIhAVhvbYiL7kW5BN9pkLOrYioSIinVtgn3oGpjBHXJPQZY89vAwi4pA/0vVBrWoNLJWt5sHcdWcF+kTWFA/t33ZZtBnfa8cIDxUr9ThGM9O+xEBVcmnFOiFORyqtao+0wkF+U68yoSUloy2YQNPTbRbGhoh06WmrkKMyf1RMGoTwynIYu0CjksyI27GxfTy47MlA0+Ua4flpSCaQSSCWQSiCVQCqBVAJntQRSwuKsHp60cakEUgk8EyTQChUFVsFLKC/PBpAwL9PGUt+QEojFWNgDSvBSa6y91/DLp2cBwKBvxssAsAPQay02/FoBoAEoA8ACpIDoAbCALECOgB5YKyIvYwl+Ji3l22VvAD8ICcZ2ryqeIISomFAFuIPMAERqxX1J2olV9kFVwEKsPAGDaTf6AOEBGAIZwzWJXc3n0zFXibr1hBf3Xxff2NPjlnqydmOmZA1mq2GPvCy8c8PYLTej3FHltKh88CW/9lhAzK06xVgCEJOrgRA57YUQYf9OdV4pltH5C6Vgx0E7wt9TqrZSYdveDRkrvkXHzQnxQ7dM7HS8d9AjdHOFeOcCwxRK3/5DT8mdtW3/+EjvuQK+vqbvu11rtDGSvWphtvHNvxFE+QOtczvb/73agA7jcUHYFTMHAO4BkbuWK2sPLe/wFwchLHrDWpJQuUVWnOqg/71OgJCBZDigi+SUi7mpFZK1gfnD/Ifw+44TXPjV2k+lALzjjQUBAIEIyMp6gbxZL7gm4B/eXaw9eEgxX6kQHIwVoXAgnMjFADjL/MfaGwJnBwlzcw1/aXx6sSLSoSzCAuB+Xbnr8nMteVvc/twb7/1g32r1ULHaGFHYr+jh/Tsn77lkIq9zsr7n7opc90Jh75AmnYWxZ7yVfjwB+7+pyvicSjgz+gnJQYgm7vEW+utE5T1utDjYzOy0fA/nhvgX9Qc5cb/XqL5bdXGw9KkLG9nzsc+vZf3DpYHyP0EeIR/GBvKGcH4nQ1Z8UsfhAfNV1SmFL6r+xJVfCEWSfUX/s27igYJnDvKFnN65RlDYCyIh5KFynJxg25oYbI1zbF8vVFpzToneFaVJn9+y7JBnR+WxkBWEbXrXR29CdkleIjENA6uluOJ5CudV97OaY0RvEx9qnSsOIqfwPw3HdWfk+aS4THa/IrMtyfViUiTHvKb0klwySoV8xn/dVbu6Pq9M6KS2XBa67fGk2MiG5yX6h8fMhqJwbZde23dV30X1w19XTotnibRIPGTk8aRwUasJKSrHECuzLbCyo4EV3Wtbiz0DVsPPWCWl2xDB1qdwZN+pZPLdLm+2QZgxr76simchxG+yT54Uhgw0HhVsZix59kHeQyKQU4Wx3qqgA9ep0meelfS72vxbK2qFfqKB6B3XgVzDAATiDMKCMFbtXjnJfUioTY4KkYZ8RvKwoI3Hy7E9Yz+oJNzzOybnv3neg0enz/2t+U4S5gRN3rhb+hNLf8zvlJJ05JCICjuMwz7pyHb9TwZtRX2y6lq/VxwpS8ZzlPokcpTfoo63Tsb1ZuSZgzfdXLXqN/qKYZx6V5zyUKQnpBJIJZBKIJVAKoFUAk+SBFLC4kkSfHrbVAKpBFIJdJEAQJIBIxIQmnfl1icAKeAH203ehfYQUCRifboSFUZU9M9YXQI0ENYJAA0LTMB/9vFcA+DnWIAJPiEFAA4BSEw4Jr5jNW1iS59JhaQdjA3jRfwOrDeNtwRgCOCmsUKnD7SNc0zIHoAU2kef2MY+ABXARwBn+gQRw3fjkZNkcm3tW9eXp2HS9TM5Vp3XKggTKshq+6BtR3OlYOAqTavhPm+lUguLX6nGvXcGYeZ4DP7HoSHoDWQUsdABFzst5iEsHmmN+y913h/SQsryIeWw+FBvHFQ8xQ9SaBdjsWzIPk47HlLs0ORydOmztgPu/bPqdwpIBdwHeC8JouzZk/+uxVo4fXA1OPA/tG3DPVttgJx4gyrgPnMMUHoDAG/aK/mWm3bmH5Q1g/AzAp+Dn1I7mSMnWyAjmB/IAnIBEnJJFtShwg3VnB9es04WQIl1OYClrOeTmP4Qfj9+EjeBiEAepnAec5GwOsxXPCg+1NrJHKdC+ECKQjgBwrNGTaiaADrMYcBXAFXm7bJi3k9tm1nasTLQ48s6/UGFh8KLZl3Rtmu++NrnH1QYKZJwz2mVn5dHxasFS+LtQP9IaryZtTljzzrxm61j+U7ZQLhJdluVpuQK6QFRgyxe60Ylq1i/TWBuXbUkLVOG6LgJKWPyiyiHhn1Qy9W9brS0y4lqU4OlTw5n/GP/ScesS1685Z3X7vkBVcbvOlXk2U7S8x3CirX8/+ie36XGaHzsahzLttyKIIl3rpES8b/pO1b0hJH6G/1/Y+QPLNhOs2DFmWJY2z4nvqAZR9ngF176e2eClGQ+MwbMqW0Ck5X22JWFfKRt7o68ElP4TlSUI4M8Lizm6mom4zaUM7lRzGfwfJqRP81iRoSWHHDqg/2FE4amasv50C7WVREZrFt/pUp+EEPMrRO9cs2cc0fh3ESXlNy8ORqsZiEUS04h6cS4v2hVnLzli2k5dtmIdaQ4ZnnKmMD+5R4es92L5vhS/2r17fVcZkDeF4vyxvCffduD4Yu8ex0RFRTzzOS3DfOLtYP1j3ZCPvEs57fPVmQF+oGOfkLa7cdVayq4UbrTtKrytuJ85iPjwRzEoAEdRFchpzASMAQxc5v1jOPXGqdHK6SFSMNIc5bcLqwD64oIm59aGex56P6LznnoT9/orHbm9Ok8/iT/Zx1LvO70eC9rJZ+Xbj+oTvBjL6tVzhEhMSZCa5EURMpvonU7Xs4oN40UZTWbccrKX4GBhzXUXwhLFZwu0pJKIJVAKoFUAqkEUgmkEnhqSCAlLJ4a45S2MpVAKoFnjgQMacHLeRKyqPXCagAaXrjNMQm58QwEpAEaQEeoJpE2QBwgIWAaXhaAXMjMgB8GOAJY5HwsfLF6fjwICxt5YfMAACAASURBVDM+3J/vgKsAwADRWIli9UmhDbSTNjLeACe0CWCJNtIfQBQsQNlPXwm1AgDLtem/saA2XhxnAmRrNe8Z+SFvCndsNRgczjoNr+iWlSjXmapHhU8oJBRAKQTT4y1jAKZ7Vblft/JrW4zMAXlVFA65hZFtkbvw+uYsupSYmasCBtL248QoVrxc6/VHViEasFRHzwjf9AVV9HR/j7vn/Mv6fr50x+of/mM5PAQoiCXyZp4T//kktIZ+vedAbscXRVw4O/35ETWOsFLfrQpYyHwBQNwsDwPtBICfUMUiGnIHryqIAMsk0uW7YsdDWuDx8CXVO1UBP/HEeLvqurwRJ2g39+ssgJ20l1BPtBn5YhFOsufOAkhsQj4Z0PVBoY53KZDTvymMzP09lRpEz4e6taORzxKLf0KW3egFlXu+rlW3avq/aiceXayJtA9ZEObodIBLdIPzIWQ+bcXBG3xv3CoVXx4VGt9WmKoshAXyNQXC4nwvXHi1F8xqn39pb/Xrr1LC7nXW6Vs03iSO/msdw7podMOQ+STt1mgmfQn+bOyNtG05avY/HAc9eQXKyVtOs9fyKr5tB4wPADSyv1kVYJswTStOdrkU1UdrwcrFq/7SFbHtVaKoNm6966NvtM382ErAJ7HPhGZi3VbC5LgSxvahQLSEQiotFXLuimj2YRGlExLMqDqzIG+nQ8pXcZ8Ijpl8LlMmp4yIRDN3T+KWGw/RmDdFWvCMwdOG5+Wbt7qQCMXsZGbEou5WjhnlurC2B0tWWeQEpMXxsi6QWfcrXnzPwRmtOhfuOjoXZ4PA6VupjA8PlkdES4ha0DNMwLtIG3iQnGRBCDfIPfS1PcQXhOFm5d2iIu7XKjca160D0WFrNbrfGhdpAYHGcxeCgST0zB0ILOg5SAzWOnSi3WuFXCydhFpThOEvKyzU9j2HZwtTO0e95aFe5uC6IjKGe+BuNAtBdJrz7Pg1W14WhrQoySMu6zgiY+JYnpWWvsuXzI4d5R+ytQ9XOTlbOU0RXEHBs2ddxz2Sy9okeklCk/3QNeeeSW/SrdQn3ZdKIJVAKoFUAqkEUgmkEnjMEkgJi8cswvQCqQRSCaQSOOMSMC+oxjKaGxjw+3SApjPewCfxgsZKHPACAB8gC8ABjwWsrPFewEoZMALAC8txQlAATuK1wLEAX8ZTwYC4Z7pLAAOQFCYngbGMhaAwYWMAEQgXA0ACoEasewBYns2Aa1iBEmaHZMCcR9x3CA/6DWgLVATIiZ6AIHFPQ2id6f487a+n/BXGW6UgY9UFhX8CYGz6cfZikRiMEQAnwG+sY636958K3n1K4kPHAdbQ7VMp6DReEISCenjKydUM4KrQIgnxuQUAi55CENApgDhCQkFa4DXwNs/uGbqy/zc/fWf5PR9Z9u+FcHiVKvpJgRRpQzC3bPIfae+1AmfvrtvZlQW3n3wMsoKP0X1C/jBX0W8s4JkHAI4Tqug+9/gnVUBXPCvoLwQeRARzfQ3Abit4DbQS3kJcMIcgNyAssMhnvCGHWC8gGTZ4N6y/2ob/sNQ3ScE3hJHpOLoT1mW+o19fULz78vbpxfCeS/dNy4PivzSzmb/Y5L6Arhssu7doI9ehvxCbkJ6se6dLViREkOTLOoa8/8iy3Y8ocfTPOnHlRU7MkpaU9mdWEkbIjhVCyD9iNbMTeGFI5ps+wiAi8ERgHf89VcYXfSR0FKAzMoOY7XoBLNpbel7xBu6rZobusJ38jPIQJwbmWMzTdpMzAXIjITrY6eTn/eaDV3OgF/t9bDekymMiJ1thoSA+QrWNeTOtEGy2EiHnZQUvHYyLTdcqu7bdUw8iJS+Ph2SAMNnfk1+o1JqTmhfH5HGB95yvHARJW0ma3K0o1E/X7R0bGSjCtqEL71eFeHy5Ks+hTQtkBWXG24xD7H7qxbOHrL5K1RpYLF84PLny273l2j2eFT3sbI93OBNWUXB7XgENq3pK3iOJXyyKAu8O5mK3xbVbB1l7btEoHoxmrAPxjHU4OmrtEWnRoyfh92gfz9FPqOJVwXXRMXLVdHaknUTrJCv+Hx0faWymi9W6t+vY/KGl4X70FA8snsftBSIUHUVvHhBpgafFSf1mk35sJn+e6egm86EpYoIQUA8oV8U2VVsEWKSJ1adQYysiLMra72tTWVksFpp+NOsF9rLynpTyWS8lK7ZS8nRfKoFUAqkEUgmkEkglcNZJICUszrohSRuUSiCVwDNVAl08JdpfdB8TcPI0kimAmCEtDOkAuGkADsA5gCGAZUAKrKABENiGpTHIC14WADfrwLUzLCMzdgANAAUArlhf88lYmlBRAK+0me2AKYSzglhJYqirTqhCwvA/gCpgC0A2oBMgrYn3zSeV57oht85wl54Rl2Os0JcekRar8qxAlowH2xiPJ2Ie0gbuqfA2CSFFOKMTFfTsL1XxJMBbAt1IiBXKu/T9BASLCUUFyEefCcUCIEe4JXT5fMfO/M6lvT8X3b76O58rh4d/Vtt+RJVcBSdDVgCYY9kNcI9nEQD04lRmuDrwCkXuuTYJt8R8BgiEbOS+kAAHVT+qytwAVF3r0JqeA7qyPenrCUIaQVzQx5KIC/IgQGRCuDCeXBNQk1BReDI8EQVSBrkh24W+Us0fXlg9MLt9iHWKcXzbY2wEID+kE4TsV42sThY83ezeLdKCtfMOeVNM99Rv+t/NzMSNXjD/IrkmbMxDYbtWM7PHCrwxIb6KuiQvjC0IC+YXZBJ5NljLWBPx6CHsFfsoJwJ/E2+iYOXCSDUh6AQas431k2I87ZLrtMvjXR9NHJfQB2TGfpccAmfCy6JFpLCGoOO0oU85LRpRZC8FYewXi5nZrBIm1xr+BdmMq3B01kyzGZJ8u9KjPDOBqgiJxww4t8IUVSUT9B9PAHKOIBvGjrl8xso15Tuty51HrPJA3opEDxV2KT33Unix7cQXSxW+W6vMHfpkHhyTRJ4tn4ZTuX+g87+oURqMFq3bw7t0napVFFGxU9e6UttZH3hWQjTzzGdNe8EpdO4fW2P1OX2ig0lIxtB173vw/N2V6R3DhKziGUxOjc7yDm3guZ54M0nW/snMO+nZVs0jn4X5LRGJlBDPa9fUzyAK47pSoe/SljhyoorIiWXp1kGFFPNdz1mtVJvlbMYLHzy0cKK5cwriSQ9NJZBKIJVAKoFUAqkEUgk8/hJICYvHX8bpHVIJpBJIJZBK4MxJADAJkAOLWSphYAB3AbgAMAF4+Q4YCRGAhSXHA35CEkBsUAFGAQBOGBP8MTTdAAQATdwHMJI2YBVKmzCpxEIcIuWtqoRT4blMxcIea2r6iMU7AC7gCwCtAc0N0UEfkQvAE7IAwDUhxB5D85+Rp6I7yJJwXFe05MlY3NMatycK9GGcD6p+SBXd/dVNRgMwDfAR3fqyqiFVTolYIRGrLLcBtn9aFSt0yDX0itA5v6v6H1Xf4trZ371y4J2r95c/8PHZ5jchGdBt7kk4p27EBeTAx1XRVYg29BMwL/FeUQVQtv5M13nH3KfoA7IHEId0od8QHCaZNfMF0NfUdeCztp9UaXlc1ERccA/WAcYcoBxvBPrM/GQO0WcK7QT05pN5eyYKQDFzH4+qRcXHP3LRPQcbd1+2D7lAVLGu/cIWN8Lbx3i4cBi5GfBM+LaqITvpGzJD5tEmuQ1OuS8t0gL5HFzu/d7S/NBP9oVO7y0Tkz/6lZ7aTQDfEEtJPpJIueEDl3zXWcuNVpJcF5sUyDF0GYt11jpkA5FEn06KkGqRAowlczTxNMNqXbh54rHYBghvNYfZR0V2rMN4bWzlmXRC+bV5OTEnTTirJKSfrOOPhVGYqSrLgnIRLCm0jxu58azC/sg6PsyJsEieUY9DKB/mEM9LQHVIFGRPYnV0nrl/WoUE3UrYbY0rdNQuX7nO6aRynNh7FPMp8bdZJ3rWV8qW3h3rGhJp7sufIF62JiNptdRrJjpkLcaL1iu1vanLQ1KQ1wrPLJ6XFBOC7UR9IiwdHh7kqGDN4jsFlu1bqstKut04NJFcFm8t/LmYr6x9z++4OOfiEcIahjfXmXhuoD/mt0RdurEiskv5tW1NKnsytqJMEPKvtShPiznplu/Glq+8J/7UXOmMEG8nEmC6P5VAKoFUAqkEUgmkEkglcCYlkBIWZ1Ka6bVSCaQSSCWQSuDxlIBJzAmABQgHYAdAhfU2AAEWoybkEiADgBeADy/6WHUTEoLtgM+ArYasMF4bj6ntm+QSIRc29wepA9jlvpAWJs8G7YeUANigP4ZEAUTif6yM2ccxbONcAJ7XqwKiAMwArhnLdPoCQMK9DPj2mPr1DDqZ30RY96M3JiE7wB6gVE0eCmcCdDpZcSYga2vMP6BPgLjv7TgZkPdXVNGtl6oCQAJkA/CfTluZO8wlgET6z1xBT7/R+v4W7u9Y3p9f2PuTUWnl4Y/Xwhlkg7x+WZWk26B56CbhnQjfhMcQJAChngCi+TSkW2cb+Z85SWWOo+/tv1O7eQ6dTj/phvG4aIi4YM5AzNAXk1PGrDVGFqwtBsBMzt+k0Ea8XCZUAe07CQ4IHKy3P6xKvHvmN0TOzNjsciBSwReBg5zYD3HyG5vch7YawoJx/9+qEJ8kC0e+6AFgP2Nz2jLarJOtPCEiuf5/9s4DTIpia8MEySBXRUAEyWHJOeckgiCICigGUBEDBkTEhCKogKiggCTJgigSFBAkB8ksOecsUVFy/M87TvM3w+zubGTD1/epO7PdVdVVb9fM4PnqnNP3fJKrZ23T/JlTSa5eGGkhn8ZbrgqeGQmTk5pQ8eq1xCkqm6n6tF0/aqLFHjuPdw2CBIIR64W1zbqD2zgriEcINs56CM/4ne+8yHgj8LljDh5vDW8JzxhCwkYfPBtEOZ4LYhz3On/p8lWzhV/lu/+4/V6cPXLiNHmeL5tocS06dsZ7d/xfsbXGZ4zfEcRGQn3hzVLayx7PxYC9Ekqe3Z6o5LkdZi1P5xEpUprWYnv+bbJRgc4s9fsTnbKSPrF9okywyGVRyHKZ+X69vdYxigii4fHQ8H1GiBQIhDwPfl9Zf3wO+TzD6PK37Zq4J8L3I+Ig1zh8BQs80PhOYa3P4xn73jC8f3uFL0Q4R5Djt+k287Yg0fafiZNacpH/Htyl8xcvn7V/SXhynkSFh1B4x6r6IiACIiACIiACIhAVBCRYRAVF9SECIiACIhBTBBxDFP/RjrEfQwX/YY7Rj5BJD1jBEIaxlbANGL8IDYXBn9886mGU4TrGQgyjnvj30Xg4xmdugQEYMQHDFecxatawgmGT807eAnYqY0TiHOPEOIGxl/BQxN8mGSkGT4wizJ95YqjGaOF4cbhZReP04k3XjoAFP+cZYcRzkpzH9EQdgy1eQ12s9LbCM23iXQMYqXn+GD7xjoiMWMHcWGPdreDpgyDo/BsRLuy+Hm/lESomTpSkX5n0n83d8G/vNScvrXOMuhjiCZ3CWPZYQTjDsMc8eEVYwXDn14LpJ6STY+CNCe7cC+MjuTSc7wXmgTGdfB0cXIOLE7YNAzMh53hFiGBH9SArfJ8gMjJfzlEfcYFkv8ut8DmFA8/OERcwiCbq3c5zH9Ye10g2zTOlNPXWJdE2AtBwKzyX2lYIZ4V3CJ5jtMUjiO+ZiApXnkEEeJy9miT1zquJUqbbm+W7fQV2l2EN8Z3MOP79N03t90+la/i2eVlcs7BR60zcYB05nmaIQHiAEHYHhs53mLOTPMAh3FAtqkRa2DqhoRLjvREFhl/H0Myr83z4DYOZc5Bv4MLlK9fzEV33FAkjZFBEWDkhsUjGzXxZk45AybjmW8G7j/XP55pnyrM9nSTR1R0mQgWlvHppYzLLcJ766vk7Ul2zGFaJkp7PePlv6iZOZjo9XhU3HMzGnS0itFF7g3NdtW+/q3s8lNJ7TPM2wmuM5D/5sojPLRDvEPFDOwiXVtJbAWGC0E5jrdCW7zzWIoISPDz8vcXdpxNCj1H48yxj9NWt8J2ZiLBkgYSFCmPcnsuOcMF7W5eOx841y43CeD1Cq5M7JZD+VEcEREAEREAEREAEYisBCRax9cloXCIgAiIgAr4EHJECAy0GfkQHQlo4hkGMD5gy3LkpKtrf/Ef9fisYFwifg7EBjwT+A5/fwSS4QZiHRNRsBfUZtdfzgls4YZqc8Tn5JjBOYmTEOOqEIsEwhOGEsbP7mN3TnqSbVghxgdlnt7fAwUnq6xhQuIfTf7TMy/fhxIO/WReIXRileR4wxVgcopE9BubMs8PwvMEKhjGeNePByMmaZswYyKnjGNduGlaACcK5F/dh3gh/GJCPecNF8bnCwwIRwhO3PXGipJuKpHvzwb3nJs3Yc86TWBbvBGcnMeNjrbJ2eY/3QKxch94QUdfM04KD8bIGHLGP+bKTGsGB9wiCGGQRC9k9jScJbFgzObzv4YdAw2eU7yQ8HTi47hZh6A/Dpm/4LqcOwirfb3wHzLNS3dsf64D1CV8ETtaBYwAnHJQjVEQrb2/yZ8Zu90tS5Xzy/Ov/zPDOzszHP+N7ivEkOpDpS8JCsVM9SbLLhxdacm4EQHc4PtaGM96oEFijSrBgLMzN/VvifYyRenGPz3kPA+c+vuOP1mfozITcFmZUd0QjhBrWLs+Q3xiEO9Y7n29+l/bYcE9aeKe7LQLRHSZe3nc1cZL9x25LnzzFbZd2FLy4t37SRFc9CUFuOgIUKywXRaJr9knkF/OafQNf49Nkn4JrjrTj/5uOs4h5HHy28PLxPfh8fGeFz20pKyOtsD7ZBMDnls8yArXHO8HvHP7/JL+1jkcWYm1jV33WOZ9RRM4oWUMhJOV2RG33+kHIYCie8TvtokPwCoOPLouACIiACIiACIhApAhIsIgUPjUWAREQARGIQQLOTm4nTAOGLnbDY7Rjt24RKxjzMIixSxohg/9ox6CHcREPDOJbYwikLYZET+ik6BIr/LDBqIJBiDEyVgo7O3NYwRjEeDnHrnqMp4RMYawYX9i1TULaalboh3bMm4M+CXuFkRnjKYz4jU9qQkkim19kQqR4b5EgXuCE0R2Dl3PECLswRIWLlkAbwzUmP8QrPguOAOYxTAUoSoT1EJkrnxPWE++5zzVEC3u9YEZqQhS5E81OyZ6qcbHG+Z7CqE8yX9Yqh6cdb2KrUBECCObsft6OGOTkxuFzyzmET0fMghUH4oQjQPDq5FNwBAnMrtTFMByI9wPtMJ7yOWZN/mplnhVEE8ZAX5xH1HAMrFFlsA8Bj9/TrEuO9H/e9U6ie4p/dp3h6v3pGKfl17hW8myqUofNw8ITz9+8aa5aovXE3tBS4blXiHWjwAPC3bevsBAlY3R14rvOfI3aYRnLo3o8Tn/ucTm/JQjqeFtwzeN5cjWRZVNPlHj7xcRJkiW/dinFnVf+TZ7nwqEU6a+ePmVixUyrc8JWJJ+Vp61VimtnPZ+NDInT2+/c5UQXr/2V6HjiuxNlsfOJLAdFosQmF9DjVVsdeFFwXDMpAOHiupwX9sp2wivS3BErCEvHZxVPRoQ0flv5rOBlwXkEWj6XzJV/C4Qo+oYAnBHy74lPvf3iCcWB0MPnkt9nftcRRfjcR/gIKyl3hDtWQxEQAREQAREQARGIpQQkWMTSB6NhiYAIiIAI3ETAMVmwE5IdkRhPiLPNvkuMePymsSuUUFAYC9hNyY5LTzx1b30ME4Rpye69jrEiSnZAhuN5OcZFxsucCD9B2WMFowoCC2MnljghOTCKIFwwb+aFIEEfCDQ1ve1IlIpAM88KuzpJoorpx5OE+T8HkujxIAnHvGN1VR+Df4yIFOEEwlpxh8uJDqMm/RPPnXXD2kIM5DPjHKxT1h07iJ1jrQkZuUzU2O0SJ6JjbOHEFb7q5mkR0uHZxez1wMDo6ISQ47z7u+Oc11vjpn68eTIcg+V1MSfAEXq9GDyfZ74fMMw6972+EzyqkmoHOCZ3NXaSswM/hxWMwB6Ts60JxojIat9NppgmTnXcBIrr3iRRKVZEYMyBNOH3JUCfgLC7i+0GZz/rx/m9Zd26je1O6DxPqKPnSky/tmRJUJLcFw7xvPmd5bdnt63Q5Gb+X3PtUqILlnNi37V/E92Z5FKi+6+dst+j04kOJz5teXeSJyqVOFmio9eOJsp09UyivBbqKZV985yxaFKX7X/pb5AOw0bs1MAjBIFxpbcgLLKBAe80xohIwfcbv6f8e8Ej/Ib02b1+2yETPW9tzr4j4d8fiDqEleLfE7Dic8B3JSEc4ZHc2jlhIBFxA5+NaoqACIiACIiACIhAAiUgwSKBPnhNWwREQATiIAEnzBE7FjGEIVI4wgWGfHZ5Y3xAjGAnr+3s9SQNJX8Fhgl2QmJsJNY7Oz4dw4slOI1xgz7GIIQIQkpQECgwciCwID7gCUICXQyBnGPczJdktVg7MPyRT4D4+BQMyBjZSRKc2wrGEXJeYDxxQo7EOSOyjV2Hl4BLUInO58ga4rNCyDVyv/A5uy5YeMNDsU6rWFnoeji7zECdza7jFRQvD5eg4eYf0LPwMYb6b+M1iPqB57u33DeE1C3hbc8aUYJ78z3G95djFHa8bNhhz/cvu9rJ3YHQGpcOR5AK6BnHpYlF1VgdgbJChc2OwHvFPGf47fnHpB6LFmXCxLVEyRJnsffXEh2zEE87E6dNlNF+yJPZt0ywiReZrv5t+blP2to5n6iw/YKZw4b9v3llWH3n97mM9cdv+29W+E3MbwUh9Vkr5IXhdx1Bf5gVEogjSCA0IZ443kd4ODBGzjsi35kwRYrAQfGd+bsVfp/Jj8Fa5z2/xdwPsQSRRIcIiIAIiIAIiIAIiECABCRYBAhK1URABERABGIFAf7jHyMEBlUM+fOsEMIG4YKC4QIDvWMcw9uCsFEYNjAYsPOSHZcYoTCwYWhwQprE5ASd3fIY+zDsOSF4iJWP6MDYmCthq9jRznvEB4wuhLdgjggvGGAw7FAPoyEGEgzMznVnd+ytmGNM8tS9ooaAY5xlXRJGjc/aDYdXtFhsJ8kPQ8JnJyxZFzNgv27X8fTRkXAI8P2FcuHk23Bmjicb1/gu3mDrIq59B/FZiI2eVrF6ZXk9ZzzfIyZenEn8QKJr9uoJj5akvuf9PxYSKgm/eBb+abNn5Zwx0eKCRwDFsI/Axe87Ar0nj44VfrPxVCCUE9fpj3XF+kKkyGEFUQPvRO7NdScPiUfw8wqOkRb7QvCOIAcI/77g/qx7xsaGAcbNhgn997ZB0CECIiACIiACIiAC4SGgf0CFh5bqioAIiIAI3GoCeFlgpODgFSMYBn6ECbwq+BtD6yorGDbY5ciOX8I/sFscgwevjlCAUcSTFPgWTMwxDnNvjB1OolMMMwgWiCvEsGd8/M3OUcZLslDmw284u91ph5cF4SdIyI04s8l7HiawOOZNLC4D3C140HHslggOrJ8QPxNmfL5q4gSZXV+xgmjB0drKVjs/yK4TDkVHwiDAdykGWr6TnPwazByhmGt8h3mScMfBQ94VkXhoTtgvcpY43XjDgvkKB6ctbBq/006eKqrz+8530ADveX7nKHy3sK7GWHHCPDkeFE4ODue7K8aenzdxOWNb6h0n9+bfI4esyMsxEutITUVABERABERABBImAQkWCfO5a9YiIAIiEBcJOMYMx6vACRGFQQBxglBJGOsJV1PXCkYRDBt4YhBGCmMa3hgIGngjEGYpUokwwwPRckj4q46O4CR6xsDBuDDc8IqRA4MHuzZJqE38erwrKlvBo4L6e6wQ3qqxd+7Ml5BSiB4kSuUgrBS/98ftXmeVyyI8Ty3h1HWF+GGh4qnEa0kTIAh1cpXr7sP+vmzXptq5B610tVLCSg8rae38Z3bdCQ2UcCAmzJnyPcsueHbFu8Pe8Pz5DuM1rq4Fj8E7ihN6J8xVEvasfUUMxyPHeXV+QJ0QafzN+gp3iLawhxKxGt4QWZfN28LJfYJQ5xFrXPl9Ita5WomACIiACIiACIhAAiMQ04lGExheTVcEREAERCCqCJixna4cDwsM94gPjvdEDXuPYZUk1Q9YcXb27rb3nnAUVtg5jhGfnBHszMSIz3uMbJdutSGfPBreMRHqiRBRGAAZO6Guqlqp732/z3ueYBrkGWBuBa0gzLDrFAbMCwEHUYZdn7TBQ8Oz0/lWz5Ux6Ih9BLw5CfhcIPzhrYNQNs3KTYKFM3prw2cJkXCWa0Yd7X0/Ey2cBNWxb7IaUZQSIMk24cLo1JtwG9ELEYvv1wXOtSi9qToTAREQAREQAREQAREQARGIlwTkYREvH6smJQIiIALxkgAGfcKOYEgl1wPG/Pus4GGAQIFoQcJLdjRi8Kc+BjQSATtJqfGoICcE1wmXRNil2BQmiVAWGHkRZBzPEEQJ3pNolOsLrOSxUttKee/4nR2dhbxcSExaxwoiBQlv4cBvvnuXqv2pQwRuIuAkpSXMCp8TJx68X1RmiL5oBmriz79l5XNvpZ72es7Oj1BOi4SxwnwECdYN3zfE8D8YF8SKbqOJcHbT4fm+lIdFwljDmqUIiIAIiIAIiIAIiEDsIeAYOGLPiDQSERABERABEfBPwPFAILQTnhVOkk12eDsCxGx7j2fBWiuIGogbCBbkeHjMShMreGYQSoIwJvRzNZZ4HDihLRBViPtOqCvmzG/1Iit4kBS2wu71DlaqeTFxnblw4GmBmJHRSlkrTqJx+iT5J7kwkps3h37/vcD0chMB1iGfJ8QxQpOFuVYQLawesea/cvX2qb3/zEQLcsboSCAEvF46rB9C+SCyHvaei2sE5IUe156YxisCIiACIiACIiACIhBvCMjDIt48Sk1EBERABBIEAQQGdu2Sk4LfsDJW8CYg3BPCBAmmCbZPCCQMrhhSy1lB5CCJJ7ku2DlOUmHasJs8MeGYYpFowZjwssDghxCR3QrhoQjTQ7goPETcBx4UGIVJcuskJOc67WFFefrEmQAAIABJREFUQnJ4IeIQRgpvlNg0Z5/p6M9bRcCVx4LPGZ8vhL0wBQvGa21Pm2H6PXvL5+9Z73p82V7T2/kX7RXx7IYkuL55MW7VvHXfKCfAmuE7l+cdmzzYwjNRxp5Y3hXhQaa6IiACIiACIiACIiACIhA1BCRYRA1H9SICIiACIhBNBFy5K9jxys5dwkLlsIIBHy8KDGMY+TGU4lFBmCTCJhEGCrGC83hj4KEQZIVd49TH4wBj2plYIlY4BN1GXXJOsEsZ0YHkxszXfeCJgScFBwIMggxzgxO5KzA4420Bq7lWEDEcjnHVkOiDQH9GAwEMznw+SPTumww3xNuRaNvEiVe8bdp4K7a013usfOFdgwhmOuI3Ab5b+D7iWd8gUsXWaZsw4W9ocWLssZWpxiUCIiACIiACIiACIiACESUQ0K65iHaudiIgAiIgAiIQWQImJjhJojG0I044YZLwqBhlZYoVvCYIm7TfCt4JhE7CuM+ubmdnNwmE8UJA0CDXA8Z9DFKx7bfQ2ZWM2HDcCnk28I5AcOF1pYspYgwH+ThWe98vtdcfrfxlhbBRzBVuWbyFsFDufBau7vRWBDwEWHt467BOwmW0NdECI/XrVl51saxl77+3Qsgo8rPEts+cHnvUEXBC9yF0SZyKOq7qSQREQAREQAREQAREQAQSDAF5WCSYR62JioAIiECcJ4AhDJEBI31mK+zaxhCPBwFGePI3UAehgp3h260c8dbhXAUrGP/JeYGXhpOsO1EsCgnlPCQncTiGXUJbMR+EiobeeROyh3OEvCJMFGIN4Z6qWqlkBeEGgYZQUXDAw4T3tHF2PYfLEO0MTK8JggDrhCPcggWNvJ4Wg7xrt7+9brRCWLK23vKMvf5kBXFRR/wjwPcSggXfXTpEQAREQAREQAREQAREQAREIFwEtMMtXLhUWQREQARE4BYTINQRXhIYVDHqk9sB8YHfM4QIdoXjbUDuBkQNrmMUZcc4bRAwNnvfE24JgSO2JN32Rcv8COFEaJXUVhApyNERbIXwTog091lBqEB84Lpz4FVC0m5eCYFFLgzqwMcpnjwWvjfV3yLgJcC6wksn4JBQbnImWvCZIxE3wmJPK+5/cw63v2dZ+KisVhLH0aTMWij+CfA9g1DB8/ccylWipSICIiACIiACIiACIiACIhAeAjJUhIeW6oqACIiACMQ4AZ8cFhjuia2PsR5DKB4XhJjBcE9YKM4hUOyyQjJuElJjoC9pBYGCvzHeI3LwilHtvIWduuX5HLzz9OWLQMMud+Zb1DtPxt7ASh7v/BEqCB1F3g7yXOBxQZgsDIe0I3QWc2X+hJTa7b2GgHMpluXv8J2//o7jBBAkbAoIh1WsjLaCp4/7qGt/rLDCelRS7rj/vJkBz/z6s5RgEccfqoYvAiIgAiIgAiIgAiIgAjFMQCGhYhi4bicCIiACIhBhAk7uCoyfua0QDopd4AgUeBKQo4Gk24gPGPWpj4cCYaAII4XxnzBQGO4x4LPjm93jsTk0kiOkMA+8Q5hnESt4XfA3O5mzWylgZZaVhVYet4JAg4DDXDdYISQWfZGImzaw0CEC0U7AjNV8vk6bcDHDXsls/KWVh1w3JjcLeVe6W5nnXdu3XECMdjDx9AZecSI2f6fGU/KalgiIgAiIgAiIgAiIgAjEHwIKCRV/nqVmIgIiIAIJgQAiBCLFn95CbHxyNPCKJwHGea4hXLCTm2S/Na0QRooY+k5YJAQAvCtiTYx1b3JxEoy7ixNehZjwCC97rZBce6oVxAsnBBYbEAiBxd/MzRFv5tt7cl8gUBAiisKcZRA2CDpilABrDs8nBDW8LdxHeftjkhU8g8jDwudV/0aN0cejm4mACIiACIiACIiACIiACIhA7CAgD4vY8Rw0ChEQAREQgRAIYMC3wyImXXOM94RAIi/DHV6jJsZ48lfstIKYgVjBNZJLYwjldasVBAs8KkjSjVHfk/shDoREwtDrxINHuCAHB38XsoI4Qwgo5sg1jplWSLqNN8UO75w5hycK9RA1nOOG0C2u83orAtFFgHX4hxXClXW0QkgoPC84KlshP8s2K++aV8Y0e/XkZlFYoeh6HOpXBERABERABERABERABERABGIXAeWwiF3PQ6MRAREQAREIgYDpFey4piBQkMeC3BWIExyEiELQIEwShnrOExefPA94FBAaKasVvDE4SMxNvQsmWMQaLwt/U/fmtmDe5OtAmHE8K8jRwd+5rNxvZbEVQuvks0K4LOrjUUEYrH1WyHPBXNmsAENEm8txQLDxh0Xn4gEBEyRYo4QzI0xUDT9T+tTOTbCC8OYkl79eTSJGPFgEmoIIiIAIiIAIiIAIiIAIiIAI+BCQh4WWhAiIgAiIQFwhgCCBtwEFTwEM8AgUGN8xZmKAxziPFwVHTiuZrBAaijoY6/HMIH8FYgU7t+NKrHXGiVcFrxTHy6Sgd254lyDC7LFC8mKMv8wdRnhgkPOC9szb8aq4KrHCu1L0cqsI8DkmEXxjK495X0ko7xzv2hsKa7udFRLL814hzW7VE/PeN03adLdnyZY9x+VLly7t27Nz+5XLl2O18HuLcen2IiACIiACIiACIiACIiAC4SAgD4twwFJVERABERCBW0fA62ngJN7GswCvA0fEIBE3f5NsmwTb2awgXOBZQZiZE1bI/YDAQWgohItzcclgb/Nn7s7vNvNmHniWsPkAcQJBglBQTj6LIHs/x8uC/BeIORh7HZFG3hW3bjnrzj4EzNuCzy/hyvCcmmylcAiQnvReP2seFo44KZ4xRMB0ivSdun3R9/5GDze77bZknvByZ07/+8/YYQO+Gfhl9y6XTcGIoaHoNiIgAiIgAiIgAiIgAiIgAvGUgASLePpgNS0REAERiG8EXIIFU8NQ5uSkYGfvPVbwqCAUUmorhEDC0wDPihxWiJtPQm4EDMQOjPsIFnFmp7Zr/o6HBAbeu6w4Xhfk5uD9X1YQcBAsECiov9sKOS7g4NkJHZfmznh1xG8CJli4J8jnmFBneBD96Gfm4+zc71ZmW0F8vGLiRVzxloqzD9K+MxIPGDN5ZqHipcv279X1gxV/LJiTMnXqNHUaNH7kiWdfen3u71Mnd2jTsmmcnaAGLgIiIAIiIAIiIAIiIAIiECsIKCRUrHgMGoQIiIAIiECABK57B1h9wiIRA98pGO8JMUOOB+oRBgmBgr+5hucFbTgfV42b7nHzHgHCyUdB+CdECcQKwkAhXCDa4FnBnJ0jrs49wCWiavGAAJ/TTVYIdVbBSicrdawgRnI08xbe97Yy2QSPLfZ6Q7go5biI2pVQs17DJmUrV6/19kvPNPv91wnXhaT1wSuW7t6xbUvnnt8Mrt/ksSemTfzx+6i9s3oTAREQAREQAREQAREQARFISATkYZGQnrbmKgIiIAJxmIDXw8CZAb9fGOopeExQSLSN1wEJuREx/rSCWMF76mHAx6jv5ILAyyDOGO995g8HJzwWc+NIZ4X54EEBD94zf/525unxxohL847DS1ZDjyQBr9cF65z1nNVKGysdQ+gWYQ5h4zcrvD9vgkWc8aCKJKoYaf7F4O8n5C9UtHjDSkVz2/fRTd+dQyfMWJjSXC4er1+lVIwMSDcRAREQAREQAREQAREQARGIlwQw7OgQAREQAREQgbhGAGMZ8euJl85ubDwN2F1NrgoSS/MebwuMnfxNSCQEjOvx1eOB0d7J34EgQcGbAk8KRArmTMHjAqOtEzZKYkVcW+kJeLx4SBDqyQoiI94WH1ghb0tbK2t80Nxpfw+ystzKMis1TfBIb4W8NjqigEChYiXL7Niycb0/sYLuZ06Z+FO+oEJFU6RMRUgvHSIgAiIgAiIgAiIgAiIgAiIQIQIKCRUhbGokAiIgAiIQCwg4O3wxyGOwx6iJcIHB3gmT5AjzGO7jtNHeBBZ/yJ05JfJjRHQn6I5T3iSxYG1pCLGTAJ/jXVYGWxlmpZaV8lbqWSnrHTL5bCgzrSBgnDXRgvBF2614QsYp30XEHu4dd96V4YodIbWeOHbEkJVLFs27cP4cIrIOERABERABERABERABERABEYgQAYWEihA2NRIBERABEYgtBHySUTvDQqjAsOaETeK8x9MgHnhWxBb0GocI3FICJkTwOSdnyx1WHrTyqJXqIQxqqZ3fZ6WPlY1WCBmFyKkjQAIzV207dPjA/r1PPVSLvCI6REAEREAEREAEREAEREAERCBaCEiwiBas6lQEREAERCCmCbiEC7+3llAR009E9xOBmCPgFS/S2h0LWPnUCt4XHHhf+XoUEy4NAeMlK+S2wXMD74vrHks0VNLuG5/fgDGTZxYtVa5C5aAst1+1I+aeru4kAiIgAiIgAiIgAiIgAiKQkAgoh0VCetqaqwiIgAjEYwKETEKUCKnE46lraiIgAv95UP1jhRwWhIjKYiXIytNWxlpBpOCgzv+8dQgvhWCB5wX5McpZIRcGSb61qcdnVS1fvGBOqtSp0xQvXb6SFpwIiIAIiIAIiIAIiIAIiIAIRBcB/cdYdJFVvyIgAiIgAiIgAiIgAreMgNfrAu+K1FbYpPOQlSpWWoUwKMSLX60ctELi7s1W9lq5ZOUG7wvaJzQPjDz5Cxb+adbS9d8P6d+7V5dOb9yyB6sbi4AIiIAIiIAIiIAIiIAIxGsCEizi9ePV5ERABERABERABERABCDgFTAQL/CgyGelo5UmYdD5ya4jYhyxssPKYSvkvria0AQLOCFYpEmTLl39CoVyhGdVZciY+Z6rV69cOXn82NHwtFNdERABERABERABERABERCBhEdAIaES3jPXjEVABERABERABEQgwREwgQGR4bSVkzZ5PCiesJLbCsIFnhT+DhJ5d7Uyw0pPK09ZIfdFIxNAilnJaiW9lWReQSRec5028cfv78maLXvpClWqBzpRC9OXeOjP0xc0f6bNK4G2UT0REAEREAEREAEREAEREIGES0AeFgn32WvmIiACIiACIiACIpCgCZjIwL+F2cCTxkoGK6WsvGqlsgvMdnuf1w+oc3YOb4vjVuZYQdTYYIVE35w7a4XcGtdMJCGkVJw/7sqQMdP0FZv3z50+ZVLHF59+LJAJFS1VtsKISbMWd2jTsuns336ZEEgb1REBERABERABERABERABEUi4BIjrq0MEREAEREAEREAEREAEEhwBr5BwxYQLknFTdlv5xcrdVtJbSWmlvpWP/cBJZecoJPHOY6WNq84kbz+L6MP6J5QUOTI4EEmuxEUR48Txo0cQHWo90OhhwjwdP/on8wr1KF+lZh0qBC9fvDCsurouAiIgAiIgAiIgAiIgAiIgAvKw0BoQAREQAREQAREQAREQAR8CJjJwhn8rJ7OSxQq5LxAwCAtF7otcfqCdtnP7rdCYZN2ZrWS1csjKTiuEo9plZbEV6l60ggcHx3kreG1weDwzvCVWJfguVb5ytSE/TZvXv9cnnQf36UG4rFCPnt+O+LFQ8VJlGlQonDOsumnSprv9zOl/PeDDcyS97bbbLEXGlWt2hKed6oqACIiACIiACIiACIiACMQ+AhIsYt8z0YhEQAREQAREQAREQARiEQGveMGI+LdzUiuIF4SRutf7SgipFt73iA05vHVCmsX3duF2Vx3EDcSLmVYQMDDaI478beVfK4SYOuPqjDBTt4zQxHmrtqRMmSpVg4qFc161wz0QclZ0+LD7Vzly581/8eKFCyXKVKhsWsKV1V4Pi8tXLl/eumHd6mH9v+rhbvfgIy2e6tzzm8E1iua8G9Ei/f/uuLNt+3c/Kl6mfOUjhw8d6PNp57d379i62d0mT/6Chdt3/vSLshWr1jxtbd55uVWLJQvm/O7UYSwffzlg+LgRg/ptWLNqeUjA0qRNm+6MdRDZdrRPkjRp0rc+6tF7yfxZMxbMmj7F6ROvlAeaPPbEqqWL5o8dOuDrsB5efavbvFXbdrnyFij4z99/nZw/67df/5j7+2+L5vw+Lay2ui4CIiACIiACIiACIiACcZmAQkLF5aensYuACIiACIiACIiACEQ7AZc4wA5+clRQzpqQgZCAiLHUygArqAh4VWS0EmSlpJVMVg5aIT9GQW9bwkzdYeWKFYQKxAiECsInIYbss/KJFcSAP6yssYKHBl4ZhKA6bPdGzGA8p7ztET0Yi8fLIDoFjQljhg9u/8EnvSrVqPPAwtkzpnI/5zAdI3VQ0eKlzpoAgGCQ/o477zqwb8+ue7Lelz1ZsmTJ8YI4fuTITaGkChUtWTqpuUpcNVeJbDly5Rk0bsqcTPfcm3Xvrh3bqtau9+CaFUsWuQULEn9/M2L81L9OHD82Zui3feo2fLjZu5/1/rZhpaIkUvcchYuXKosQgmDhHqP7fbc+g0flzJOvwBMNqpWJbDvaFylRuhwJxjNnuTebI1g89tTzL73zyReeMSBcWGStwzOnTPzJ35gQPLp+NXAEggXixDfdP3ond/4ChejTHEmSSbAI6UnqvAiIgAiIgAiIgAiIQHwhIMEivjxJzUMEREAEREAEREAERCBGCXjzUDhhiBAOTpmQcMBeEQ5Iwk1Cb0QMhIcUVopaIUQU3hPVrBAiChGC63gP4KlRzAoG/RNWCEVV2gpCxiYrw73tm9mr4+WB0DHeCvk3clhBAPnHxsF1hBAn9BTnuc9VG/cNXhF2LlzHr+PHjHjtnS7dGzd/6llfweLc2bNnWj98fxU6xLuiWp36jT7/sONrbm8DfzcrWa5i1Q2rVy5LnjxFioFjf52FB0fbFo1qL/9j/hxED7wMnHZZst6X44vB30/Yv2fnjucfa1DjlF07dGDf3rc//vzr28014x87Qd2ylavXOvXXyROb1q1e6e+edR5s8miDh5u1nDh2xBD39Yi2ow8EC16Dl/2Xs6NQsZJlOnbp0WfujCmTECk++XrI6Op1GzwUkmDRofNnXz7Q+NHHP3vvzZd/HDm4P30gzjz65HMv4p0RrgelyiIgAiIgAiIgAiIgAiIQBwlIsIiDD01DFgEREAEREAEREAERiJ0EXCKGIwrgheEc1z0LTFDAI4PwUuTIIMk3B4Z1wkwds9LHSksr6awgfKy3stUKoajwsqAenh6IH45IUsP791l7xdPgiJWjVvDw4NUTZsruvdrGSdsbjhQmEjz7Svt3pk36acyeHdu2+F53/v775InjyxcvmFO5Zt366Uwh+NcUAn918bTg/Ma1/gUDp80dd2W4O29Q4aIDv+re5f3ufQamthBNzzatV3Xnts0bqYPo4O7//R5fDzRng2RvPNuiMWIF18yxIzWvVyzklFOXfBuEgvINW8V1PBle6vC+JwcHHiPu/iPajj4KFC6OV00iBAru8UGPrwfZNNa9/eIzzS5dunjxlbc//OTuTJkRom46ylaqVrN5qxfafde316eOWEGl8lVq1CFHh7wrQlqROi8CIiACIiACIiACIhCfCPAfPzpEQAREQAREQAREQAREQARikIAJBlesXLSCF8QeK3utbLCCZ8ZqKxOtPG7lUSuNrHxnBcFjlRXyPwy1glcGuRdI2J3dSh4rCBW8prWC2IEggsDhJPK+094XMtHihv8OwLPh62Hjfn382ZdeS5I4SZj/jYCHAG0QLULCVrh46bKHD+zfe+LYkT9DQ1uyXKWqhI9KkSJFytoNGj/y3qvPtXTECt92GO8rVK1Zl4TfB/fvxavEc+QvXLSEeVnscXJRJLGjaMky5TdvWBPs794PPPRIC/JsbNu0fq07v0VE2zn3KGDjIIzVgb27dz7c4unnyLPxYfu2zyBWUIewTv7GY3pLmg979ftux9ZNGwZ91eNjd52K1evU27xhbbCl6cCLR4cIiIAIiIAIiIAIiIAIxGsC8rCI149XkxMBERABERABERABEYjtBLz5JpzQUgzXeX/O3p8zcYEQR4SZonjCHdmxwsooK3dZQfRAnNhlJZsVwlBhGKcuHh7kt8BrI72VQt72eGxcPzCWFy5RplybZg1q7tq+hfBToR5L5s9GWPGEXfrNPDL8VSbM0+rlSzyhkUI7CKOEBwH5JqaMHzvyj7kzfwup/lNtX+uAh8fYYQO/cerksBwUtR94qCmeCc45klWnSZvu9u3m3eDbl6XKuK3N6506c9537BFtR1/JU6RMmTN3vgITLMQUYs6z7Tq898PwQX23b9noYW0pPJJnMPeKdauWL/Ed08OPP/M8oa6eeqhWBUfcoM5dGTJmQgT5fkj/3mFx1HUREAEREAEREAEREAERiA8EJFjEh6eoOYiACIiACIiACIiACMRbAi5Bwy1q4DFBforTJmgwd4QJPA7c+Rqo7yTidgQPvDLOu/NYkMuBJM+dXm7dYuPaYISQMI8/Dx3Yj/dEUOFinhBIvgfGd5Jmm2CxKKzO8hUsUozwSZZ+4s6+PT9+L6T6GS2TdbnK1WuP+LZ3zwvnzyHmJLo3W/ac/UZN+G3v7h3bhtt5p23BoiXI/ZHIBIsbhBnOPfRYy1b35cydl/e+OTgi2o6+8uQPKsw81gUvX9LosSeeMcEk3aDe3a97S2TNnjM31/fv2bXDPUe8S5o93ebl4OWLF64PXkEC9+tHxRq163GdpONhcdR1ERABERABERABERABERABERABERABERABERABERABEYjTBMbPXraBEt5J9B3587TFW/9ENLnpQAAxIeVa3gKFioTV78xV2w5Rl/wVodVt+OjjT1Mvd76gQnhJNH2iVZtFmw+emrpkw27EEXfbN97v9vnyXccvUM99ntwX05Zs3EM/Czbu/wsxICra0UcTCwFFv4SBmjhv1ZbWr7z5jrtvwl1xHU8S9/kqte5vwPlaDzR62Hf+3fsP+4Frd5lnRlgcdV0EREAEREAEREAEREAE4gOBMOPTxodJag4iIAIiIAIiIAIiIAIiIAI3E8C4jgAw+YdR5MQI13HcclOQewERwLdhkZJly5NzgZwMoXWKV0WGjJnvoc44C58UWl1yXZw4fvQIIZImL1i9DYFj8bxZM1rUq1zyyOGDJB6/fjCnA3t277Qc3DckF8fz4c4MGTIeP/rnYXJXXLMjKtrRRz5LHI7nB54UzOuHYQOuh63iOuGmeN22acNa9z3rPfRoC8Jczf196mT3ebhWqFqrLrk6wsoDEq4Hp8oiIAIiIAIiIAIiIAIiEIsJSLCIxQ9HQxMBERABERABERABERCB6CRQuHipsvS/cd1qdyipgG6ZMlWq1Fc9x5Urvg1IeE2uBl9BwLdeHq8Hxub1a1Y5uR5Cunnx0uUrkdOhW5/BoxAonnu0fvWOLz792D+n/nbyelxvSqiofXt2bnf3RQ6J59q99d740cMGpr/jzrvWBy+/IfwSdSPajrb5ChYutmv71k3Nn2nzyqjBfb88e+bMDd4nlt6iEPkpdm/fSlguz4GHR6XqtestmD19Cnk83OOtZOGgbjflY+3KZYsDeiCqJAIiIAIiIAIiIAIiIALxgIAEi3jwEDUFERABERABERABERABEYgIgTsy3J2RdifNcyG87e/LkTvPsSOHDyFZuNuSfBrj/YY1K5eH1Wf+QkWKU2fGLz+PC6suYZ/IsfFkwxrlnm1ar+qqpYvmh9Tmbst3YZrGPvf1pi1bvYBQsXDOjKmIF+t88kVQN6LtaIv4Yk4RyYOKlij144hB/XzHljt/UKGdWzdvdCfVJpcGY1q15Oa51G3YtBmCjz9hJSxWui4CIiACIiACIiACIiACcZWABIu4+uQ0bhEQAREQAREQAREQARGIJIHz586epYs77/pPuAj0uNOEDguBVAwvCt82ufLmDyKc0aZ1a1aF1V+BQsVKUGfO9F8nhlY3efIUKQg/tWLxgrmEcgqtbgpz/UiTNm26E0eP/OnUswTYt7d57e0Pxgzt3yfzPfdm47xv8uuItqMvEoLjDUHOjvGjvhtw5vTpf91jhEf2XHnybdmwNth93vEw2b5lwzr3+cxZsmYjoTkeGP6ElbC46roIiIAIiIAIiIAIiIAIxFUCEizi6pPTuEVABERABERABERABEQgkgSc8ESVatR5IDxdEfaIhNZTJ4wb7dvOBAtProZd27dsCqtP8lEgHPiKB77tbrecEJy7dPHChbD6TJ0mTVrqnD17+npIpjavv/3B1WtXrw7v37tnrnz/5ZIw55Ab8l5EtB195SlQ0JNc/PLlS5fGDht4Q+4KzuNJgWjhm9Mji8Wg8jeWdp0++uzQgX17Ll44f94350VY89d1ERABERABERABERABEYjLBCRYxOWnp7GLgAiIgAiIgAiIgAiIQCQILF+8YA75IJq3atsuR558BQLpKn+hosWffvH1jpvXrw1eaLkXfNtkyZo9B+fciaILFC5WAg8Jd13CMuU0bwy8JsK679kz/3o8FvCCCKtuCgtJRR2z9Z/jlXs/8exLr/ft3uXdM5YJnDwVlvbiJAmy3X1FtB19kLyc17nTp0wiobfvGAkHxbld224UcVKnTZeO86ZzXHLaFC1VtgIhtc5ZEgy8VBBBuJYkadKkYc1d10VABERABERABERABEQgrhOQYBHXn6DGLwIiIAIiIAIiIAIiIAIRJECi54/feuW5lClTphry07R5ZSpWrRFaV4WKlSzTf/TEGVcuX7nc5a2Xn/XNX0FbPC94TZU6rcfTocHDzVqOmbZgVanylau5+0aswOuAhNthDZ8E1ggBTgglpz6hn1q93L7TMyagOOcw9DvvLUrTnT36Dx+3bfOGtZN/HD2M8+ksdtNRE2l87xnRdvTjCBITx44Y4m8uJNzmvE3hoPv6qb9PnuTvLNn+E3nuznRPlu59h439qtv7byFcrF21bDE5Lng2Pb8d8WNYnHRdBERABERABERABERABOI6Ac9/TOgQAREQAREQAREQAREQARFImAQWz58949VWjzXs1nvQyEHjpszB42H2tF9+3rxhTfDJ48eOmv5wW9a5AOmFAAAgAElEQVTsOXPXbtD4kYZNWzx13jwXOr38TPOtG9et8Uds767t2zjf4cPPvjxx7OiRFq1eaLdozu/T/pg78zd3fbwI+HvtymWLAyH/2+TxY/GUQKDg3iXKVqj8yBOtXyB3RBcTXZw+/jH3CTwoHnvquZeeeuHVDogA7Z97vAkJrKmTOEmSJJZi4h/fe0a0Hf3kzJM/aN/unduXLpw7099ccuf7z8Pi75MnjruvW7LteYzrrS49+syeNvnnJ59v137ujCmTzBNjI3kx/rVBjZw8e4kNOcnnH3V6PRBOqiMCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACcZoAngdt27/z0bQlG/es3v/PNd+ydPuRs+zyJ6RSaBPFa2L4xJl/0D5436mr3fsNHWuRnFL7tnnj/W6fT5y3aguJpQMBR6LvXxet3eGMa9Wevy5/9d3YSUFFipX0bf/qO126U2/hpgN/V6xW63739U++HjJ65e6TlwhtFVXtvp86f0W1OvUbhTSPYRN+X/T7yq03eFc4dZ9/teP7cGK83foMHkXop+p1GzzE38yxe/9hP5A0PBBGqiMCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiAC8YoAokSVWvc3aNC0+ZN1HmzyaIkyFSo7SakDnSgCAyGbQqpfukKV6k7uh0D7JO8F7SpUrVmX/kNqh0cCgoQ/Qz9z+XLImIl3ZciYybd9RNuFNX7COmW6596sIdXDCyRvUOGiXMdjZODYX2at2vv3lUdatn4hrL51XQREQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREQASilEDh4qXKTl2yYTfeFRPmrNgUpZ2rMxEQAREQAREQAREQARGIAwSUdDsOPCQNUQREQAREQAREQAREQAREIH4TaNG67atDJ8xYuHr5kkV7d+3YtimAZOTxm4hmJwIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiEGMECJv1+YCRP5GvouXzL7+RPHmKFCt2n7j4+LMvvhZjg9CNREAEREAEREAEREAEREAEREAEREAEREAEREAEREAEREAEEi6B+3Lmzjtx7srNc9fuPlamYtUakAgqUrwUIaGKlylfKeGS0cxFQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREQARihEDOPPmDZgVvP/zrH+t2Zs2eM7dz0+atXmiHt0XKVKlSx8hAdBMREAEREAEREAEREAEREAEREAEREAEREAEREAEREAEREIGESSBV6tRpflm4Zvus1Tv+vDdb9pxuCj2/HfHj2N8WBidMMpq1CIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIhAjBFo2/6djwj7VK1O/UbumyZJmjTp/A37Tnbq1qtvjA1GNxIBERABERABERABERABERABERABERABERABERABERABEUiYBAgDRe4K39mXrVSt5n9CxgMNEyYZzVoEREAEREAEREAERCChE0iS0AFo/iIgAiIgAiIgAiIgAiIgAiIQUwRuuy1ZMsJAbd+ycb3vPZu0ePq5c2fPnlm6cN6smBqP7iMCIiACIiACIiACIiACsYmABIvY9DQ0FhEQAREQAREQAREQAREQgXhN4MqVy5cvXjh//vb0/7vDPdGgIsVK1n2wyWNTJ/ww+sL5c+fiNQRNTgREQAREQAREQAREQAREQAREQAREQAREQAREQAREQARE4NYT6DVw1Pjlu45fKFmuUtWUqVKlrlit1v2/r9x6cOn2I2ezZs+Z+9aPUCMQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREQARGI9wQy3XNv1imL1+8iX4VTVu39+0qjR594Jt5PXhMUAREQAREQAREQAREQgVAIJBYdERABERABERABERABERABERCBmCWQNt3t6clZEVSkeMlTf5088ctPo4dvXr82OGZHobuJgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIQAQIpL/jzrsi0CxGmmTOkjVbVNwoRcpUqXLkyVcgKvqKaB/p/3fHnXmDChfNkTtv/sR2RLQftRMBERABERABERABERABERABERABERABERABERABERCBeEegULGSZVbv/+datTr1G8W2yZUsV6kqYytTsWqNyI6te7+hY7/7efqCyPYT3vZJkiZN2qTF08+N/W1hcPC+U1eZD+X7qfNXIKKEt7+YrD/q17nLXnrr/a4xeU/dSwREQAREQASig0CS6OhUfYqACIiACIiACIiACIiACIiACIiACEQtgSIlSpejx0sXL1yI2p4j31v1uv+JKAgXkemtcPFSZe9v9Ejz82fPnolMP+Ftm/nerPeNnDx7yQc9vh505PDB/V3ffrVN++ceb7Jv987tBYuWKF2gcNES4e0zpurfbu4gcJMnSEwR131EQAREQASik8Bt0dm5+hYBERABERABERABERABERABERABEYgaAoQooqeNa4NXRE2PUddLibIVq9Bb0VJlK0Sm11c6dv6E9qf//eefyPQTnrZZ78uRC4+Oa3a0erhu5bUrly122ufMmz/o5bc+6HZw397d4ekzJuvmL1S0OPfbuXXzxpi8r+4lAiIgAiIgAtFBQB4W0UFVfYqACIiACIiACIiACIiACIiACMQ6AmnSpk3XvNUL7ZLedtv1zXt3ZciYKXuuPPli3WD9DChfwSLFDu7fu/vU33+djE3jtWhJqR0PhMjs9C9doUr1clVq1GZuZ8+c/jcm5sia+Hr4T1OuXrl65ZnGdSq6xQruX7x0+UpzZ0yZdPzon4djYjwRuUf+QkX+Eyy2bZFgERGAaiMCIiACIiACIiACIiACIiACIiACIiACIiACIiACMU2gzoNNHiUnQZvXO3Xm3uQs+HnO8o1dvvx2WEyPJbz3Y6xLtx8526P/8HHhbRvd9ctWqlYTrlMWr9/Fa848+YMics8Rk2YtdvJGvNn5sy8j0kd423Tu+c3gZTuOnnO8FNztg4oULwXzbDly5QlvvzFZv+tXA0es3H3yUrJkyZPH5H11LxEQAREQARGIDgLysIgOqupTBERABERABERABERABERABEQg1hGYN2Pq5AN7d+9s/fIbnTJmznJv42ZPtsa4/sOwAd/EusH6DCiXjZPEz5vWrV4Z28ZaslxFT96Kn0cPHchr0ZJlyod3jBWr165HOKktG9aupu2Z09EfEor7kWR7wFfdu2zduG6Ne8zJk6dI8VGvft8NtGv79+zaEd75xGT9oKLFS+3ZtX3rpUsXL8bkfXUvERABERABEYgOAhIsooOq+hQBERABERABERABERABERABEYh1BDDoDurToyuG/45devQhX8IvP30/fN/uXTvIYxDrBuwaUIEixUryZ2wULEqUqVD5/LlzZ3/58fvhjDEieSzatn/3o6t2jBsxuB99nDkd/SGhXn+va8+9u3ZsGznw616+z/697r0H/H3yxPERA/p8HpvXBeG4cubOV2Dbpg1rY/M4NTYREAEREAERCJSAkm4HSkr1REAEREAEREAEREAEREAEREAE4jQBwiqd+uvkiYsXL1yoVf+hpkzmwYebP/nQYy1bYSyvVzYo27Ejhw/FxkkWLFKiFEmhTbBYFZvGd9ttyZIVLVWuwqb1q1edOH70CB4s5LEIzxgr1ajzQJESpcvNnDLxpyOHDuz/T7D4N1qTbpcsV6kqQkunl1u3uHL58mX3eJ9/teP75SpXr/14/aqlWBfhmUtM1yWUFeva8UyJ6fvrfiIgAiIgAiIQ1QQkWEQ1UfUnAiIgAiIgAiIgAiIgAiIgAiIQ6whUqFqz7lsf9eidM2/+oIsXzp9ngBiq2V3/56GD+9evXrEstooVjJV8CngDRLchP7wPLsg8P9jlvz54xVLarrPX+xs+3AwvlgvmdhFIf3hXIMYM7tOzq5MvIro9LJ547qXXEVdmTpnwo3uMj7Rs/cKz7d58t3XTelVPHj92NJDx38o6hYqVLMP9TbAIvpXj0L1FQAREQAREIKoIKCRUVJFUPyIgAiIgAiIgAiIgAiIgAiIgArGSAPkIvh7x05R9lovgqUY1yx+wN2fPnDmd9LbbbmMH/Y8jB/ffvH5NlHsulCpfuVrBoiVKRxYKO+gLFC5WYuPa4BWR7Suq2+OpQJ/rVi1fwivCD1wRMgK5V+WadevjkTFn+q8Tt2/ZuD5V6tRpaHf+3JkzgbSPSJ1M99ybtXqd+o3GjRjUz+1BUb/JY090/Ljn12+/1Kp5bAy95W+usdXzJiLPRW1EQAREQAREQAREQAREQAREQAREQAREQAREQAREIEEQcAzhhPtZsfvExXwFixT7fur8FcH7Tl1t9OgTz0Q1hMbNn3p29f5/rs1du/tYZPvOk79gYfpq3uqFdhHpK0PGzPfcmeHujBFpG1ab3kPH/cLYuAd1ER/4Gw+GsNpyfdSvc5fxDPIWKFSEv5s+0aoN7ctWqlYzkPYRqfPCG+98uHzX8Qu3p//fHU57woKxLqJyLUQnd2fcP89ZvnHS/OCtEeFwq9vgmXNfztx5b/U4dH8REAEREAEREAEREAEREAEREAEREAEREAEREAERiHEC6cxCvWzH0XMkW+bmmbNkzTZz1bZDq/b8ddkJRRRVg2r9ypvvYHgfOmHGwsj2iTGdvoqULFM+vH0ltuOXhWu2v9ThvY/D2zas+vQ9f8O+k1MWr9/l1CWnBYw/6zt0TFjt8a5gXj2/HXE9LBNCh2eultMirPYRuZ7EjmlLNu7pNWj0z077Nq936rxy98lLDR5u1jIiffprE53cnfth8F+19+8rn3w9ZHRUjTsm+/nw875Dvvt5+oKYvKfuJQIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAKxggDG6joPNnk0WbLkyZ0BkbT4nU++6Jc6TZq0UTlIDNa58wUVct8rov2/++mX/TGoJ0+RMmV4+yhaqmwFBIBaDzR6OLxtw6qPVwR9d+szeJS77vCJM/9AJAmrPd4VGNxz5S1Q0Kn7bLsO79InXiVhtY/I9XJVatSm/xr3P9j4rgwZM/Ue+sPkRZsPnqpYvXa9iPQXUpvo5O7cEwErMp43UTnf8PZFmDa4v/3x51+Ht63qi4AIiIAIxG8CymERv5+vZicCIiACIiACIiACIiACIiACIuAlQL6CmVMm/nTp0sWLDpStG9et+ey9N18mp0VUgiKJ9M5tmze67xXR/gsVK1XGulrnJAsPTz/lq9SsQ/3g5Ysj7enhe99S5StV49yalUv/cF9bF7x8CR4rFnHpzpDGWqlGnQcIHzV98vixu7Zv2eTUS5EihUeUOWcPJDzzDLRuw6Ytnjr1918nEZR+nrtiUzXLZXHi2NEj2bLnyh0V4pIzjujk7tyjQKFiJXi/YfXKZYHOP7bUK2weNGnSprs9OtZlbJmjxiECIiACIhAxAhIsIsZNrURABERABERABERABERABERABETALwEM3+EJ3xSa5wQ70fMVLFxs45qVyyOCO0/+oMKHLMv4XyeORzqXhu/9S5StWIVza1fcKFis9SbgLlSsZJmQxkweiSuXL18e8OWnH7nrpLA4R/x9/ty5sxGZb2ht4FzdPCtmTZ00HrFk9/atmxfN+X3a3ydPHO/UrVffEZNnL/nfnXdlCK0PruM9kfnerPeFVi86uTv3LVC4aImLFy9c2Lpx/ZrwsAp0DuHp07cughDJ10Pqw/Gg2RDAukbYiOhYCFEW0bZqJwIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAKxgkCSpEmTvt211zdVa9d70D0gQiuR/6BF67avhjTQJ59/pT2hegg3FVIdjLnPtXvrvVnB2w9Td+xvC4P9GcvJ5cB1dzJoQhm1bf/OR+QAqFLr/gbue2AofuujHr37jZrw21ffjZ00b92e47NX7zzSa+Co8ZTu/Yf90OqlN96OCsjk/1iwcf9f3NPd392Z7snCmElw7u8+eFdwvXPPbwb7Xkc44Fp4QnTxjPoM+/HXb0aMn+ok7/Z332p1HmhI3/7CP9EH4am+GPz9hJDYtHq5fSdCc9EHhXVAHgnqRxX3O+7KcDc5Vr4b/9v8F998t0toz4mk8YTVos5dd2fKTOgwcqa80rHzJyF5i4Q2h5DuVb/JY0+M/GXO0kWbD/1D/g8+F+Qf8Vcfrxqe6x9bDv+7bOex86xxp17jZk+27jd64nQStU+ct2oLydaddUkeE56973MnKTf9sGboh8/lUy+82mGkiUvMFQ8Z33FQh3n+vnLrQZ7pl0PGTPTlUaZi1RrvfdZ7QGh8GYvv2o6Kz436EAEREAERCJ1AiGq3wImACIiACIiACIiACIiACIiACIhAQiWAUND8mTavZM5yb7YFs6ZPgcNjTz3/EvkueI9wcfzokcOEmPJldPTIn4c4l/W+HLkIOeV7Ha+J3sPG/VK+So06c6b/OvHUXydPPPz4M88/1abdm193/+gdd/1C5gnA3+u9YX+Klylf6ashYychbhB2qpEl5H6hecNaK5csnEc9DOhBRYuXOnv69L8YW9Pfcedd5mCx656s92VPZlZb2hw/cuRwZJ9r1uw5c2fImPkePBTo093fsSOHD/158MA+Z+y+93rxzfe64BkwqHePmxKBW0QoT0ioQDws2D3/3mdffdu4+VPPOvcglFTHF59+zN/8MG6fOf3vPyv+WDDH9zrPeNqEcaMffKTFUwhNvs8tqEixku3e/vDTLRvWrZ47Y8qkmvUebMIa2LRu9cqhfb/4LCq482wx4CM+ML6S5SpVnfHLhHHukFnOuDHK48UxYezIITny5CsweNyUOTxrQpuVKFOhsjn5JP+q2/tvuecZ1hx8mXCPrl8NHIFgwXP+xtZm7vwFCvG5ML0tGefcbTLah2XIT9PmsS5+Hf/9iKDCxUu+aMnep078YfThA/v34plCu7On//0XUesfC82V+d5s97EuE1t+mdRp0t6URwYBis8LawzGCFNlK1WryZrOmClzlkeffLbt/JnTfnHGwZroNWjU+Kq1H2jIZ/NaomvX7m/YtFndRg83m/rzD9dzrTzz4usdfdetey4FChcrwVzeeaX14wtnz5ga2c+L2ouACIiACIiACIiACIiACIiACIiACIiACIiACIhAhAm0fP7lN9hF/6SJCHRCeCN217Nb+4HGjz7O7vBPvh4y2t8NMGTTFkOyv+tdvvx2GO3rPfRIC+c6xtFlO46e8w0P9VnfoWMWbjrwN+IDxlt2rv8wfdFqElXnK1ikGPfp0X/4OH/3wXDNdV8vkQhDcTXE44O+2cnur7/u/YaOxbPD95rDBi8Qf+0+/ea771fsPnE9x0hIY8UwzU59xjBw7C+z8gYVLsrO/zlrdh19ueMH3fy1Y8c94wqpT7xV6O/VTh995lunY5eefbiGoZ1rqVKnTgN3f2wjwh0j/JJtR87wfBEEELtYb6wL5uY7npymVjCepk+0aoO3wqT5wVtpw7hgsHT7kbMIDu524ZkD7ajPOkWoc/opXaFKde7rXrtc43ng7YEXBsZ+zjlJ2WvWa9jEPQ68i1jr7T/4pFdYa5F1snzX8QumZaQjQfqqPX9dfuK5l17n88BcnRBiTj8dPuz+FeNr0uLp5zhHPbyMmItTh7Eu3vrn6ZC8pEw7SfLjzCXr8M7InCVrtrDGqOsiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiEK0EuvUZPArDJ54EGH4RCcZMW7jKCS0zdcmG3YNsV7u/QRCSZ9Hmg6f8hZNxDPa+RnF2nzviiLvPKYvX7/p2zOTf2V0+ecHqbRPnrtx8u8Xdcepg5CZcj79xPP7si68xB2fHflQC+7BXv+/oG68Af/1iDOb6vdmy53SuYwj+ec7yjRjl78xwd0Z/7QjJxPWwxvp+9z4D6Z+wPvRLfYQKzmFs9m2P0Z9r7LYPqW/GRB3CFvnWQRxBQAhrXFwPL3eELdbL3LW7jzlhxBCuMM4zHtaM731rN2j8CNc+HzDyp/kb9p3MYmqFU6fvyJ+ncQ1PB3e78MwBAQWxwlf8YW0zLksrkd7dd+tX3nyHe9Z5sMmjznknnBmhuNx1HaHt/kaPNA+L5/jZyzYM/nHq3GZPt3nZV+TzbVusdLmK1HG8oJzriDftO3/6hfM3nzXGSh4Tf/fHo4TrcAxrfLouAiIgAiIQ9QSUdDvqmapHERABERABERABERABERABERCBOE6AhMZ7d+3YdmDv7p0P225tkgR/2L7tM5cuXfTs/ie0TUhTJOH2htUrl/uGnCG0TYePuvc+cvjggUF9enR1t19niapHDfrmulGVaxjQMfivX71i2SsdP/zENvdnfbNNy6b/nPr7L6ct4XQsytEpf2MpXLx0WULxnDh25M+ofhzFS5evdPHC+fMb1wSv8Nc38+G8O/l4g6bNn8QzZMzQ/n1OHj921F87QkLRb2jjZcc/ngWE+Pn03TdevGoHu/YfaPzY47RbPG/WTYJDxWq17r965cqVxfNnzQipbycxuW3cvyk0EeGLuIfjYRHa+MLD3ez+/+v93Q+T8QVo+/hDdZxQVPXNiwehjMTkyxbNm+17PzwsOFetbv1G3Tq99gKJ1Z06p0//8w/vT/976oZ1Eegc8FxAkNqxddOGQV/dGLarYvU69TZvWBvsXnPkrWj98pvv/DF35m/uEGn5vZ4W2zdvXO8evyMUrA9e7ldoc+oS9ix3vqBChMRq1+nDT4d/27vn9MnjQ/SQef3drj15hn0+7Xw9RwtiEF4Y2zdvuC5iFStVriJrYdvmjTcJWzB//rW3P2AMP38/bFBUf27UnwiIgAiIQNgEJFiEzUg1REAEREAEREAEREAEREAEREAEEhABdrfnzJ2vwIrFC+YiMjzbrsN7Pwwf1Hf7lv8Mr3hZZLA8A+Se8MWCwROD9brg/wz27oNcC4SY6fd51/cDydHADnXak4+CMEH9enZ9353PgL4wou/bvWO7v8dTslzFqmtXLVsc1Y8OQ3KO3Hnzk1fDEXB877F14/o1CA9mHK7ANYzGL3V4vytiy4hv+3we0pgMd8oLoQgW7I7v2KVHH+79UYeXn3VEIcJ0Od4cy/0Y+MtVqVF749rgFabt/B3Svenr8mVmdOGCb51li+bO4pxvkvPIciesWPZcefK9/9rzTzpiBWsIjwX6JkeGP0EqV97/BIsVixfO9c2jkjbt7bczB981FugcyKeCx0bXt19t436+JHtHyFu9fMki97ybtmz9AiGb+vfq1tk5z/MmJ0vwsj8WuMUUrpOb4/jRPw/7nvdl6Qgb5KM4cezokQFffPphSM+OdYG3z4gBfT4nj4dTj8Tv5C2ZN2OqiUL/HcWsLmKkP2GswcPNWrK2Ya7cFVH9zaH+REAERCAwAhIsAuOkWiIgAiIgAiIgAiIgAiIgAiIgAgmEAMmMMRojOjR67Iln0qRNl25Q7+7XE0Q7YaL279m1wxcJnhip06RJu2blzUIBogMix4zJP/8QCMrCJlhgRCdZ9E7bDv790G+vx+Gnfd6gQp7cBts2bVjr2x8G50z33JvV17gcyH3DqsMOdepgjA6pLoZ/24i/gjA91CEnCAILBuWQPEKo95+HxQW/HhaIM4SCOn/+/Ll3LRky96ANz6qNd1c8vJwE5c7YEJjIK7F04ZyZoc2N/slv4G98s3/7ZQJixyNmnA+tj/Bwr9vw4ccQQH4cObj/vN//36CO0Txbjlx5uM+64BV+vRBy5snnESwGfPnpR77jQVA6uHfPLt/zgcyBMGae8EvLFy9c73PvijVq1+P6mhU3ChbkM6Eu4gr3JHyZkzy8+/sdXvEdR8myFasEsi4JHUVb1s03Pbq8609IcvpmDAgQE8eOGOKce+GNdz4kvNPnH779uluoKli0ZGlHfHSPjWfftv27Hp5LF8yZ6ayvsD4Pui4CIiACIhC1BCRYRC1P9SYCIiACIiACIiACIiACIiACIhDHCTh5BDavW7PqiedefoNQNO4wTLnzBxViirt2bN3sO1V2emM0d0IiOdfxlshpu+J/+en74aEZXt39FSn+n2CB0b/HB2+1I4yN+7qTjHnbpvU3CRZObonVZniO6sfBDnX6DF4Wet8YsfMXLFIcgafVS+07EQZq7NBvvw5tPKF5WLRo9UI7Ejl//mHH1ywC0nWDfNPHW7XBwI9HwcH9e3f7elGwUx8j+tIFc0MVLJzcIOz+9x0jff8wfGDfoCLFS+GtEdIcAuWOqPVm50+/3LNz+9YvPn7Pk9idA++eF9u/18Xxjti8YU2w770QDbLnyptv9/atm31FBerelzN33m1b/j8EktM+kEFi5PYAABUrSURBVDlUrlm3PizHDOl/U1L0SjXqPEBfbjHunqzZsuMhMnXCOE8CenJfjJuxeE2ZilVqvPn84w/7CgMZM2e5lzYIImGtS541dWA0e9rkn0OrX6FarboLZk2fwrNn/P1GTfitbft3Pur/ebcPJv84epjTFu6Z7816n310N/j291Czlq2cXCDR4ZkU1nx1XQREQARE4D8CEiy0EkRABERABERABERABERABERABETARSCfJWgmng6GduLz/zBswDduQORh4G9/ng1FS5QpjzeE7y79GvUaNqHN779O+DEQ2BilCxUvVYaE0rOmThrvz8Br4f2Lkr+BXAO+fRYpWbY8Y/B3LZD7h1YHAYXcCmEZdTGm4/3w5ZAxEwkZNLTfF5+dO3v2TGh942FBTCbfOiQOb2uG/M3r1wYj+jjXSf784pvvdiFHwaEDe/fs8IbtcrcvVb5yNcIErfUTpstdj+fN34QL8jfGUQO/+YLwQq1feqNTSHMIlHub1zt1xnjf+5MPOrpDEz3Z5pX2GPTnz5z6C/fYsWXTDfkfOJcpy73ZEGCW/TH/ptwWzIG8GP7WJm3DmkO9hx5t8ffJE8fnujw+aIf3QYWqteoiCLlzohDeievnDPB3P09fMPCHX2fz2XmiQfUySy1a1c3rskx5zq1dufSPsNahCYOFqTPOhCLffDDutnhgIDTw3Lp+NXDEpHmrthQsWqJ0++cebzL4657d3HX57PLZ2rtr+1b3eeZHGC5y1nA+JM+WsMas6yIgAiIgApEnIMEi8gzVgwiIgAiIgAiIgAiIgAiIgAiIQDwikK9g4WJmz9xECKdRg/t+6Y6JzzQtvUUhYvuzw9132hjz16y42RhbrnL1Wuz+dsLmhIUrh90EYzzCAOFw/NXPF1Sk2L7dO7f7y4dR1BJ/4+URmqE3rDH4u07YJELqkHg5LPFhrTfxNjvlj/556OBPo4YOCOueyVOmTGmRnjyhntzH021f7YDo0eezzm+75/Tim+91ueOuDHd/a/kNYObvmZQsX6kq4b1gGdr9nR395N/wV4/n9+OIwf3L2rN0vFt86wXCnfGytlZbaKX5M6d5hAkODO8kr+a85WXfxzzxLvC9x3058+TlnL+5lqlYtQbXLOn7svDOAUN+peq16y2YPX2KrzdPJQsHhQfKWp9QZyRf5z5dvvx2GALMh+1fbNX8gSolEe383R8+rBvT2G7yCnLXR0CwsFcF+Jz9NumnMaE9t2LeMViumXer39/goe/69vr0wUpFc8+dMWWSb7t7s+XIyTk+N+5rjZs/2fp/9mD+mDdzOvfcYsJYWGtV10VABERABKKHgASL6OGqXkVABERABERABERABERABERABOIogTxmYDd7afKgoiVK/ThiUD/faRASaufWzRt9E06TO4BwPGt8do9jfEUEIYQSHhGBYClcolRZ6k2dOG60v1wZJAMnFM8WEw58+yOsEPfbsGbl8kDuFZ46GPXZ3R9IqClCK/156MB++h/yda9P/CU5vmnsNrFL3twUzjXC+DR9ovULCDDLFv6X/JqD3f3NLUwUXisnLSsz3ih4ALj7xMOjaMmyFfyJSL73JrcC4o+/MEtO3TFDB3yNMb9xsydbR5T7Y089/xJJqQf37tHV6QOx4KNe/YYmS54sOeG/ChQuVgJPBrwVfO/jhC3yF7qKnBi08ZdDJaw5sHbT33HnXatMR/G9Z92GTZt58oMEL78hpwZ5UvDI6NCmZdOHqhTPi/eLr9jh7quICRab169eFVod6ufKV6Agn5tlC+fNsjztJ0Nbo5nuyZKV6192fa/D/WXyZ+3f65POeML4a5Mx8z33cv7wwf37nOt8Xp5/reMHeFIhGnkSxvtJvB6ez4nqioAIiIAIRJyABIuIs1NLERABERABERABERABERABERCBeEaAXeLsJMcwP37UdwPOnD79r3uKGFFDEgrYPU7dtT4eFlmy3ZeDdod8jOmhoSPnBdcZg796ufMXKIQxfvP6m3Mc5LJcGdxvk+XgiOrHQz4I+ly1NOSE2+57mlCwiN3sk34Y+V0gYyFBtq8nRM0HGj2MaDH++6EDnT4Ie/TxVwOGHzl0cH+3Tq+94HhHGOM97vsQ3gvPDF8RyXcsCEDszicUU2jGakQCQh1VrV3vQd8+AuX+4CMtnkJYcYdMQnghN0afTzu/vXXjujUWuajIof37bpiLcz/TFDLwHqHAPQYEM3JQLJrz+7TQxKGQ5oBQR3/bffJfYMQPKlysJKKKb6gki5h2F/lESOgdiBjHcwpkXRYoVLQEY5kz/deJYa0bxkCdH0cO6e/rDeXb9s67M2ZifZ366+QJ5xoJ4dOkTZdu5KBvvshfsGhxfwJhWGPQdREQAREQgagjIMEi6liqJxEQAREQAREQAREQAREQAREQgThOII8ZipnCZdvlP3bYwBtyV3CeXeiIAf5yQxQrVa7iieNHj7gTQtOGEEC8HvOTzDkkXIWLly6LYXnDmlV+vSTyFihclLbkbvDtwwznnhwbu7Zv2RTVj6NQsZJl2Gm/xsIWBdJ39w86tHu6ce2Kvt4oIbUl5JQ5MNwQuqlKzfsbYAyf//t/4ZMQanp8O2KcbZbP1umVVi0I1cRz4ZpFnvJ4dDhHibIVqrCb39czwPf+9R9u1tKM1rf/MHxQ37DmhbcGuSLwknDXDYR7zjz5gyzdQq55M6ZOdkJbEcbpzQ8+/WLh7BlTv7dk14gz5OxwvFN8x2MOAZ77njt35oZ8II+YFwqCjzvHR0hz8TcHS42RnfpHDh864G7XrtNHnx2yRY0I4psb43ZTCwL1RkAMJMxZIOsSDxPGsHjerOlhPQ/GQJ1LAXhFwNYiUp12+sxgLheE4Rry9eceDyASch+xeFxh3VPXRUAEREAEoo+ABIvoY6ueRUAEREAEREAEREAEREAEREAE4hiBPPkLehL9zp0+ZZK/kDuEg+L6rm03iwGEuyFske+U2ZnOuVQWSsn3Wo7cefNjnHafZ7d/XkuoTTickHJQODkUdmzdfFPC7SxZs+egP3dyZAzAqVKnThPZx4FgQX6CsML0OPdhJ7uvJ0BoY0hqioVvDouCxUqWxkvDdIm/YPlO1159K1StWfeLru++6fC20ETZ6Nc32XmJMhUqbzNRh1BHTlJt3/tjSG//wSe95lmiad/QUTwbPGrcbRJb6CkEFN+wRoFwL1isRGn6Wu/NMZHbMqd/PnDUeAtRtPeD19s8xbVMlnXb31ycMThzdAsmJId/8oV2b+7ZsW0LHhbu8QY6h9TmZUA7N/+ipcpWILwYSbXxjEDIow6iEa9m+//X9JMbhJuQni+eRr7rkvBWhJXybZO/UJHiPPNAxAPGQHtHyAltfRH+yR1mq1O3Xn1PmsiIUOTktwjknpH9HKm9CIiACIhAyAQkWGh1iIAIiIAIiIAIiIAIiIAIiIAIiICXgCNITBw7Yog/KCTc5rw5Pxx0X2dne5ESZco5hmj3tf17du/kb3IuuM/z9w/TF61+qFnLVu7zGIjx4li5ZOG8kB4MdTC8HrPt8L518FLgXKrUadPy2sC8B8ZMW7CqVPnK1SLzoDH25rJYRcHLAgsHFZF7IUiYg8UNHhaEQEL04Nr73fsMfOTJZ9sSKmus5ZNw7mEaTwrenz3z7w0hvMzDovLGtcErBo2bOueb4T9NQQxyjwtjfu+hP0w2o/fpbm+/9oLvmN/99Mv+wyfO/OPODHdn5Bo78h9+/Onn165attjXayQQ7tfDOf114nj+QkWLD/lp2jzm1e6ZRx90RCBnLme8hnjfMe3dtWMb55wQTuTu+LBXv+8IZdb70w86+oZmCnQOp/4+6ckVkSXbf4LX3ZYconvfYWO/6vb+WwgXzBnhhzH3/HbEj9RhLHi3uLkyHtYcY3KPHTHKvS4JDzV2+qLgFq3bvuo7R+ZGrotA1pAvD6cNYlXXrwaOwGvCOXfe3Cuc9yQ+r2Xhxr74+N03eZaEGePaUR8Pk0DGoDoiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiEOUERv4yZ+nkBau3OV4Rvjf4fMDIn1bv/+faXRkyZnJfw1OC86++06X7mGkLV/nmOOg3euJ0rrOju2K1Wvc/267Du0u3Hzk7a/WOPzGCu/siKTN1MWiHNME5a3Ydnbduzw05DJy69R56pAXtP+s7dEyHD7t/tWrPX5e/NmN9SHMKFGLBoiVK0+/9jR5pHmib8NZbvPXP018M/n6Cu93EuSs3r9x98tKvi9bu4P5fDhkz0dnh79Rr9XL7Tlz7ZsT4qY7xnN37nHukZesX6IP3A8ZMnvlA40cfp3Ts0rPPos0HT/36x7qdOfLkK+BvrA0fffxp2k2Ys2IT912wcf9fS7YdOYM3jW/9QLjfb8mr6W/ako17eP70hWHd3RdJzedv2Hdy4aYDf/vLlYE4Nnft7mMzVmw5gNG9//eTZtCnr0Dg9BnoHBAQgveduvrdz9MXPP7si6/9tnTTXhiRw4L+WbN8NngOztqsVueBhlzr1nvQSNY14gOs/I0HAYT++Yy1eb1TZ9YwHJyQac54ERhoT16PQNYPIsryXccvfD91/gqSjjdo2vzJb8dM/p0+xs34Yw05TJx+GB/new0a/TNj+fjLAcOdawiIXCtbuXqtQO6rOiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIQrQQwelarU79RSDcZNuH3Rb+v3HqDdwV1ic2/bOex8xg8ESec3dpOP4QVwsDMdaeMnDx7iZN7wX2/tz/+/GuMqRh4/Y0D4QGD9cR5q7b4u453Bl4B3Id+uvcbOhYjeGTBYQhesfvERV+BJbL9utvPXr3zCON1n6tZr2ETzmPgRhBifr73ZH79Rk34bdmOo+ccbwhHQEBogfPY3xYGu/k7/fk+K3ffsHaeB3MfOPaXWU6Cb98xBMIdLxXGiVAxYtKsxU5ydd++qtdt8BBiypudP/vSH18EF0Qc5xl37vnNYMfDw7d+eObw/Ksd32fNeESIPoNHIQwxFv5G+Oref9gP5Ppw7kHfeKi4uY6eMm95rfoPNfU3bkJvOXUR9vyF6UJ0YG5uz4iw1tiTbdq96R7Db8s27Xu67Wtv+XrU8Jmat37vCeoijLnDamXLkSuPR8ywEF1h3U/XRUAEREAEREAEREAEREAEREAEREAEREAEREAEROCWE2A3t7+Y+wyMvBJODgx/AyWHBMZfDP9BRYqVDGky5FQg9FJok7X8yDlDEjScdhju3bvLIwuPPAnFSperGNl+QmuPtwGMI3oPt9Ee7wBEBrfRmudTsmzFKghI4fE4gSMJmwMZV1RxRywIbYyW6iI7xv2QcnP4jjXQObCunBwphJlCpFm19+8reKqENP+gIsVLMRaM/mExQtz7n4X5CqkenjH0FVY/vtfhgEcK+Vp8PXDcdbk3uUP89Y/wE9o8wzsm1RcBERABERABERABERABERABERABERABERABERABERCBRHgwEBJIKCJGoHDxUmWnLtmw2wmJFbFe1EoEREAEREAEwkdASbfDx0u1RUAEREAEREAEREAEREAEREAEREAEYjkBdtjnL1Sk+OYNa4Nj+VBj5fDI9TB0woyFq5cvWURS603r1wSUADtWTkaDEgEREAEREAEREAEREAEREAEREAEREAEREAEREAEREIFbRYDQT57EzZaU+laNIS7el7BRJJYnX0XL519+g3BahNUiCXdcnI/GLAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAK3lECDh5u1RLAoWqpshVs6kDh0cxKTT5y7cjMJ3ctUrFqDoZObAo7Fy5SvFIemoqGKgAiIgAjEYQK3xeGxa+giIAIiIAIiIAIiIAIiIAIiIAIiIAIicBOBfAWLFLt65coVi2W0VnjCJpAzT/6gwT9OmXPu3LmzTzaqWf7A3t07aUWSdThu2bB2ddi9qIYIiIAIiIAIRJ6ABIvIM1QPIiACIiACIiACIiACIiACIiACIiACsYhA3qDCRffs2r71vBngY9GwYuVQUqVOnabPsHG/JEqcOHHb5g1rH9y/d7cz0JJlK1bZtnnDOnGMlY9OgxIBERCBeElASbfj5WPVpERABERABERABERABERABERABEQg4RLIW6Bgka0b169JuAQCn/nTbV97K1uOXHm6dny1jVusIHF5uSo1aq9dtWxx4L2ppgiIgAiIgAhEjoAEi8jxU2sREAEREAEREAEREAEREAEREAEREIFYROD29P+7I0PGzPcoHFRgD6VB0xZP7tmxbcv8mdN+cbcoXb5yNVgumT97RmA9qZYIiIAIiIAIRJ6ABIvIM1QPIiACIiACIiACIiACIiACIiACIiACsYRAngKFijAUQhnFkiHF2mHcdluyZPdmy55z+5aN630H2aTF08+dO3v2zNKF82bF2gloYCIgAiIgAvGOgASLePdINSEREAEREAEREAEREAEREAEREAERSLgE8noFi+2bN0qwCGMZXLly+fLFC+fP40nhrhpUpFjJug82eWzqhB9GX7AEFgl3NWnmIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIhBBAu937zNw7trdxyLYPME16zVw1Pjlu45fKFmuUtWUqVKlrlit1v2/r9x6cOn2I2ezZs+ZO8EB0YRFQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREICoIjJ4yb/mgcVPmREVfCaGPTPfcm3XK4vW7Vu//55pTVu39+0qjR594JiHMX3MUAREQARGIXQRui13D0WhEQAREQAREQAREQAREQAREQAREQAREIGIEkiRNmjRvgYJFJowZMThiPSS8VkcOHzzQ/P5KJchZEVSkeMlTf5088ctPo4dvXr82OOHR0IxFQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREIAoI3HFXhrvxFshXsEixKOhOXYiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACPzfRkNgNARGWggAAKJoYnTvO13VAAAAAElFTkSuQmCC"},{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOydd3gc1dm375nZXtV7taplyUVyr7KxKQYDBgOhkxDCy5dAKqRBCkkIqZA34SUQEkJJINSYZgM2tsG9d1m2el+tpC3aom0z3x9ryziAkYnBTjT3dZ1L2p2ZM2dmd357zvM85zmCRqPZoyhKCSoqKiofgSAIDYIkSYFYLGY8041RUVE5e5EkKSie6UaoqKj8Z6CKhYqKyohQxUJFRWVEqGKhoqIyIlSxUFFRGRGqWKioqIwIVSxUVFRGhCoWKioqI0IVCxUVlRGhioWKisqIUMVCRUVlRKhioaKiMiJUsVBRURkRqlioqKiMCFUsVFRURoQqFioqKiNCFQsVFZURoYqFiorKiFDFQkVFZUSoYqGiojIiNGe6ASqnhslsQavVoqAQCgYJhUJnukkqowRVLM5idAYzU+csYNqsuZRXjsdutxEJh/D7fIgaDRaLFVEUaGs4xIZ33uTN1/5JIKiKh8qng7oUwFmIJTGV62/9OvPPqWX7+tVsWreGA/t24x5wISvKCftqtHqKx1ZxzkWXU1s7h/vuvJVdew6coZar/LciSVIQSZICgKKWs6NUTlug/OPtTcrnrr1W0es0p3Rsbsl45fnVm5W0ZNsZvw61/HcVSZICkiiK31cURYvKGaegYjI//cV93HXzlWxYv5FYTD6l470DDvRJuYzJsOAKafn9k8+jj3k5cKDuU2qxymhBFMWoarM4i/jyd3/KA3ffTmt71ykdJ4gSNrsdAYhGwiQnpXDrndfw6t8e46obbuHNt9Z84JhwaIhAIHCaWq4yGlDF4mxBa6cs18qmbXtP+dC03BK+88MfIwjx16JGx4QJ47Fqo6QXVvCj3z78gWOO7FrPQ//7+3+31SqjCdVmcXYUQZegvLpuoyKchrqSCyqVRx9/XAGtsnztxjN+bWr5zy+SJAXUoKyzBCXsZl9DH5desvjfristLQuHowtjUib+AcdpaJ2KCqgGzrOIHZvf4//d8yuqKorp7mjD5XJ9onryx00kP8mIw6eQk2rinVXvnOaWqow2VAPnWYa7t4Pbrjifcy6+ktt/8Bsy0lNoaz5Ce3MTvY5u+p199DsduAecOHt7GfR6P7QenVYiGpGZUDOV3Vs3A6DRm7njuz/k6d//jN5+z2d5WSr/JahicZYRi4Z566Wneeulp9HpjeQVlZBXMIb0zCyKK6qYmjSf5LR0EpOSMZvNdDQf5o0X/8aqt94eriMalZEkkZlz53L/l38HwOJrbmXqzNm075vD8y++9iFnFigZN56+rhZcruNiYrZY8fsGP7yxgojJZCTg93/oZoM5gYuWLuX1558mGIqc9Lr1BhMWq5l+p/PkN0jlzKEaOP9ziyhplJKqGuW3T76qfOlLXxh+v2zKQuWx515V/vTkU8PvXfGlO5U3tx9R3ti4R3nlvZ1K1djiE+q69fu/VR5+8jnluTfXKTaTTgEUS0qO8sLb7yoaAcWWWaTce/99Jxyz6KpblW9/99sKoFx04x3KogUzT9h+9++fUf722rvKRRcuVBBE5Ss/elB5feMepXpCxQn7Xf7Fbygvrt6sPPrcCuWhxx47LUZetZzeoho4/8ORY1GO7NvBj7/zdRZefNnw+12tjVRUT+elpx4bfu/5R3/Fjr11/OjLV/PiKyspKhkzvE1vTeOCc6bwlRuvpMMVIiPFDsC5S69h3St/J6pAemYuFqP5fWcXWHb1dbz09ycAKBxTioA0vDVn7BRK0zS89trb6I0GLrj6NnKsUX73vw8xffqs4f1mLr6GhbMmcN3iOdx27aXc/5OfoBzdNv+8C0/j3VL5d1HF4r+A5NQMvAP9w68He1s50tDEnt27h98rmzyfXFuMnXvryMrKobuzc3jbZTf+D77ebipnnk+KJkBjhxNJZ+Kq629kx+YNAKSkZzIYcA8fUzq5loJkiYbWnvj2jBO3L73mJl597imsKQkIooWbbryK+390D0aDhcGgDzhqR7nruzz24M8IhiIsueF2zl80F4DyKedw7XVXfQp3S+WToorF2Yio4dJrbiI5KeFjd80qLOfun/yMxx9+f4CVzCsvvcR1X7gFAL05gW//8Cc8+JPvE40pmM1mhvxBAAorp3LJ4vlYCyZw++238N2v3EJMhhu/+gMyk20oMRkQWLj4YnJzi+L1mWzcdc+PiYbjdghLcibTpk0h7+j2iikLmDIul+XLXyM5OZ2LrvkCL//5AdyDQTRaPYoSA+AL3/wxuRlJBHyDaPQmLr7sCuRoDFGj5xvf/wEP//rnp+mGqpwO1FmnZyOCyLIv3MHlV15Ff3cLe3Zso7W5iT5nL4qiYDTbyMkvZNL0OWSlJ/Lw/T9k85ZtJ1Sh0Zv5zV9fwNNRT27ZJNa9/Gf++viTAFxwzZe5eNF0NmzeycXLruDer95E3qRFXLZkAa8vX864KfNIt8g8v3wVt9xyE+09LmRPO7b8STib9jCmcgpvPPk7yuZdgTEyQG7ZeN586RmWXfd51q9dQ83UKXz/tutobuvi/sdfZVy+jWXnzicUlSmtmce9995DQ0sPJryseGcrN3/xRsIxCUWJsvrvjxBJLqMkFe794b1n4OarfBiSJAVVsTiLEQSR/JKxVE6YRF5hERaLBUGASGiIjpZG9u3cyqG6OpR/mbZ+DEmrp3raLAb7Ojl0qP79NTP73IvJzkhm7cpXcPT2AVBRM4uJEyfQ09bAutVvE5MViismYrfo2bltC3qjjZrpM+hsOkRLSyuSVk/NjNk4Wg/T2tpOdkEphYV57N66Ad/RnktuUTlCxEdbW8fw2UurarCZtOzcugVZUUjLykUOB1m47BbKCrOpGF/OFy+/kMGAmpvjbEGdoq6Ws6pcc9vdyvr9TUpVRckZb4taTiyqN0TlrEHU6Jk+bx5P/+F+9h08cqabo/IhqGKhclaw7JZvUllWiKu//+N3VjkjqGKhcsaxJGdz5eUX8szTTyMK6lfybEX9ZFTOOJde/yVWPPMIXv8QAsKZbo7KR6CKhcqZRdBw4UUXsvyFF9BIOiLyyeeQqJw5VLFQOaPkltcw2L6PPk8Ag81G4H1RoCpnF6pYqJxRxk6oZu/OrQCkp2fg7FaT9ZytqGKhckZJzUilt7MdECgpLaKxoelMN0nlI1DFQuWM4h5wk56dy8S5FxF21NE/OHSmm6TyEajh3ipnFHNCGvf94TFMUpT7vn07zW2dH3+QymeOOjdERUVlREiSFFSHISoqKiNCFQsVFZURoYqFiorKiFDFQkVFZUSoYqGiojIiVLFQUVEZEapYqKiojAhRURRVMFRUVE6KoiiSqCiKmkBARUXlpCiKoqYlUlFRGRmqWKioqIwIVSxUVFRGhCoWKioqI0IVC5VRiSCodv1TRRWLj6CwpIyZtQspKR93ppty2pE0GqqnzTpt9Y2vnnLa6vo0kTQarrj+Zhacv4TZC84jMTnlA/tYbXbKKyecgdad/WjOdAPOVgqKSlmz8lWycvM/1fOIooQsxz7Vc/wrU2bMISbLp6UuQRBISc84LXWdKpIkEYuN/N4lpaSya9smGg4d/Mh9CopL6e5oPx3N+69jVPQsRFEkITHplI6JRaPo9Hq62ls/pVbFyR9TBIBOr/9Uz3MMQRAor5pIT2f8gTCZzf9WfYnJKbgHBoZfz5q/CKPJTM3009dzeT86vR5BEBAEgcSU1FM6trh0LO0tJ8/xmZqWwUBf74jqs5/id+o/nVEhFlqdDqs94ZSO2b19MxNqpg2/zszJA8BgNKHT6zEYTYiiiE5vwJaQCIBOpycjK2fE5xAEAXtiEoIgkJaRdUrt+6RUVU+hfv9eBvqcWG12liy7hoSkZExmCxqNhqzcfExmC/aj15SQeHSbVkvp2Eog/gudkZWDRqOloKiE5oZ6zBYrAJvWrcZssbBzy0bMFismiwVbQiIGg/G0XKPVlgCCgN5gxGY7tc80NT2T8dVTqZk+C0EQ0Wi05OQXMr56KqIkUTN9NonJKciyTMX4SSSnpJ20vsSkDw5j/psZFcMQrVZHcmoaOp0evcGA1+MmNDREJBwmGosCHH0dwmqzI4giXreL5NT4l2XuwguQ5Rgms4XSsZXEYlFEUaShvo6K8ZPIyS/gj7/5OecsvhhFUVi5/IURtctoMhGNRjGaTIytmsjipVdhtdkJ+H0EAj4sFhuDXg+O7k58Xi8et4tAwIfP6yUY8CMIIkkpKfEHx55AMBAAFPy+QQa9nng9fv/w+XR6PWazFY97AFEUESWJaDR+LdPmzEev11NYUsaurZuwJySyf/cOikrHYjKbCfh99Pc5kSSJq276Enu2b2FMSTk6vZ6ps+ZhMBhZ/tzTTJ+7gImTp/PSM09QNbEGUZLYvmk9M+edgyzLvPXqS+j1BvIKi/D7fcixGJJGgyzLaDQajCYzBqMRs9mCyWJlKBhAkiTC4TBDwQDpmdlsevcdLFYbN/zPHbgH+gmFhpBECZ3egG/QQzgUoruzA0d3J61NR3D19wHQ3dnOto3vDt+PwpIKps2u5bknH2PhBRezffN6ysaNp7i8AkVRKB1XxeZ338FqsyNKElqdDp1OjyzLWKw2UlLTaGk8fJq+pWc/o0IsFEUZFoqklFTSs7KJhMMM9DkJDQ3h8bgYCgQAmDxzLmtWvgqA3+fDbLEgx2J0trcgiiJZuXks/8fTVE6sISMrB0d3J37fIDn5hVisNvbt2g6A2WIlISkZq81OanoGGo2WhKRk9AYDWq2OWCxGZnYuzQ31hIaGaDh0gFWv/xNJklAUBQBJo8VitWGzJ2Cx2khMTmZMSRkGkwlREACBwUEPHtcAA/19+Lze+MMSDhMaCp4wns8rLOaCS6+grbmRwpJSklPT2LtzG4f272Ggz0lqWgZ7d27FaDLTfKSerNw8xlZOYNUby1l00VIO7d9LVm68d+Xzeti/ewd5BWNYcMHF/Ol3v2TGvHPILRhDwO8jJT0Dj6uf4vJxPPq7XzCmpByTycy+3TsACIWGaDxcR0Z2LoXFpRjNFixWK6HgEJFoBL9vkGAwQDgcRlFkREmDKIokJqeQk1+I2Wyhv9fBlvfWDAuzAgjH/h4dpuj1huHr1+p0RMLhE74X5ZUTWPX6P1FkGVlRsNrs7N+1jQk10xjo7+O91StRlLj42hISsdkS0Op0SJKELSGRzOxcBFFEOU32n7OdUSMWBpOJrRvWfey++vfZDoxGI5k5+XR1tFI2bgLvrlpx1OWm0Od0UD11Ji/+7XEmz5xDSlo6q1e8wkCfEwC/bxC/bxCAQ/v3fOi5Zsw7h97uLvRGI5FwCEVRiEajw9tjsRgDoaERj6FPRnJqGq+9+AydbS1YbXZKxo4jr2AMbUfH8PbERHp7ukjPzGbcxGrWr36L6XPnk51XgNPRTZ/TwbgJ1aRlZrNv13bGVk3k4J6dNBw6QDgcIhwaorxyAgG/j8b6gwwFg7Q2HSEWjZJfWMSqN5bj9RxfbUyWZbraW0/ZJqTV6ujp6kCSJOyJScPCCnGhgPjnrQDBwPFeVWFxKW3NjSfUFQz46enqICExGUdXJxdfcS1/ffhBEpNT2bD2baKR+FKKsVgMV3/fcA8F4oK06KKlo0YoACRBEO4BpDPdkE8TrU5LfmExzQ31H7tvNBqlctJk8gqL6Wxvoa25iamz5tFQf5DwUJC25kZMZjM9nR0EAwE62pqx2RPo6WxjwuTpRMLhEx6Kk1E2bjyN9QeJRaPDQ6NPg5rps+nr7aGjtXn4Gu0JSQSDAaomTaa18QgajRYFaDh0AKPJTGd7Czl5hSQlp7J1wzrmLVqMq7+PlLR00rNycPZ04/N68Lhd8TojEWz2BBzdXXi9bjwu13DvLRKJUDVpMgG/f1hAPylJKal0trciyzJOR8+I60vPzKascjx5BUXDHi6PayA+jAmHqJ42i66ONhoP12EyWygprzipMVQURYwmM709Xf/W9fynIAiCjCAIIeKi/F9bNBqNkpCUfMbb8a9FFMUz3oZTLTNrF578miSNAiiCKCrCp3B9JrPljN+D49cqnfE2fFZFEITwqPCGRKNR3AP9p3SM3W4nLy8Pq9X6KbUq3hX/LBABzWkKWBTFk39lJCneSf20uucBv+9TqfeTIJ9CjMd/A6NCLD4JycnJ1NbWcskll2AwGD7+AECj0ZCRkcH48eMpKipCp9N9yq0cGRoRFmSB9t/8tEVR/FjRjYRDw/+PpvH8aGBU2Cw+CVqtlmnTppGdnY3L5aK7u/uk+9vtdmbPns3SpUuZPHkysizj9XrxeDyfUYsh7g/4IDEF0oyQbYZ2/4fuMiIURaG35+T3QeW/E0EQ5FHhDfkkDAwM4HK5SE9Pp7i4mF27dn3osEEQBEpKSpg3bx7jx49Hp9PR09ODLMu43SMzdJ6APQ1xxhKUQ1tQWvZjtGjIG2tHK8t4XAZ6qi4nsu55cDtObMeYiUhaLdH6bQBkldqYuCgb0Wxhle8qdvd2cm3d/9JHDHsC2M2wfj8MhT+sER+PTgO1E6B2IogCOD3wzw3QeAr2PkEQ0OoMRKPhk3bpBQHe5/RQOUOoYvERRKNRVqxYgd/vJxQKYTAYCByNxTiGKIqUlpYyc+ZMNBoNfr+foaEhmpub2b59O16v99ROqtWjuemnSJKA/pJbWNj5I6bMiZCTJBOMWPlN790USQrC1GnMeOpGXmqScYdBKByP9q4nQJAQ7rmQwhwfN/5yCptebKHNfh55c+dAIIDolNmU8Tt63HGRiMbg1gdgd+PHN+0YGgmmlMGdV8K0sbBuDxzphPJcWPsbeH4d/PyZuHh8HIkp6VROqaWj5QjNdTtPcIOW58K150B1Ceh1sPkgPLYCWnpO7ZaqnD5GlVgIgkBSUhIajQaXy0U4fPKf1d7eXvbu3YvBYECr1X5gu9FoJDc3F1mWMRgMrFu3jv379+NwOD627g9DnHohmRkGvtJzG8GSG/ln1l1kPvE5Vtf303r+fSTn7OZrY//KdyofYdK4PL5W2cKvGhN47qZHiL72R4SUHBKXLOOqJXtY/fgR1r/Uhf5nC/lx4KdQYOEB4Ye0/OLvrNnhRFbg8+fByz+GL/wa1uz++PZZjfDLL8EFU+HhV+JC0+eJm8sBspLhjqWw8n647udQ13aSa5Ukpsy7kJp5S+hsqcfR3oh/MN4Tm1Qcr+O9ffDie9DVDxdNh/UPwtU/hff2n/KtVTkNjCqbhSRJFBUVsXTpUux2Oz6fD5/v5NZ1t9uN1+vF7/ef8MsH8Z6FRqPB6/Wyb98+du/ezcDAwCnNhBxGZ8B8/Xf4qvQHzDVp9LX18qZ7MRuffoOmfgO+S39I28++Tufq3SROmMBrAwm8+cZWCi+7CZPVSuTpH+MNhin+8hcx7n+NdY8dZNnVZcg1FzJ14z3sOBIhWjadw4cFhhoPEo1G2dkA+1vgL9+K/20aNkfEbR/vz/mQmwpPfgfy02HZj2H5JgiETryEwSCs2gkxGR7+GqzYCgMfEQYhiCJFFTWkZOTiGXBycOd6opEwqXb4xz3w6GvwzT/CziPQ0AVvbIXth+GWxfFzhKMfXq/Kp4MgCPKoEgtFUTAajdTU1FBSUsLEiRNpbW09qW1BURQikcgHhAKORlgODNDV1YXT6Twh+vLj0Gg0WK1WYrEYsiwjlUyisDSLEnkTTUN6nvjBTkIF02FwACExHSEpg9gbj9LhhB6/leLrL0O395+sqP4RNXuf5I95B3DlGtlXfAvKM7/n4ZsHCU1ZxvJ3w7z6+xXU73Qza0EaOcVXMy41gY6WBoaCfpq74w/ko9+IP4wdzg8mhkmywl/vgsEAXHc/tDtPfm27GiAYgt/cBhsPgsP14fe1v7cTd38v+7etw+XswqiLH+Pxw/f/ApF/0dxWB7y+BaIyqI6Wz5ZRJxYAXq+XUChETk4ORqMRk8mEw+H4yB6GIMTHz5fMlri0NoX54yPUlMgYddA9AJGo8qFC8lHo9XqKioq47LLLuO2223C5XHR1dRFNzqG8wIes9/LCr/bh90QQMscgmKyI5dNQmvehHNoKQMznIbjo61y+wM2W6Dns+909eHPtLLijHK83g9oJIsH6vdwbuYfA6heQOw5TYJT5fLqXotpllOaX0NvTTfPhAwC09kJDJzzyDdhxBDreF12ekQh//lbcxnHLgzrCYgIGo5VwOHhSq+Oeo3aQX34pbtP4MMPnUMBHd1sDg+4+Uuzwh9vj9pBbH/xom0dMFYozwqj0hsiyzJYtW2hra2P27NlEIhFycnLwer0nGDCtRjhvMkyvgKrKcWRPvI3k3OlEhry0N2zmas0QjqZ3eX3lu6zaKXO446PPKQgCdrudzMxMli5dymWXXcbEiRMRBIFAIMChQ/UMpVtQBhp56ZH9hALxn1S5cTeaK+9CtCZS2LMf65xFHNq3nUFnO74t63nunK9RIW4j64ZMqq4pwtRwkF8lfo/LQ09j7I0hlaYy0bGecybA9SWwYvthxKmbyUyegMiJvaAV20D5Azz1HXh3LyzfCGYDfGMZtPfCLQ9oyCqZyaRZ5+L3e9n05gs4Oho+8ppjMvzfK3CgJS427+yCXz8PRzqO2zgANJLCnCr4xRehow/OufPDeyIqZx5BEISQoihnR/TQZ4xGoyErKwtBEOjt7SUYDCIAc8fDrZelUDx2OoptBpljryCmaNFoNKSkpBAIBIhGIxALEnXv4OCaH/DaqoP8eSX4gieew2KxUFVVxfTp05k/fz61tbWYzWYEQaCvr4+f/OQnPP74X4kVV6Fr24Fn4H2GAFFCc+0PMBqM3JBlIC2zgO0b3uGtF/5EyJaK7qq7+FzlSuaWDTAteBhXXS8PvABvRxcRu/pH3NjwR27tfor9A/DUEXinE8bOqWbSlHPoOFjP4QN7GejvOyEqMi0BblgES2eDXgv/WAu/ewmQjMxdcgMzF11O0O9l5T/+yL4tq0Z0n7NT4K6r4Pwp0NwDPQPxnookQlFW3B7y6Ovwh+Xx4ctnjXB0+RxFUbssH4UgCJFRLRbHEAQBRVEQBVg2D667MI+cGfdjTB5PZmYOkiTR3d2NVqslNTUVn8+HzWbD4/EwMDCARR+h4d3vsnPzSn7xrELfUY+pJElUV1dTU1PD/Pnz0Wg0VFdX09PTw8svv8zq1as5dOgQfr+f4xOsP4goaTh/6TXUzL2Afbt2svrlxxl0H58BaTXF4x7cvvgvuk6nJ6ooCNEwogCR9z0DKQVWMidfgNzQiNPRjX9w8EMnY4lHzRaycvwelU2aw8xzryAWjfDa0w/Q33Py9HOCKJKQnA4KuPq6SU+Mezry0iDBEh/i1bXC1kPQ8xn2JiSNDrM1FZM1GXtSFiZbCoIi4Olvx9PfgcfVRSQc+PiKRhGqWPwL1y+CGy4pxVL+PawZk1EUhYKCAiRJorOzk1AoRCAQoKmpiUWLFmE0GvH5fIRCIXzeAbq2/YC6Hcu556/gGow/YBUVFeTn51NcXEwgECAYDLJnzx6am5sJBAIjsnfotZCSZGT61HKUiI/mxma6+6MMBuKxErICkaOjCqPZwsSpc8Geyu5VLxP0nRjrkZxjQimsYV5hOekpKax6Y/lJc1K+H63OQFZhOUGfl97OZj5K3I5hsSWx7EvfwWA08+Kff4Gz6yS+1M8ASaMjNbOI6vNKMFiSGXQWImoMSBoNIBAODOLubsLn7qWzZSeDbjWo4xiCIERGnYHzo5g3Hr731UuQs++gqHIBycnJaLVatFotjY2N6PV6srOzicViWCwWotEoCQkJ6HQ6DAYDeoOJxNz5SIEDZJqaWL8v/hAPDAzQ39/Prl272LFjB3v37sXhcBA5mivhoxCEeJRlbmr8r6M/yv5DDto6BojJMiJgMkCiNW6ALcmOCwdaOxdc+SUqJs8hEA7RefjEoAR7mgEhPY9EdGx+5y2WXXcz2ze+NyJ3rxyL4unvwT84sm6AKElMnreElKwx+DwDtDWMLEBCZzAydtJMEpLTGHT3fzJX9L9gNCcydvLFlE6Zw7iFbhJzHXidEtGQnWg0jCRpkIU+kvL6MZhsGLQ5eFydRCOfTtqA/zRGpTfkw0i0wH1fKSJh3J20OaJUVVWh1+sxGo3IsozL5SIxMRGLxUIsFiM5ORmDwYDuaNYkv99Pa2srObn5JOTUohl4EYdzkMauuIswGAwSCoWIxWIj6kmkJcS9AjZTPPbB4Y67CyHegxgMxGMavIF4D6arPx4clWKHNLtCQkoWSSlptHiCtO3ayPt7AJnFiZhK59G+ZRNCLEJD/UFqz72Qg3t3Ht1D4KPmmJwq0WiEYCCAzmCkqW4nfd0j61nkjSnnss9/neLKyQS8Tro7/70eicmSTNWMZSRmFiIrWroOa+g6LKKRSkHWICCgM/eQUtiFIhsom9tJ0CdDKAdXXzvKZ5x9/WxEFYujXHsOLF56C9bc85kyZSqhUAidTocgCLhcLjIyMgiFQgwMDDA4OIjFYkGSJDo6OrBareh0OiwWC1qtFkEy4HS6KDRtZOW2D8YKfByJlviYvsMJ9e0jO15WIBSJuxu7+qIcPngAybWF5kAUl2MAwsetrhXTKpk+cQnF+UU0HNhBS+NhFi6+mL07txK1piDOWoqQOxYl4IHA+4YwehNCRgHEohA50Qgr5JTHu0Khfxnna/X0Swaatr1Db9uRD85ClY45404UUL1eR2nFRCw2Gy31e+lqO3lG7pMhCCLjpi0ha2wx6WUNyHIPsVAuAmkga4Z7DpEhGOwPoyiNJOUo2DKC+AcUJCUHd1/bB9o42lDFgrh78Ds3JJE9+fvkFIyjra2NjRs3Ul5eDsRnn8qyjM/nQ6fTEY1GMZlMGI1GQqEQ+qOp6RVFIRwOYzKZiIgpeJufp881RMP74wskzcfOigpHBXoGBLwBsOugIhFyzfG/Oo3AoCGJWOhYvqKjaHRgT4FIGBQZa5qOivk2xkxJREzLJNDeRSD56VIAACAASURBVCgQRdKKZIzNJdk2FovJSm9nC47ONgb6ncxffCkHIwY0/Y0Ibftg7GzobkQjRzHpRIxzLsUgCSh544g52iAWH0YJOWVIlbPQ5peg6M0ovceNnkLZFLAlEzEnIg90xYXmKNryGtIuvpiEmmoinS1E/ccFLeDz0dlSz5H926nfv2s4vd0nwZqQwYyleeTXtGBN9WBLtWCywaAzEVGUkLQ6dEaFYOgNUgudGO0hfP0WAm6JmNJPLJBK0BdgKHiK83z+y1DFgniv4qILF2MuuAqj0YTb7SYvLw+TyYQgCEiSRENDA3l5eUQiEcxmM/398ZwOqampw5mnm5ubMZvN8eUBDBa8g34KjJt4a/tx4yOKfPLpkyYb0vX3Is24mEvzmvnOHSnMu66Iq+foWZwrcGDJwwQu/gaatFzEvWsIy8Tdq1+4H83V30csqWZS2gFuuK8aQVFo3dKBpayQy27NoGFHP2JOCYEI1K9di6vPQUt7K0NeFwN9TuYvvRpzmYdLL49Se3kGaRkmpiVn89OsIyycM4Hx4wp4UPM6U8syKBiTz0ylCZ1GhPmLWfq5GOfXuhCnXYSrvp2QwwkGM+aZF2Nt2slQfw+U1ICzDRQZKSOHGd++gmuXdFJeJZJz4QKK83w073ISDctgT2Ewo5S+lsNE/cc9NXoRZqSBJwyhEXo588ZMpuKcGBqjH6/DROfeqcgxA5EhY9xlqigE/O1EwkP4ndX0NEUwW4uIDpmxJJoIh5yEvHbc/aN74aFRKRb/Gsr8jWVQNvkqtIlTAejv78disWAymYazPtntdlwuFzabbXjIYTQaEUUxPs1aqyUpKQm9Xo9Wq8XhcNDnjjAlbS1PvzXEYPDE8+t0OoxGIzqdDq1WezRMXEBadieZ6RYuKT1E08xbcOxby6Z3utlJIptqv0xY1JL7j69wZM53+ZnxXTYc7iecPwHNZV8jcu+lmBdfy9R5et57cBV1rzRg0+bQeEBDZ0MHU76+lF6Pmd7V7+Htc9Ld1siQIkJKNlJiCgUXTOCWGhtT179K1eE2IqkCzTWLWflGA8+a5rF7+Uv8bZ+PXYc76ciZTpH7IDMungqXLuDGwy/R8Ld9uJxOMm76HM617xFJKmLa1HnMrp5GoK+TfskIRgt4+8j+3FVccH6ILX/ZxGs/38KRJjPZNXksWmpl5zv9UDkfXD2IRZNQetsQYxHGJcJDs+GcHHihGUIjGJ5ptAZyi6uw57hJykyhY9c0wkMGwgENinLUZS5HEcQIGSURDBYFo3EMovYgCdntePqc+D1BCOXh7DkyqufJj5oITpPJRG5uLunp6SQmJuJ0OmlsbKS3txebWcFoL8E1OIhGo8Fms5GamoooigSDQSKRCCaTid7eXkwmE2azedhIGYvFEEURv98fT4JrtwOg0+kIx3SYEgow6uPTOe12O1lZWRQWFjJ27FjKysqw2Wx0dnby0ksvsbfHgzillq/a7sGJxAuNl7H19x1xu4HWjT19ErdPeJrP3+FD6nibprLF/G3BYa4zz8K/dy1VVTHGlm9h+XvjMW/7DYtrc8mbfSuVmFl54BAxfzKV9h20Bo7PhhV9/dQkham9ZAxZYzZh6ZzNAy/08U4HuGI7ufwPY2hZcCWO9fuRu45myPKGEXbW0TzjZsZNG0/H7/7C4W0NfLEMrnJv5k+DtQQvm8DGujyGelrQlo+noHQ89a88jTDrcjRWK9MuyqT59X+y4dkOptVehqLRsfYNGfvFCUy542I2PbUXpXU/AgrZlVX8zLqZOZnwagvcuzPesxgJBqMNYwKEvFV014cIDw1hTPAS8svI0XSQRQSNg9yxh8gsDROLyDia6tizIou0wjBR/zhC3hii5EdAGOVWi1EyRd1sNlNdXc306dOJRqN4vV4SExPZsGEDkugmFvHTN9iHwWAgJycnnjna6WRoaIj09HQ8Hg/BYHA4Vb/mfYviHDN8HpsYBnFhSEpOQQjFA720Wi1z585l9uzZlJaWkpqaSmJiIunp6cNC09kQZLxhHW1dLv76QBOhm9oQkjJRAl5ISCcY0fPMt98i6b4JzDJs4XvKVaS74YILqlizezdLvjaOV/7vWQwXPc6KBy3scxTSZkolzZJAWdMh+l5ew/z/l8eRtU6a9zcwKVnhi+VQWx5m1eXpPPXLbWxNSWGLpoo+qxtD0E3T69tZekUfv3tgzQn30+A8wCVLxrL56Uc48sZeALY7IdOoMEu/g8zLl7JAbmDzP54g2DwZz0AvctCHRhSYdNM8ioQdPPTQQUTBQl5pFRZbIp1vL+fV1Rmcd106loeWMz0bbi45iGPipXRv2MuSFQEOueFUYiyj0RBBr0hCVjvRUDoanZ6gBzRaK7EYCCIg21HwMdgvY00xkF6kI7+6j32rshEwkJKdi6NhN8qol4pRMkVdEAQyMjLQaDRoNBoaGxvp6+ujvb2dS2dGSMioICl/IX6/n6SkJGRZRqfTkZycHJ8d2d9Peno6VqsVr9eLVqtFFEVkWSYQCDA0NERiYiJ6vZ66ujoyMjLweQewuJ/g0VcGcQ3G7RtFRUUEg8HhoYfH4+HAgQOsXbeOVhnSvet4+dFD+NxhhDETQKtHadmPWL0QISmLvueeZEiWMEwpod1yHkP7n2fTxG9x/cw9WOvryHTUYZsyh60bOvjTXw5jTsvH0dVK/YY3KS6uoqJiGhZrC18VWrmhFNb2CKyeNJZun8KrDx2iraWFC2/5Bn2WTK688noMUTvpFYM07e5lsD/uAZG0Ipd/uwrB72LVQ7tO6Jn7olB3pJvsOaV8KbCa64zdNLW0sKvViSAJLLwAFiySef6e9fQ0DBIJh4hFhpBlmcYd6zDXr+fCxQJfSXFzbUKA9Z0xfnvYzKv9CfR295zy4xqNhElKKUKJTSfkt1I0cyM9LfWEfTlotEYURUYQ9PS3JhAJ6YhGHSSk60nMUmjZHSMxdRKRUABPTzPOrtGz8tiHMWqGIX6/n3feeYeNGzciiiLhcJhgML5il2sQfM59mEuO34rW1lYOHDjABRdcwNDQ0HAv4lhdiqKQnJyMw+EgISGBxMRETCYTiqJgsVgQBIHIYCMeVw9D4eOT19rb24e9K4qiIMsyoVCIfpcL+1U3s+XtFvzueB9b3vwqmivvRN7wEuKYCcQ2LQfgvWebKKxOI6XCTfC2P2MxaCgM7+cG+340Vyj8qW4538u9m6qs23mnYDbVGx9iGoe5sGAaWc/eTdGt99HeK3D+E+8y6boKxtQuYPl3XkeOKXjcLiwJCRg760hbtJCstHQObm1i0S1lPHHXVrR6iSVfHUfu2AQe++pm5NgHH19lKIBn5cusWpCF8yWBu6oVLp9rY311OYU1qTz7w/Uc2exEFEAnyrjr3qPUvZn7SsOckw3rmzpZnZvHdQ85cYcB40HEaReBpx/6TtXIqODsPkxqXgXhyABafYSCiTLu7r242vPRavNBENAZUvH32THaexjo8hOLClhsM+LGT1cvXlc3o911CqOkZwHxNHlDQ0MEg8Gjy+LFP3xRgIrMLsK2CygYU4JGo8FsNmMymYYjBzMyMoYzZQ0MDKDVajGbzXR1dZGWlnbCKmYJCQl4vV52rriTfXWtLN94NCRblofnkrhcLtxuNx6PB5/PhyAoGEoqGNi8DSV2tKPt7kXIG4tm2bcQ88YSfe4XEAqgyHBgXTc1+c149cmc5/ojtf6NPLVe5ut/gNChwwwl5dJy1a8p6NrE11v/lwxtiO6uLv68ycHKQ7uY9vXbKJmbgzQulxeegb5IBorPBbJMSkkV/fu20NFUT78+gTVPvUjNBalULMgne+lFFORH+dt3N+Ns88fdwKl5CNklcVfq0TiLoDdC7Q3F9BiMbEtJJ/nqcaQGApy7agcLgv1cUwS3jIVvjIfrS6HSHmNPP9y9HZ7dMMiUa0poagzh7pdhyI/S341YNgU0WvD0cSpEIyGS0wox2fOJhDuomGelYLyAy9FPyJNPLBpBlDRImigZZT1o9CG8vTLuzhSUmMRgbwftTdtGfSSnIAjyqJ8botfGM0WZi25m/hW/JRaLodFocLvduFwuCgoK0Ol0RCIRPB4PiYmJw8MUWZZxOBzEYjFyc3NRFIVAIMDGd99gaNcN/P5lmXV7R9YObdkkIof3xN2rx5C0CIVV8Qe5p3n4bVEUjwZZKiAraDXxoKzjCGBJgIAXQY4d/00UJVBksopt3HL793hq3S6a1m8Cdx/CuJkISZnk6GSmJut54ak/I6TmgtGKfuAIZUtn4DGMoafBw9C6V0COIYyZgJCcjeLqQcwohLqNxPq7ETUC536xjOmXF+IeUHjz0Xoa1rWQqFEosUOmCXojGvqLZtOjTcXTfJho4/ElHsdePAnKplO/N4TibEfZtTp+rSY7BAfhFCMqC8vmkDt2BmklPiZe2IK3L8LuV8ehkfIIh/zIsRiiJGFL85FVuZkhbwLOFonu/Ul0NGynq3UEOQf/y1HnhhCfpamRoDKzleTSawkEjwda6fV6TCYTTqcTvV4/bLM4NjdEFMXhaE+DwUBPTw+7du2i/+DDDPY38ejr8fpHgtzfwwe6uooMA93gi2fyEmwppOaXMnX+hRjzSvHKIhG/l9ixHHMmG0JmEUJSJrh6hgOnAEjNQ5x+EUJ6Id6mdra+vZrP3XQHO9asQPG5obsZpauRUNshps2qZdfWTSiBQYTccqJuN70uE+7tu4gFAnF7StCPWDQRXf0mSlPshNsOES6fhdLXgRIK0bDby8YD2exuzqInmIZsScHf1Uq7Hw56RNpyZ+AcgsCBrVA4AbS6eMZyvQlXyaU4V69F2b0GIS0XQacHjzMeZvkJ3JcB/wBWSyo6i5eU/CDrn7JjNI1DEEQ0Wh2iqEEQRSJBA7a0Ppq2JODuEGmt205Ph5rwE0ZpnMWH0eKAeeOCZOWPwxNKJCEhge7ubkwmExaLhaGhISKRCAaDAYfDgcFgIBiMB08YDAasViu9vb3xFHsN72J2P8HDr8i0OD7mxKeIrmAcNYuuYPaU2aTbLDTW7SKQVhQXBkVBqJoLkgQKiJVz4hGT3j4w2xGnLEbZtoK8xARKF30O94CTAXTUji/nwK748gFEwyhyjNnzz2XL+rVxsRrsR6ycg2C2obTsB7cDQaNDrJqHvP9dqkqKuen/fZOCwiL2vPc2clE1isuBUDwJORAgvG0VSvshxLyxoDeBx4mQPw4hLR9l59sQ8qN0NyKOnQGSBrFyDkpPM0r91vj5+7sQCioRdIa4YHwCYtEwfq8TrZJDy07Q6UsRJQ2xaIiQ34MoaUABT3cLnfvDDHQMcHjvelzOltP0yf3nM2oMnB+Hfyie1Wnc1DdJr55CNBpFkqRhQTCbzfT19ZGUlER+fv5w5m6j0QhAIBDA7/fjd7dh6P1f1u+NsnFks75PiZglEWfjflxpKcRiMkFHO0q0DaGkBsXRgmC0IO98CwClvQ5xwgIwWhDsqSiHtyH6XUweX03x2HJSMr7M6i0bKUoVqZo0hX1HBSMWixGNRY8nggn6kLevjNsnjoZrK+2HUNoPAeBOshGOREnLzMUWC9IbGEScfC5Ky36U9vrhYZW8402EsmmIc64AQYy389hwIhZB3rYCoXJOfNhRv+X4RUdCKAc2IJ1/M7IgoLQe+ET3zuft5eDOlSQk5WBN8GI0JyBK2rjIihKRcBCfx4Grr5WA36VOHvsQVLE4ys4G+On/ruS3v64lJM7GYLAjyzJ+vx+tVovdbsfj8WC1Wmlvb8dkMg0HYQUCAXo7DzCw4y4O1Dv5v1c+nWA/GYG6bWtx1+9EUWIMelzxEwUGEcumIje9b2w95EfevgIhqwQlFkVpqyOmyHQ2HyKnoASpZT/CvrW86mjla9+7l7p9u4YTDkf+dRmDkzw47c0NvPLsX7HZE/B5XSid7Sg6wwmT1wCIRVEObkAx2SA8BNF/OUc4iHJU6D5AOEhszd8RZ1yK0tsWt1t8AqKRIfocDfQ5jqYDPBrNKyCoWbJGwKgehgiCQGJiIhD3lhxpj9BYt5HplVaMJhvOgSFEKZ7Twmg04vV6kSSJhIQE7HY7iqLg7O1hy1sPMnjgp+w+2M2vnz+eIt9ut5Ofn09OTg6pqamkp6cPR4AqinLKeRqEzDEo3Y0MOjsZdL9vzVHvQNwI2t91okopcnwY4jpuD+lua6Lp0G4a9+8g4OxCURRcA/1MmTWPI3Xx8fn46ikc2LNzRAv/yrJMd0cbLU2HGTraE3v/hLEPEAmdkoFSEo82PRxEcfUgZBcjDnSdZjFW3aIfx6gehhwL1MrKysLv93PkyBFisRgrNnro/Mr9fOvm1UyaNAF3sByyZ2FLyic1NZWBgYH4ZDJnNx2NWwkc+Q2x9h28sgmef/d9k8aIi8WMGTMoKSmhrKyMMWPGDGfX6u7u5plnnmH9+vV0dnYedeUKiNOXIM25HGnt3yjuXEXNRAOluQpmIcp2g4ZBOcyRVmgbjAdBASBH44bQo0hakbzKRDKLrQz5ojTt7EfxBZlTBcXZUY50tLGtHo7Nozy0fw8LL7yU8mk5VNQmUVippbqlmB1v1WEVFSqToCoJUo2QqAetCciCzEKImgys7U/nnXV+6rf2ndJDbE3WozdpcHUHiEWPH5iWAAur4zk7k2xw5yPxBYvsg92ck+HncKLI/n51mPBZM2pdp4mJieTn5w9n2G5oaDjhl14rwdRymFUJNeVGUvOmk5Q1CXtKEQgiA456dmz4J2+sa2HDAXB+yNIjVquV6upqFi1aREVFBaWlpWRkZJCQkDBs91i5ciW33norTqcTsXA8lm//lWubf8E7k7/FJbYnSdYcIhwBm1UiGkrjuvCLJLX46dkMLx2GF5thYw8ce9YyS2xc8s1K0gutNO7oIyVFS25FAvld9eT3NbO3CXLTRIqzFNbuUfjhX+PrgFTXjuP2X97EC089TmbiBKacl0T/ujUs23uQcCwezt0dgvnTYOJskIzQJ9p5O6GacF8EbZKOt9e4efbHu4hGPl4xpi3NZ8lXxzHQFSAalnny21sZdA5x9QK459p4wp9n18DbO6C5G+ZmwHcnwREPfGMTDKla8ZkiCEJkVPYs8vLyKCsrw2q10tTURGdn5weGBJEYbDgQL5nJISYVrSU9cQ2SFM9Utb8FDrae3DYxODjIxo0bOXToEMnJyRQVFVFdXc38+fPJzc0lOTkZr9dLamoqAZcT+zlLWcTzTF/YRnfTIzwycDNDd85HDslklOSQt9jC4IzJJB7ZSG11hN56uH8qDEbg57ugIzOZa38+mS0vt/LM3TuYXRTiqzdC8xYL23Mn87s1Mlte6WHitHlkpZmYm7WWVb90880ndEz8VhYtO33sf/IQCxYozMyYxKqp2XxnywCvv9qDTh9faCi1GH70AvgiImP/33iW/6WTLX9r4Loagdpv15ByfzWv3reLxv6PtgFULcjkgtvG8vT3ttO4o49zPl/KLb+fQfrmTZw3dog7HoJ3dsd7ablmeGQOLMyGB/bBIwdVoThTjLqehc1mY86cOWRkZBCNRlm/fj1NTU0fme7u2JKH0WiUlpaWD11J/VSQJAmTyURWVhbZ2dnodDp27txJX18fqd97iKtLXmXXm3VseKkD4Z5Xif39J6R6Hcy88DqavINUVryHxzFIpbOOS2fBZXdDbSr8z5Ikdlw+nbeeaGDd00f4zlUK1y+EXz0HT74FpgwL//PwTJb/opXZ87+J0WRizT//gs2/hjvvK2ZPfyKGNWaW2Lpp7HDwrP5ctrat5Yp7JvH41zby1Xleakria5i298G5t5RRPjOdR7+yETmixZ6SQWaCm6U/qKBWcvLKg4d5dDP4/8V8kZhp5Jbfz2Dj882s/0c80CzBCnf/pozk4iR++fnN1LUq2LRweSHcNRHqvBp+slfPnu4A8iieJn4mGXVBWYIgUFZWRlpaGtnZ2WzZsoXDhw+f1NBoMBioqalhzJgxdHR0MDR0POxXkqThSM6RciyjVn9/P83NzTQ1NcWzcCUnk3b++QysXs7G55uQIzJCSja6jAIKhAgzltxEVnIGa599lXNvy+f/HuhhTLqG685VeLzBhunmKejWNnBZeyO1ixQWToGbfgEvr4+vC+p3hwkMRjjn86W07zViMJiRu/aSITiRFo3nWu1eUpyt/Lqhkh+saKBo0izeWb6WvhYvt/92ElP1XVz+/Rg9Lqicl8HCm8t47t5dDHQOUTP3QibPW4Kjd4h3XthOxrJKbpgf4qakQerboPWo80KrF7nynkk423ys/GM9KPFlDJ64C7JlF7uNxRyuC1At+3l8PszJhG9sEnhLP4es6vMIDQVx9/ee9P6qfDqMOgOnIAh4PB4cDgcNDQ00NDR8bJZtrVZLWloawPBksmPYbDaKioowGAw0NDTgcDhOaSlDYFhoDGUVDNXvZPvypuMR3343cl4FXU0yTtGA5B2gIGci2fK5/PLJZWx+rY6U1A3c9YiVtX9vpHd9E1fdDpMD8NvHYM/h43Z+SYD2Ne2YryukSvcKCztjJBd1cuCCKlZvc3LT3z386dsK6UMKQ5EovkEPiVa4vryXikAz/zRNI2dGEwtnplE4IZkX799D6z4XOr2RrIJSMnLG4HJ2cnDHWp68exfGB6ZwyeIIb5T08sDf4cFdAhOvLSGt0Mof/2cDgqJw7uT48obr9sLdf5apnbuf275XycJn+vi/nTEer4fBmMDCaSXkl9cQkxXaG+uInczbovKpMap6FscybTudTnp6egiFPn75K6PRSG1tLYqi0N7ejst1PA2+JEkUFhayYMECcnNzh+eKnKpgAEjFE/Bs2Ux04H0uUVlGuuzrhMbOon7lUxx84fcUFo1h2/r1JFQfwROrRy5NxLmhiS/kNXPRNPjjSvjeX/5/e/cW2+ZZBnD8/34+xP7s+JiDEztO0jRJ16bptmxrt45O7ZjQBtoQF90FnSYx7YICRbsACQkk7nfFBTdjEhJCiEkgEKoEQoJN3Ua7tWvT09qmztFxjo4Tn882F+lh6Q51u7RJmud3Eyvf5+RNFD9+877v8zzwSie80Q/9Hni8CV7rhVe6oDCbxvxyDydH5zn7dC+XolV+/8szDE1WOHYOfv59B8/2xdi1w88vvnMVtx0O/2qR8FSZjl0eYlMZ/v7mBSYvLa/oVqpVcukUJpOB4QsfE52ZZHE6y/incYz7HyHtd7LrKRv9L/SwdcDLB2+eosmU5tevwo9fgr/+C95/D376ELzakOGit4E/J+y8fXRhuXRetUqpXMLucDMbDhEZG0K2Ou8/SSSrgcvl4tChQ/h8Pt555x3Onz+/4rrb7ebgwYMMDAxQLpd56623OHPmzB1/HxXcTjV86XMrptq+gwBUPvwblIs0t/hp7+rm2Ref470TbzM7lmDsbAyzYbnQzvUzHorlIr/f7YCgHeayy+0E/nAVHLtb2bm/hSsn5jj/7jS51M136t6eAE/1pmnr7ObimY/59ylWlAWEmx3crjMYTZjMdeSzmRWHm5xNFp54KUjLVgc+leSH7SM0GIvUKVBhmLoIxQQs5uEvI/CnECT0Ol77zZO8feQ4iej1H0Zh1esp5LOUS3dfvFfcPelIVoPGxkZef/11DAYDR48e/cJA0NzczKFDh9i7dy9KKY4cOUI4fG8KvCqlCLR34nC6eHT3U/zxd7+9q5nMl7HqNuqdTpLxONlMetW+rgKsdeDRoc0KVsBqhLMLMJ9dWYDX7qmjmC+Tv3V1VKyZTbfAeTe8Xi+9vb1omkYoFGJm5vMt7dLpNNFolMOHD9Pb20skEmFwcHBVX8SfVcjnmJ4MYzSa+Pb3XubyhXMUizUWpryNUrFIsVAgn8ve/uY7VCxDIgeTSRhNLp+ZSBTh1ho6hWyZclGOX68nknVaA6fTSVtbG0tLSwwODl5rYvx5yeTNfIXTp0/fdpfl67iewzEdCRMJT/CDH72Bw+VmNDS0KgHqXo1bbFyyZlGD64uYHo+Hc+fOrdg6vZXZbCYQCJDP54lEIvdtjEopHn5sDwdeeJGx0BD/+ec/WPrsQmmNPA1NtAbaWJifYzqyuftkiJVkzaJGSimUUl/7QNb9EOzs4pnnXsCq68xEJjl1/H1mpiZrGnv7lm4WY1GS8eWdjnv1b5TYeCRYPMCUUnR09fDonr00+Vool0osLkSZjoQZHwkRi86TzaRXBBFN09jx8ACjoSsM7Hmaj95/F7e3kVh0niZfC/OzMxTyeSxWK9lMGuO1LvO6zU50bpa2ji3MRCZXbf1ErB8SLDYRpRQWq47b24DNZke32zGb6yiVioyGhnA43UyMhnj48T2MDF3G29iM0+0mn8uhaRpW3UYyEaexuYVYdI65mWl8/gCBYCe5bIax4au4PV4uXzy3qrsoYn3YtIlkm1G1WiWbSX/pCzkQ7Lj2SNHoayE8OkJTSyuDJ0+w75vPc+r4MXq291PvcBKdm2HXY7s5/dGHtAaCzM/OYNV1LLougeIBJrshAgDdXo+/rZ2l2AK5bBaHy83C/BzpVJI6i5VKpYLT5WY0dAWlFKlEnPjSIpMTY5TLJSy6jY6uboaHLtVUNEdsLLIbIlaFwWBg56NPkMtmuHzh7O2fIDYcpVRRW+tBiI3PYtVxe7xMT06s9VDEPSQzCyHEbcnMQghRMwkWYl3wNjahrpXmv5WmGeh+aMcXXtv9jf3Y7PUAPL53H/Z6x4rrwc6tPPPc85jMXzx5bt+yFeO1Prbiq0mwEGtOt9l47Sc/w6rbbnyu3um68djl8ZCMxwFQ2so/WU3TaPG3oTSNbTt2USjcrFFiMBhxuT2MXL1yoxfKrc93ujyUvqIA0q33b2aydSrWXLFY5OypjyiVirg9DRiNRnTdRrFQoK2zi3qHi2q1SqlU4ukD3yI8NnLj5GmTrxWUwtvQRDqdYnJ8FN1mx+ly4w+209ziZ3josrrrQgAAAp5JREFUEp3dvVQrZfbs28/48FVaA0Hy+RyBji2USyXqHU5MZjMWixWn27P80eXmyX0HiEyM0eoPguLaIbQspWKROouFcmlzpNFL1qlYNwqFPMHOLloDQez1TsyWOnz+AOHRYfoeeQyjyUwqGadSqTA3MwWA0+3BYDBi1XXq6iwUcjli0Xn6B3bTs72PxYUog6dO0L2tD6tuY2F+jlQyga7b6B94AqPRSHOLH5PJjNWqMxWeoGNrDw6Xi9ZAO4V8nnRqOZu4Z3sf+VyO1rYgdRYLjb4WNM1AMhFfy1/bfaOUqsgcS6wbrf4g46Mhspk0xUIBg2Ygk06TSSVJJeJYrTZmp29m8waCHYTHhslls1w8+wko2LZzF5VKmZnIJNVqFbfHy9xMhFwui8/vZ3YqQqBjC7rNznQkzOT4KIV8nsVYlG19/WQzaUwmM4VigYXoHLGFeRp9LRw/9l98rX4uDn4CQM9DfcxsssxcmVmIdSOTTpHL5chlsyhYnuaXS8Si85SKRZKJJbyNzSwuRIHlYsepRJzo3CylUulGluz05ARmcx3+tnbS6RTxxRgOp4tYNIrD6cRitXL+zEly2QzNLQEuXxikfUs34yMh9uw7wOjVy5hMZmILURqbfMxNT5FMLFGpVLDa7GhKEQmP3VUZgI1KTnCKB1bP9p0MX/n0jgr59G7ficPl5uT/jt3DkW1Mcs5CPLDupvG02WIhlUzc/sZNSmmalqtUKnVrPRAhVpVSX91bUtwRTdPymlJq/Zd/EuJOSaBYVbIbIoSomQQLIURNJFgIIWoiwUIIURMJFkKImkiwEELURIKFEKImEiyEEDWRYCGEqIkECyFETSRYCCFqIsFCCFETCRZCiJoYlVIhg8Gwda0HIoRYv5RSw/8HvrA7rwnTVDMAAAAASUVORK5CYII="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydCbhNVRvHv0qj5nlQUsk8D6WSSlKSFBoMaaBBaaCohEioEIWIZMqsRJlnIvM8z1OJaKAI1bd+11natn3O2fuce91z7/2f51nPuffstdfwW2uvvff7rvd9//c/fURABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABERABDI6gZMyOgD1XwREQAREQAREQAREQAREIOUIZMp08skXXXLZ5f/++88/Bw8ePJByNalkERABERABERABERABERABERABERABERABERABERABERABEXAROPW0009v1u6Tz+ds2HVgwZbf/yUNmzJ/Ve2XGjY+I3PmMwVMBERABERABERABERABERABNwEThASERABERABERABERABERABEUhuAg2bf/DR/Q/XePLbof37bNuyacPFl15+RYlSpctefW32HDt/+vGHV5+pUXnxvNkzk7telScCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACSQROypQp0/QV23574922ndxISpUpV2H8/DU/zl7/818lS5e9V8hEQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREIEUIXHLZFVlQSOQvUryEVwWXXp7lyi8nzln+/Zqf/sxXqOgNKdIIFSoCIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACIiACJ598yimRKKDUGL9g7faRM5dtPOvsc84VMREQAREQAREQAREQAREQAREQAREQAREQAREQAREQAREQARFIFQI3lry9DMG4X2/RpmOqNECVioAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiIAIiAAEWnfq0X/exl8OEYxbRERABERABERABERABERABERABERABERABERABERABERABEQgVQhkz5U3P1YWjd/76NNUaYAqFQEREAEREAEREAEREAEREAEREAEREAERSBkC+AwnmGnKlK5Sk5PAGZkznxnNx3ty1qeyREAERCBRCXTtP3w8Abgzn3nmWcnRxixZs10bqZxEuldGa2ty8FAZiUvgnPPOvyBxW6eWiYAIiIAIiIAIiIAIiIAIiIAIiICDwMuN3nn/s6GjpwaB8kSdVxpOXbbllyDnZLS8LTp061OhSrXHU7vfH/ca8m3/UdPmp3Y70kv9V193fU6C90phl15G1LsfJ2XKlGnA6OkLSpe7v1L67mli9u7yLFddPeK7xeuuynZtdj8txHri/U96DTrl1NNOi5T/3kqP1MDK4r4qVWv6KTdSnnyFit5AWdfnzlcgXL5EuVf6aWu8PHR+4hLIU6BwMeZqqTLlKiRuK9UyERABERABERABETi+BE48vtWpNhEQAREQgSAEbipVuuyJJ5wYaK0ucuMtpfb+/vtvQerJSHkRst374MPV//770KHU7jeCqoMHDvyV2u1IL/XfeMttd16W5cqsp51xRub00if141gC2a69PmeOPPkLnnfBhReJz/EnUOymW283Ootr/jEfP7U/+Xy918uUf6BKoeIlbomUf+q4USMOHTp48NbSd5f3U26kPNwHOb7399/C3gsT5V7pp63x8tD5iUuA5wBad/DAX3oWSNxhUstEQAREQAREQASOM4FAQrDj3DZVJwIiIAIZmgDuKrJlz5Fr3eoVy4KAyFuwSPElC+bMCnJORsrLbkb6u2jurBmp2e+LLrnsctxALF04b3ZqtiM91V3QCEQPGg3Q1o0b1qWnfqkvRxNgnPllw5pVK8Tm+BMwOvSk94dfdu3c4af27Lny5CffxZdedkWk/Ht+/+3X5YsWzEUh4qfcSHnyGiHw7p937vhh6+aN4fIlyr3ST1vj5aHzE5cAFki0btmi+XMSt5VqmQiIgAiIgAiIgAgcXwKZjm91qk0EREAERMAvgWtz5MqTKdPJJwdRWOAHO0kIvmCuFBZhQOfOX7joL7t+3mnkWOv9jkVK5Ls+d94kVyXLlyyYlxLlZ8QyCxS+ocS6VSuWsUs7PfX/7HPOPY9d2EbHleXff//37/YftmyeOWXiWGOckyF35BYoXLzEv+azatnihelpnNNKX/7bCX7CCX7afO75F1xIvpOML69o+VcsXTg/f5HiJS6+9PIrdmz/YVu0/OGOH1ZGhL8PJtK9MlpbY2Wg89IGAdyWbduyacNvv/6yO220+OhW4iKuQNEbbsLizdyS9nMPXjBn5vS02Be1WQREQAREQAREIHEIRH1xSJymqiUiIAIikLEI5MidryA9Xrty+RK/PUfwQd4lC6WwCMcsT8HCxSIJsvyyjjdfzrwFClHGsoXaVRkvS86/4KJLLr30iixXzZgyfkxylJcIZaCwfPGNt1s9/PjTL5xyyqmnOtvUt1unD9s2f6NeIrTzeLeBHelbNq5fu9dsyT/edau+//3vQMiN3VnnnHPuH2YQojGxc9fPeG1cu3ol5WGNEavC4kJz8iWXXZFlSJ8eXcK1LVHulX7aGo2vjqddAieedNJJ2XPmzjfFuENLa73gntv4vY8+LVXmnvvcbX/5yUfunzJu5PC01ie1VwREQAREQAREIHEISGGROGOhloiACIjAUQRy5S9YhB/WrFzmW2GRv3DxG01ohkMrlixSIGeP+WQ8mZyYM0+BQr26dPggtadbrrwFCv+xd++eTevXrErttqSH+s2wFqUf6cWtBnO1zad9hyIMwsrq64F9P//RbMPNnPnMs9jJOu6brwanh3EL2gfT/bOzXnPd9aO/HtI/6LnKnzwEjNe1A5R0/gUXXbx929bNfkvdvm1L1Lx2l/lpp59xht9y3fnyFy52I79FUtwnyr3ST1tj5aDzEp/ANdflyHXqaaefvnzxgrmJ39r/Wnj+hRdd3Hv4hJlYV0yfOHbklPGjRvz2y+5dxhjw/NNPPyPz99MmjUtL/VFbRUAEREAEREAEEo+AFBaJNyZqkQiIgAgkEcidr1CRnT/9+MOvu3f97BcJO4+NbHPxX/v37fN7TkbKd+31ufIYOVjm5Yvnp7pwIGe+goVXLVu0wG/g2ow0TrH0NXf+wwqL9BIT5Mnn67+BsuLLfj27vfvGy89qnhyeFbnMdXOC+SxdOFexX2K5UJLhHGspgdDST3H//P3337jw2rA2esyRfX/++Qdl7jd/+CnbKw/3QepbtnBe2JgAiXKv9NPWWDnovMQnkDNfgcK0Mq0pLN79qHtfYwR1ZdN6zz0xfPAXPROftFooAiIgAiIgAiKQ1ggo6HZaGzG1VwREIEMQMK6+MxHjYOXSxQv8dhi3Gznz5i+0dKECbodjZgNuE9jVL9eUyMcuxCuuzJptWRrbVZkSLJKrzJx5CxY2ero/165avjS5ykytci69PMuVtV9u0Hj2d1Mmtnj9pWekrPhvJLBM4r/0ophKrTkWT73EAOJ81jE/5RBTBhdeWJRFy282mydZVljFRbT8XscLmBgYuJYK54Iqke6V0doaS/91TtohwMYUlGtGYZFmYlmVKf9AlRtL3l7m0w7vvyNlRdqZa2qpCIiACIiACKQ1AlJYpLURU3tFQAQyBAEsAXATsNIEIPXbYXbqnXzyKackQnwGv20+3vnYzYpf9F0/7/jpeNftrA/rCv5X/IrkGwWUdQQwZzd38pWaOiU9XuflhriEeqdB3doIs1KnFYlZaw4T+wUBeBBlbmL2JO226pfdhxUWmc88+2w/vTjhhBNPXLl0kS/l+xmZzzyTMv3Eu/Cqm5gAufMXLhrJHVSi3Cv9tNUPX+VJuwSMxViRTevXrvYTCyZRevn0yw2bbFy3ZlX3jz94N1HapHaIgAiIgAiIgAikPwJSWKS/MVWPREAE0gEBE287KX6F8Rjk2xLA+sJeumCeXKWEmQNYWMQa3+Pqa7PnKFm67L3JMb2spceyReFdliRHPSlVBtYh15hIodHKx1Lo9rLlK2IxEC1vPMfPPf+CCwmya1zApPm5j8uy8pWqPvbNkP69t27euD4eLunxXBRTa4zbuwN/7d+fyP1LzvUi0fr5q/FVj9VP5rPOiqqwgAOuo0x2X4rESy67PAsKKdwhxtLv63PlzY+VRqT7YKLcK/20NRYGOidtEEBhldMoYNNS3KXCxW8qeV2O3Hm7f/R+C+KlRSKdntfAtDHD1EoREAEREAERSNsEpLBI2+On1ouACKRTAjbgdpAXWawH2KW3cd3qlekUS1zdOuXU007LnjNPviBWK7ZChPMDx85Y9FHPwd9g/RJXQ8zJKKQIULl104Z1sZSV3QjlYjkvuc5p+fFnXwyZMGtp0w86dodruHKbtf3k83bd+31Vv0nLdslVt1c5BYrccBO/B1HwpWR74ikbBY/ZZH7WoN7dP4mnnPR47llnn3NuNhOk1qyLvhW5qcEhudeL1OhDpDqxYvpl184dflxC3XjrHXdRljH+O9VPPy674qqsxghuS6xu0LgPUk8k14iJcq/001bitTR5/+Nug8bNXIxS1smQ64FYAi+92fw9P2yVJ7EIEHA7SbkWYzyeytWffGbEd4vXlQhdY7Z3WOc9W++Nt3lewf1Zcva6fOVHH+PZZeyIrwZFKje118DUfkZKTuapXdaFF196md94RandVnf9XF9XZbs2e6K1S+0RAREQARHwR0AKC3+clEsEREAEjiuBXMYfP66Lft6x/Ue/FectWLQ4QUblQsabWC7jMosd/7FYWJx1zjnn4m4LNyVBxiTc2OUpUKRYrPEr7n3w4eoDRk9fkCnTySf7nRvJna9JvWcfJ4ZAxUcee6pTn6Gj2CnqVYd9yd2Qwkq0gsVuvJn6EyGYerysUVjgf3/FkoVpxqd5vH32e35+E5sAYVyiB6hN7vXCL5/jme/HbVs3n39B9KDbN99W5m7axbj5aR+xm2JV5FJ+3oJFimN9s9pY4YSrL1HulX7aisugBx6tWQtl+z0Vq1R19qlR6/Zdyj3wUDXWDD9slSexCPxnaTk/bHD4SC1+5a1322S56uprqtV6/mVnvgerPfH0M6+80RSL0LN9xpnxQwblWaky5SqM++arwQcPHjgQ6ZzUXAMT4RnJD8+0kIcx7zF09NRHHn/6hbTQXncbGzb/4KOmbTp9lhbbrjaLgAiIgAiY9wdBEAEREAERSCwCCHbYHRYkFsU5551/AW56FIg2/FgiHOKo8aXuOy6ILW3R3FkzKpQsmL3cjXmu/s34Q4lnxiDEv/SKLFfF6g7q3kqP1lhnpHG4TYmnHfGci8/txx8oc3P/Hl0+Klqi5G01n33pNa/y6teu+uADtxXJ2fmDFo3jqS/auYWKlbgF66J4BJ3R6jgex1H8mB3pZaZPGjfqeNSX1upgnEPXsK94CKnVv+RcL1KrD9Hq3b5ty+aLLr3s8kj5sL4qdlPJ28mD4CtamSiFr7k+Z+7lcVjQIAQmvkk4dzWJdK+M1lZ42dgGBDofM2LoQCfD00/PnJn/B/Xu1jkaWx1PPAJ5ChYuxjxdtWzJwlha9+cfe/Zg7TS4z9HWeGZTedK8mDTmm2HJscHCts24ryrM84uf+1NqroGJ8IwUy3gm4jn5Che78cqrr7ku1jmamn3CuogA8atjvL5Ss+2qWwREQAREQAREQAREQAQSkgAuTxZs+f3fx597uYHfBt502513c452WoYnhhujiQvX7/DLNKXyseuRsSpV5p77gtaBVcWsdTv3v/Fu205Bz02J/AjYcVUybt7qH8JZWaREvc4yeSmFyedfjp2e0nWldPn5jDubWOdGSrctEcr/bMioKfM2/nIoud2cJELf0lob6jV+t83QibOXRWq3vS/N3/zbPx9+1n9YtD7iH5/5X/qeCg9Gy+t1nPgvzI/X3n6vfbjzE+Ve6aettg9YWFxuttK7+0QZCBRjYaVzUp/AF99OmdNv5LSYLemYy1aJ6+wNykGsDpN7nXyizisNuZYznxk9dk1q0U20Z6TU4pBc9T798utNWJPPu+DCi5KrzONVTuEbbr6VtqO0OF51qh4REAEREIHkJSALi+TlqdJEQAREIG4CBJWlkCAWFnnyFy4a9Jy4GxqwAF6icckU6TSsRBDAGNfc5wUsPmr2pIDbMVhXUDBt8uuCiT5GEt4jlKbMWIKj44sXIUSiWNKwu3NQr26d8HGcJ3+hpDloP+zEvPq663OGGxiEbX7dxEQaXCxnYLJ21fKlUSdBgmcoetOtSbvRY3Fb5qdrzM1TjVNnP3kTLQ+777mGTRzytQcO/PVXcrYvlnUn0noQZL2ItR/R1tOUHusfjYWFO6aCuy8oZff9+ecfuDjzY2FR7OZSd0S7j9GvcGXlzFOgEGvvkgVzZoXjGvReGam+WMeO8/y01Zb/Vf9e3X/Yunmjuz7YLpk/5/t42pES5/q9V6ZE3eHKROCa3AL8eNpPW3B/tizG+BXUPWPy+NEL5sw8RlGPW9CFc77/LrnXSe5PWDFaq59I/U/uNdBaHuc2zxmRxjHWZ6REnLPxzK9o/Tn3/AsuxMUi1r6R6jH7p/Ky9mDhFa09sSqyot3LotUb7jjB4TkWa4yYWOvVeSIgAiIgAslHQAqL5GOpkkRABEQgWQgYs/tCBBxdsWTBPIR0T9V99c3PjA/Z5u269LzoEm8XHLgW+Mk4FQ9i/s8L/MuN3nmfXcvP1X+zWbjGFzMvqY1ate8SqXNnZM58ZjghEoFZCRo6fcUPv89Y9ePeWnVfa+Qui362+bTv0G9mLFnf++sJM8cvWLudnV3JAtQUYjYEnoNZ+8olCwO7gyL2BW16qGatOpHac33ufAW69h8+fvbanftnmn6G8/lL/Ioft27ZtOvnHT/Z8m698+7y+Nl9vkHjFgRSddaDgqNj76EjO3w+aETj9z76lGMVqlR7vE3XPkM+6NJ7cLN2n3weTyBw5hSBW8MpibD4wXoh3HFcP9CmS6+48qgX3ybvd+z++dAx08IpqQaN+37xCw2btrR9ve2ue+//pN/XY/uNnDrXa46Qj0CeMOj7zeTZpLL3VXq4QCh+xdqVy5ck13zxKoeX33c+7Nqr++CRk++8t2LlcHVVr/38K5VrPPVspLYQVJvj7ILl2mIcGc+HatR6DmFTg2bvdeB/mxq1/PATrhGvMnG7U/ulho2/mjxv5Xcrf9wzyASHf/H1t1sxbu78sOs26NtJ9nfmzfuf9Bo0cMx3CwmgbgUOXMv01bpRC9cX2w/ncQTGDd9p8zFz2vk7u+a5xh998tkXo40TwpQ6rzZqzrqHBU+d1956hzUOZcvalcuSbZyDrjv07Ynn670+du6qbVj1EFDePS7R1oviRij/VusOXZ1CN/qLr22YRwsQ6mc9ha/fsY42FuGOs4YxX9zrlTP/raXvKT9z6oSx+/fv33eSWQii1YV/fNzdEb/JnZfrr/MXw8bMWrNj36TFG392BxomP3OE70gKXb/3Sj/1xTPX/bTVzQAhJNdP1wEjJrRo/2nvSALCh2s+/Tw74p1l4GqyVcce/eo3adUOhXG08UAhxTwaM2fl1mnLt/7K2sF9Ody5d9x93wNcr3M27DqA9U00YWi0+iMdD8KCvIPHf7+kmlmbbZkIwGFEO6cu2/ILzyhOIS/XKZx5bmH9jaetXufmyJOvIPU5N6ZccOHFlxAsm7UYS8wgdbLe8ozwca8h3xLvxOvcoOv6vZUeqcGaZO9DRW646VbmnPPexL2rxtN16zvri7YG2rx+5xfziHnFvQ2rFOajk088z0h+5my8a3aQcXTn9cvInuenP9zDxs9b82OvYeNnjPp++SbuywSnpgzmCBZqnfp8OQqrOPp+2mmnn2HHvHXnzwe41xXOIxj7pMUbdto1ifsU97T+o6bNb99j4HCv5xE/97Igz1O0o+LDNZ7s1Per0dTJWsnzVP3GLdvSfp51Xm/RpiPvK/GMic4VAREQAREQAREQAREQgQxLoEu/r8fxcs1DdY8vx0zDpHn8/DU/8t1nxCTPnaO45OGlwy80BKW2TMolIQz2Op8XFwTm4cpGwTJ9xbbfvF6wL7708iuGT1u4Zsaq7XtxY4Tgf96mX/++LMuVWZ3l1aj9Qj3a0LbbF1+iPJmwYN1P/M8OML99ipSPl65YXY1ccNEll3IuL1/h6sA1AwJMXv7qNWnZ9qtJc1fMXP3TH15C/slG2PZe555JvsgR5iN4onxcLfD96cBvJjrrqVz9yWdQGDC+I6YvWoswqPfwid8TeJuXeF46c+TJXzBWTrgRo95KJlCnVxm8nHK8+C23lfY6funlWa7kOAG4nccRxPM7L6Xu8/iNYy++0aw1xxCw8z/jPmnRhp3MJ/cOQdo3e/3Pf8EA5R3fzCVYc25KukZBAUHd9lqhnV4saDMCrkju3HDvwlhzfdN/lAVc1z2/Gvcd5SM8Q3E3evaKLQhmRs5ctpGXby/LCJSOCHFoG4LFhx6rXQelD+WUrVD5EXcbmS/MHX5HOMyc/X7NT39SH22y1j/WNVUkhUWLDt36IDxy11Gg6A03Ub/TBRDtsuyiuWhgHFnP4IAijfnNOUMmzFrKN8KWWOe6+7wg6w5j277HgK/hxPWL4Ib2INRzlhttvbDjY69ZrgU7hykvkpslv+sp7fE71rGypP20FyG4VxkILTl+X5WqNZlzCJEi1YWVC/lxNeXOR5wc1lOuBY5zbYz4bvE6dz6E8ayvkerxc6/0W188c91PW539wIoNjs7riOsq3DoEL5QM9jjXMgpNe340t4Lce6cs3bwbN4oo0hH+cS/nfOa4u17WPI5xvXKvZG1JqWC3QVjQTpSAtA3hJ/+jrLDXL31iXnEcBQbHENhynfPsg2KcYzwzxXqteJ33yBPP1KVcK8ilfO599lmAexvzMFqdrEsoOJzzAsGs13lB13U2YCBw5rnNrr9cP/Di3kTiPsz9O8gaSN4g84v7H889zKsGzd7vMHfD7oPMZassjvUZye+cjWfNjjZ+kY4HYUQ5fvrDuszcxhUZGx0YX+bOky/Uf4MyUEby3sEzP/c7jrHWcq/nWYPnlVebtv7Q3W7GhjnL+WwOGjVr+WbqYSMF3+5nIj/3sqDPU7QJxSOKRhRpPItxP+Aapt3cE+mXFBbxzEqdKwIiIAIiIAIiIAIikKEJIAzlRZ+dbQgd7E5Sds7x8uAW4vPgnyTIc+2mDAcR4T3l8sKHFYBxjX0NL4DsHHcLn3hhQNkQblc0L/e8BPCiguDaWSfnIojlpQGlBsfY+Udb2QXmzMuL0LAp81dZKw1cCSHg8vLbHcvkICg09UZzYeJVthWuh9s1j6IHngiTsOSgDAQN1MduSWeZWa+57np+R1DK7wjeYUf72CmPUsIpxHC3BwECFgixMAh3Dsoj6nyzZTvPwK28/CUJZh98uLpXGezS5/hd9z34kPM4L7BYynidY5UkzG0rNEZxk+Qmyuxidyt6UFZQB9eFtdhgZzfl8zvCsZRy94GA3L6033LHXeXoJ/8jTLe7Em0frQAznBAX1igIEJK5uTA3KTeStZP7+mIuIJR0rgnMOQQEbmssgg0z1+oaqxaUAgiAEFrYa8zpoxqrLl70w7nswic0bUU44O4HQsGkOR7adYsbJ9YXrBHuqVilKm2Dnde8YJ1gvaFftj2sCQgOrUDOjxDP7/URZN1BSEMbUDhRPu2CEQI0Z32R1gvOYbxQxth5jGKHtZjrizWPOhD4uPsQZD0NMtZ+WbnzcY3SVhRfXmVgIUM8CaxHsOJj7YpUl12juT858zE/EZwzVlb5aYW97nWC64q5Eq4eP/fKIPXFM9ejtdXZB9YGqyzAeol7LYLGLyfOWe6lmOQ6YmzYcU857HpGgIhiDDddVhkajhPKI+YpQj6ncoJnBO7T7vOwjqM+nlnsmsG9jDGLdX6FOy8oC8rheYP2lXvgoWr8zxrL/7CkvTauCW0m1hXXtX3usjGnYo2rEq4fKKxgzJrAcxFrAJsQeJ7AWpP22Y0N4co4rEQdOJy8XF/cd+iTVTK5z4tnXWd9oh4sbqONabRnpiDzy5ZlrUup21rrebXD7zOS3zkbz5odjVOk40EYUY7f/nC/Yhzt8wHPXMwzt0UkZRIfhbxex9xtZ61AWcl4odBC+WbXcu5HTgtsv/eyeJ6nuL/OWrtjn5cCPJ5x0bkiIAIiIAIiIAIiIAIikGEJ8GDPCwLmywj2eAmxMOzuqbvvr/yoE5B9UXELerwgoghg9zovE3aHL4JyBEvU634pRxDK7+F2WiMA4LiXBQY7tjjmDHgXLsKh/OQAACAASURBVKgwSo1oAq14JkXrTj36szMwljJuLHl7GfqRK1/BIu7zEa4jZEAA6RTsIAR55pU3mrpdNWE2T1m8iD1Y9fHa/O1UhFihHQIUr7YiuIvmniuWPjInnK6CbBkoBRBs085wVgNWGORWpGExYAVm7jZhls/LJIJzhNmRXG4gwEEhwa4/d2wQzqNt1BVLv6Odw7VG+SijrLD0hpK338lvXJ8IY51lMOcRPIUT9CPgD8fyiBVQufsrRWsXxxG60QbmpzM/LLwsH3BjRd0oXb6duXQDebxcOlEWrnfCWVUxBuyaDLcuYHnBsSxZs11rrw8UI3Y3LHW7rYiok3Xo66kLVk9esmmXW9mC6y/KZK64lUR+WIXL43fd4XqFtXtXOsonLKqc5UdaL2BCP2DEOaXNWCetu6ExxxqB/wkW6m5zkPU0yFjHw4+5Hk6ZjXDcjjNKhGjXKMJt1mj3Nc5cpB4EeLat1urLOX9Zq2CHoiRcn/zcK/3WRx2xznU/bbV9YL6jnEDZyP3D/o7VXZLQ3cPyD2s3jlmrN4TYrPFsTuB83Ahyz/dy48hv3At4RnDe0xBsYsn1ylstPnDypS9ssuA+6HSPxpjHE1DaawxjYUE57CSHB1YMCPVZR1AU2v6jxOE4/WP9cbpUqmLc9Nl7djzXivtcrNrYuU+fWPe4XpwKOLsJIlKduJajbTwT2HsO1jD8xkYS97nxrOtcV5TLM2o0DpHWwKDzy1pq1X6xwVvR6uW4n2ekIHM2njXbT3u98gRlFKQ/KLiY/37aVvWp515izL0sqpzns7mA+yPPvFg2cA1FclPq914Wz/OUVfp5KXT99F15REAEREAEEoOAYlgkxjioFSIgAiKQRODakFumW80L9OA+3T+ZPPbbry2avXv3/M7f5us3Jy58YeOndfniBfMiYeSlpv1nA0x5J5zwbNX7y6xatngh+cuZXc8Iif4+dOjQrOmTJzjLKGCcFhNY2bgVP+bll3MQBJB/6BefJ8VWsB+Eu08+b4S3k8aNGvfNV4Pt7zlClhZrVhzth/73X3/Z7Y6BkJxTImfegoUXzZs9M5Yy8xUufuNf+/ftM20+hkGlqk88jeLnk7bvNt2186cj1gTEIOn6Yatm+GN31onC5tChgwd3/7xzB37ERwzu12tIn8+OxAexAh/3GFMGbi0QaKREkNWN69asyuYRILvUXeUqWNdM4eKnoHRg/m1Ys2qF7SvnIGgI19YiN95SaqGJfcFuP3x4t27yWt1wY4NyAy4fNG3wEnPRmW9P6FqYP+u7qbGMbaRzUFC9bSw6COb9fPUH7v7NzFHy31fpsNDQXG9zf9296yj3M1wvq5cvWcT4u8tG4IpAmvEfPviLnu7jNnbBmhVLj5ln7rzMuadeePVNrrvvp00aZ48zP5hjc2ZMPRKnwh6DuZnGf95U6s6yxhvVWfVqVX3gD7OouMtG8JXfjOmKpd7xXu4xSpyrr82eg356xQrImTd/oU3r164mOOuDxhqBWABN6z37+MGDBw5Ql9n4eLIXdxRiMOj+0fstdv7041HKxT17fkta82BOH5JrrP2uOy+/+c77BB3t0LLJkZgAKH9x0+Uer0jrhbU0mz5xzEjmNL61xwwfMmDCyK+T3PmFC5QadD31O9bxctz+w5bNl2fJerW7HAS+8Bn99ZD+HDNBevecEYrb4lUnCiEEyaNMfuc1juCTne7dOrz3zrYtmzbYc3OYOUYgWOf8zV2gcFGOL1s0/xg3Zfa8aPfKIPVRZqxz3U9bbZubtf3kc+ZNi9dfeuabIf178zvXiVUQfzd53DGutmgX+bj/ovB96LFaddq/27iBQbb+yDwzUlGvscDNFFZMrRu/Vtd5T0Ohypx1ry0o2c+/8KKL333j5WftNc7u5uty5s63ZmX0tSzIHIyFBeUTOJh7FGvWa2+3bv+7WczffvX5p/iN41mvyZ7Dcnmz7lPV1jji5Fxz/WFXmVs3HWaXHB94cT8gOPwLDZq+a8JIZan/dPVKtMuWf7KB7fUcYI8zTlgefjt0QJ+Wb77yHPccuN9T8aGq5CEgt7Ot8a7rzDnW5d9+2b0rGoNIa2DQ+fXbL4fvu37iofh9RgoyZ2Nds6MxinQ8KKMg/eGexzwJ9zznbFfegkWLJ8VbczzberUbBTtKllNPPfU0lOWNXqxV3f3sa88Lci+L53nKbrJaMn92kgtMfURABERABNImASks0ua4qdUiIALplEC27IcD5Rr53K8ftXo7yaes/Rh5z9n8bQWn9vfc+QsX3bxh3ZpIL7fkxQ0LLoneeql2DausQOlgfdciDHSXUcBYWCB8PPDX/v1u5LgIQHDJOdMmjPnWebySibvA7tfObVocCZyNcO8x4yYG4TLCJmf+WdMnjedlM1rA2ViGHUUN5S6cM3N6LOfDYJlhg6DZef7hgOj139yycf3aQb27e7pTcteXr1DxG1ctW7KQXZB7fv/11/eavHZUAOIrsh7eAct4us+1u64XzTsc5Do5P1s3rV/HLjr3jvu7TRwEBM/UFU5gcLOxBiEQspkGR/ylIzBjx/zi+ccqifAfzO47xoTAo81ee/4plGVe/Slc/KaSuKAYM3zogBVLFh0TMB0XL5w39/vpU5KTB4J/duAeOHDgrxcfr1Le9o0dytbCabZLuUf9CPrDCemefuX1JgikZ02bPB6Flbu9V5lrk+vM8o7UH9w+Idxq/+5brznzYf3BNb1g9rFzHUXGXrOwILz8sMVbr/3047atXnUg4MSFjJeCDkEHQXc5b9Swwf3c5zPm2a69PidCTVx0GRckjQb0/LSjFQByzVxo5plb6MW8q/H0C/VYFwb27NbJXW5KjbOfdQfBMDuze3Xp8MGff/yx17aNHb9GEP/75DH/KZU5Fm694Bjzne85M6ZNwrUUFjptmzc6ErDWeP5JClzv5hN0PfU71vFeM0Z+udUdj4gycf3FemkVMXAycyop0LzXh13s/I7w1Xn8sWdfehWlYP/Pu35sf0cRcuc991f6Zki/JOG9/eTOXyiksFgQ1mVetHtlkPpineu0109byffYMy++igu6vt06ffhV/17dbV+5ZyOAZt2c57H25cidvyBKaATMrBXcc77s1/OI+zbWcgSXVmBvy+X6rP1yg8YzpkwYgyLNyRerP4Tii4yi2f7OPf2hmrXrcP93Bo+uUKXa41yzVsES7zyLhwXnXpsjVx7uqQjSuZ+gvHFeYyj4yDeod7fObkF/sZtK3o6iJ5rQNkgfbaygP43CGLecnd5/5631a1Yut2Xg8ou1dvOGtcc8B5CHNalBs/eSlP1OxQvXnbVEct+f4lnXqfOqbNmvX7d65VEbMML1OdIzU5D5RfncE7gn3nx7mXu8LIKcbfDzjBR0zsa6ZgeZD868KX0Ncs+jPj9B3QubIOt+njeZzyiasQDjmkdRGq7/Qe5l8TxPMRd+3rHd3KGOfteIdVx0ngiIgAiIgAiIgAiIgAhkeALWT7pXYNmXG73zPubZ7M5zgsLfMn6XI8GzfvfdLk2sCxLK9Qqkhy9aLz/KCF5x7cJ5mIC768bPNYEa7e+4PSAGB649nO4W7HHreiol/M1aFz6xBPDmBRkXAzY4tLOf1k2N9dUfbfLyoowpPq48MJ+3bmCc5+GmZ+zcVdu8yiLeRbhgz9HqjnbcupHAKsLmxcyf9hKIFBN/L/ceBAxlDriDbuJKAJcjXsEN7VhzHtYTkdpmY3qwA9srH4FAaWM410bR+h3uOPE83O7MyIsrFX4nOd21cQzf9/xuha/OslHsWbdr8PSqF1cNXm483HmpB/cwXq5vaB9zy+22A+Em7ousq5BIgh+EjeSzwWCd9Vs3Zhz3cvmAIJZjrCsEQsVVmtPNSbj5YmMS4GPdiw3zhHIRWsU6pl7n+Vl3cLuC+zIUn7YMXF/Qnvsfqv6Es9xI6wX5Puo5+BvWTYSRxBRwx7hhrWX8EIY7yw2yngYZ63hZvt22cw/3ugADGyjels/66QwA7awXpQ0u35z3C44j8GaeO9cWhLHwIzA5Loqc5bBWhFs7bb5I98qg9cU612mLn7ZynXPN4g7K6WoJFzWsecw/3DC5xxD+3GdZC1DuMJ/ccV+4j7h5U451WejlXhIXRu71ybrMu6lU6bK2HSg2GE/uV/HOL3t+rCw4n2cV3BrSHlxdwczpso9nEzgzP90xUWzME1gmV18oh/st48KzAL7/3W7QbNwM1lt3vawdjAPu7KyLL/JQho1zQtnO9Yrj8azrnE99Xu7HvOZfuGemoPPLlm1dCEWLpeDnGSnonI11zY51vgRlFLQ/zHfuy9FiodnnGaw9ovUFV2OsR9wno8WJ83svi/d5intQuODz0fqj4yIgAiIgAolDQBYWiTMWaokIiIAI/A/BJrsYhw/64piXfawjdv284yfn7mwe6hFOLl88P+yuUoTG9Zu0bMeOS+duXoRiz9Vr1My6WHG7gOE8dmKuXbViqXto7n+4+hM2WK97BxY7bmnrt18OTAqsi/Bj4JgZC9mpWL921Qed7hZsuYuNu6b5s2dMe9C4WHILDeKdFpiG46pipccO/WhlZzXjQXucu0rtORUeqva42YD/14gh/XpFK4fjKAMQNrBrbM53Uyba3cf2XIQoZnN6ntXLl3oGKmWX94IYrUSitW/b5sPuVrJkveZam7fsfQ8+/LfZNjdq2KB+7E41mz6zust5oOrhAMR2rO1xBMGrjWsj5450e8wqrNgd3LNz+/fCtY35efNtZe5md6UXf1wLsGt0pTF/8XJtFK3P4Y7jCqpStSeT3K843Znh2qj8g4/UsNfLyqVHW3ywi5cy1xkXUu6yEXBboVS4HYtcM063WuHa9/DjTz//t4E3sNfRVj0IKrF2wSLKvUOfIM4ozCizR8e2rdw7q5110Q+ul81mwXD+juCvVt3XGvEbFifOHcE2n42Ls2LxwnnVaj3/Ss9P2r/vdHNiGa03i4qzbOKg0KZvvxzgGYyb4J/s4IzVSiocSz/rTolSpe+aOn70N/QZjvjmR9HQ+YMWjb8e1PcoQWak9YI2sFt32cJ5c+4q/8BDRm50Rp9PPz4q/gV82BHqtGgLup4GGetYrxF73o7tP2yzViH2t2JmvafNznVxt7lvGaOdc9yKGM5BuYk1zheffXJU8PIbSt52J2siawvrJu5vBo6dkeTGsE61B8ru+/PPP5ztz52vUBGsBMP1Kdq9Mmh9sc512hetreRp0Pz9DqwZb9R9qqp1tcTvdRs2bck3v61wrUH8jkKDe/eyhfPn1Kj9Qj1cxs2dOW2y5cLzApse3Ncgxx994tm6uDibbe5PTo4oPlAWuddhrg2eSb6fPnk8AnLiubAxYc53Uyc2b1D3GGF7rPMtVhbUh0sn1i7cOqK4MVafjZ0u+24vW74ia+OQvj26Otcqzi1drkJSPKGp40YlBS9Prk++gkVvYL1DEf+ecb3ldnWIezTqwoWVu85Hn3imLvdQXCRaF1/kwT0l1z73J9ynOS0eOR7Pum6tL9c73D6GYxFpDQw6v2wduM3ESuuJOvVejzQGfp6Rgs7ZWNbseOZJUEZB+8P8GNCza0eec9jME66tsOTYAvNcHq0/5jEsH3lGmGemcJabHA9yL4vneQpFI3XxThGt7TouAiIgAiKQ2ASksEjs8VHrREAEMhgBBAMIAr3cD/CC4RZmm9+SdsR7ucux6HDhwgM8bhCcgjBcsPBQP2Xct8PJu3bl8iVO3AiDEYJuMm+pzt95+WfHm3Vds3j+nKN8xFqz/H1GWv3Z0NFTuw4YMQFhQbV7byvm9LfvHtoubVs2Zad8uB3osU4FhBTGlfYClAtBy8hfqNiNnOMWMuMyp/gtpUojmHHHMQhXB0KKpGOGaZtmb7zizoeLJAQnXkIKhEwIIxbN+T5FgkvbsaQO267ylas+NmnMN8MQ4mwyyi7aQL/tcXY4V3y4xpO4/3H7K85vXF+ZGBWebUXwTxnEZ9n+w9Yt4XgVLl6iJLsBnUoDZ97it9xWmvnp5f4o6Djb/JT3ZssPO5upsr9Dq6ZHCUfqN23VDiHh99MmjsMNmrvt1uJgo+t64Zo2Fk4PwxhhAYocd/sQTJpQANe4rzWvfpStUOkRXLC41wjja7swgiUvhYhljnBx3LfDjrGIctZDP7Zu3LDO7aYLBd35F154MW4WiF3hpfS43gjauNYRmqJQGvB5lyOufKiDNYVv5zrGGBcqXuKWpca9yfZtWze7+3zBhRdfggAPbsmpmLL1RFp3cM2CoBsl0Dsfdu01zAQbZ2c98T+6mVgb7raGWy/IBw/W4VXLlyw0Vln1UOY4+4NQnjXAff0HXU+DjHWs14k9D+U5FhIoHOxvlas98QzzbMrYkUn3FT47t29Pikly0cWXXOask/XkkcefeQHFx/iRw4Y4j9FvysG9HEGJsXQx7nrGPHr3LYXdQjHYci+LdB+Mdq8MUh/tjGWu23kQra233HFXuVJlylXAPdrGtatXWi4IEbGWhBVWF7jic48h7eI3GJWv9EiNTxxuGfndrlPuecbaz9z+akDvz9xllryj7L385l5bYLZ0wbzZuEczFkObEKZ3/bB1sxefeOg+twvFWOdaPCyokw0CfBM3hPgmKB+dbbmvSrWa/O90uWWPlyn/QBWemWZMGT8m1va7z+Mek6dgkWIo48Z/O2yIl1DVLMH5UaoQP8l5Puv7s2aTCfPcGQcJZeBz9d9shrLpBxNsw2texLOuo0ynHX7uT+HWwFjml+07zyBfdO/UnvmP8tprLPw+IwWZs7Gu2bHOlVgYBemPbVefrh+3RQH0ZJ1XwiqAcJ/Gc457Drr7BqMLL740aV0faNw/Rup7kHtZPM9TxFVLWq/mpszzcqzjq/NEQAREQASCE5DCIjgznSECIiACKUIAAcRlZhuj1y5rXmQwtV5qgjQ6K2f3F4JDs9v7GNcQ5MOtDz6S2Zk/Zdx/AiQEcQTF5ncj19hMGVhgOMu+4sqrs/G/O55CxUdqPHmuKZhgn16WCwWLHt6ZhRsFBHRN6z33xCP3lCwcLgifrRPBN0GaH37i6RfCBZ8NCp5yaE+sgarZAQkXt1LC+PYteTgewWF/wH4+eY2fX/Lhp93LyuT63PkKcNzIKI7ZVWmFLgtT6AVs6+YNSQFFrcICwXKeAoWLWUsfu5veGWMEVwHsqmXHvrP/vLwikFsYRrlCMFbyewWedpZjecwLE1C7zL0Vq5A/OZngigOLnL7dO36IYN62h124BOTt061jO/rndY2yAxkhgDs+xbOvvN6Und8oOLCEcu+mpQ7OZT4hGI80l9hZyzqAssed754HDgdb9bJGuc6cx7GRZrd6uHghtjza4rauYG3CumJI38+7IhgKF8jy+tx5Cxh9zXLWHFi5LWywIGLNcPJjrtH3cOOM6zSEfOEUYH6uvUh5Iq07BUJrGa6qbit77/2fdWzTsvzN+a9FkedVZrj1grx2PiOkRwkysNenR8XquMqY18HZLUgOup4GGet42VlLnotN0GDKYm7efnf5isMH9v3cKbBGiJo0z686fE+xH+IfsIZgaeKel/QbZVWLDt36IHyvVaXcbQ2eq/mQexc8ZVlrh5VhAsUfzhP5XhmkvsPjGXyu+21rnVffao6wsPvHH7xrWaHUbNDs/Q5JMaMmjh3J717rEO3iGMJdc7uY4owtwe//KSyOvs9Yd2uea0sokLNzbUF4jkuiUmXuua/2i6+9NdkoqB4oVSTnp+1bN/da42Kda/GwoM78RvPNNwpdgrc728Fz0A233HYnMb3czzk8uzAniOfhtuaJtS+cd7VZBFEwMN8/fq+Zpwu86405Ju2x1ny2vprPvvgqmzo6tGrS0Kkwfq5+o2Y8631iNn1Qfrj7U6zr+n8Ki8j3J9oZbg0MOr/cjPsZCyzGobrZaOPF388zUtA5G+uaHev8CMooaH9su7C+GdSrW2c2fVhrHneb4YkFYiRrTM6x95sVSxbO83qudZYb5F4Wz/MUbWeueD1Lxzo2Ok8EREAERCB1CEhhkTrcVasIiIAIHEPgksuvuJJdd2ZT6RFBqc1kA+R9bwL2Ok+83gTXxPwfQakXUoTK7Nrv1v6/F3WEf2+36dTj5FNOPgV3BOZFvhC7tdkZ7SzDyGWTAhr/uG3LkV3PuPSo/VKDxuyc5mWfYJ5uywWEVgj4X326eqX7SxbMjmDarwADISdCKj8BAf1MIV5c2MHttgLxcy55cG3kJRBHmM/xuWZA/JZlFBbF4fCpS2hiz89udlXyt5fQjR1jCHrh7be+IPl2mNCElG9k1UkuoYhBgMDeWsT8p7C4LjvHcTlCQFheUt1WMzbeRLjdbQgBeGGeMXlCxF2r2YxlAi/LXgJ45kipu8pVoC2R3KEFYUBe4pEgJOrd5aM29lx2kDdq3b4L7jd6fdLhA9wfcM25y77ICLic1wrHEQbcdV+lh9nljFA13Dy0iiC30tBdh43DMs/oH53HEGaWvqfCg/zmpZyzgUNN8PKB0Zgc7sfRlg6Vqj/xDIqKaRPHfItQPVw/EF4Y3cMpufIXKjLIJZCnXtw8rFu1YpnTxQ3jzLFw7p4erFozybVMco6zm0G4deeSkCC+3TuNXi1bLEeWzm3ebRJuraXMcOsFx6yi7hYThwP3R24hqHWB4bYSCLqeBhnraHMh2nGrsLgotMP20SefffHEE048cegXn3/qPNcq4q7JniPJwoYP63J14zaMdWZwnx5d3HXRb3bE17jv9hueqnT3rV7Bpe05OXIfDmYeaX2Mdq8MUt/h8Qw+1zkvWlsJAI01JQJFp2u3p8wGA37/qNXbb3DvpSyvdYh2cf/FuuKzj/5TeFhW1+bImcdrk0OBIjeU+HHrlk0k51ig4Lj2+hy5KXPLxvVr7TF7baCAL39L/mvfeql2DaeLomhzx8/xeFlQh91tzT3sGOuKylVr8sw1YeTwoe72lClfsQrPSuNHfn3MMT9tD5cnb6EixTn27VcD+zp52vxYK6EgcLsc5J6Lq0KEyM6NEuxaJwbQ2BFfDtq9a+cO+hP+/hTbus79ifUKS6hofQ+3BgadX+56jJHF7hFDvuhFHAuUM+7jfp6Rgs7ZWNfsaIzCHQ/KKGh/nPX269HlI55HsZJ1t4fnfBSfSxfOnR2tL0HuN0HuZfE8TzEXVixZMM/ve0e0Puq4CIiACIhA6hGQwiL12KtmERABETiKgJEHXsgPvxjBgBvNfebFmp3bbuG5EX4U8DL/t+cTwI+XV6dQmZdbfNd2aNmkITsLEcD+sGXzRned5xv/HewCdApNqtd+/hWzQ/is3mZHbA6jLPF64TYW4hcguJgwaviXTl/RfoZ78phvv2YHabTgin7KIk+J2w4HA108f9aRAOB+z2UXJLu/vdwwXZXtsODexn6IViY+w5MChxp/4tb9kvuc7Mb3CTvS3Ts9yYebDwS9sbi1itY2jjNOuAFCMIHw+94HH67+jRFE2Rc+6iYfMVb4rvnsS6/Rp47vN3/LXX4Bo+TBmsDL3RMMiAmCS6NoLkNQFDD3mA/uOh558pm6CHY45haw+emvVx6sQhCQjf3my0FO/9+4osHtwRvPP/Go0ZNcigLwhy2Hd4w7PxeY62XXjp+2O3975a0WH6BwYUzZSe51vZAfAdVhK6f/3L94tRFhJG6EiHPgPI6ygjHkmFdsiZx5ChRilzoC4Eh86Bs7eJ39wCLg6ZcaNu7Xo3MHo8NMEpR69YMdyYwtViCHfY7v3eOsCysKL0Ec40w+swk/ycrH+WGdsrvnw8V2iXW8neeFW3dYy8g3qHf3zl7xWJxlRFovyGdjtxAnZqDxIe5ut9357hZUBl1P/Y51cnCz9yruFcwb4kwg4HULTLGKQCl+bcgdHHVXfarOS6whPTq1a+1WlnNt43IO6xfcj0Vrq1WCRnIxF+leGbS+WOc6/YjWVpTF5HMqfVBUPP1KwyZYPwzu0/0T7tmsF15rH/OMa4p7upe7IebZNnN/dq+rCGe93NU9VLNWnZ1mE4XbUsNeG6O+Htzfy5VbtDHzczxeFqzb1jqg76cd27l3i99rlDq0gzXf3Z47y1WszD0q2eNXhCwtWSO9GKBQ4h5sNgPMdx6/w6zxKC2GfNGjq/2de0rzD7v0/OmHbVtavP7SM3aNcd+f4lnXqSspvpKJOxRtt32kNTDo/PJiQ1wp7iPOIO82n59npKBzNtY128/c9soTlFHQ/jjrtBtSvJ61jWI5F5yXm1hU0frC/YY8E0eP+Cpa3iD3sniepxg3P22P1l4dFwEREAERSH0CUlik/hioBSIgAiKQRMAGxd1vJGNOJLh2wArCBKQ9IkDmuA2KbYXJbozZrsuRC5cNCOPsi2axm269vX7jlm0RGH/RvXN7ysCs3EvQwzGzqW6vLRdXOLiR6m52beLXmYDcXgH2zjZvJbEK1tl5vXzR/LnWzDzeqVHi1tJ38WIWi1A7nxEssFtx4bxZM9ztYIcfffRyT+LVZtwM8Xs4VzIc44Ub5ZOXUADFCa524uUR6fwNRlh+kdmyRwBkvp0BhRFAIrA1Uyovu+RqPP1iffpifMqPdpdpdgneFC6wNPOY/N9NGjsqWl/OMJLyn42Q050PxUL1Wi8kxQBhrkQrx+/xW24vW44dtZNG/+fup7YR1KMM6Phe80YITq0lhNloekzsDff1gpUQbqTatWj0ajYjAKAd4QJScq1yLFqMBlzG7TD5nH3C4uEZ43Zqu7GEWrZo3hy3khAlAsy8xsrNhj7w259/7j1y3T/9csPG//z7zz8mQPr7BLA93I8fjmoDv9ndqAj5+n/e9ajYFRyHHUIQt0/sMzKfdRbH3WNNTIf6jd9NCkrNehNunfM7vpHyhVt3WMs476CP+DeR1ovDfA675Ro+uG9Pr3UDd1kIkd1zJMh6GmSsk4ObMUZKuldh8fSgCfqLwJLYHF5lE0eIHRH3pgAAIABJREFUWCUco52PP/dyAxRvQ42bMXf+INw5l3m5fvXKsOtjtHtl0Ppinet+2krMBjYSWKUk9+cPP+s/zFhebn+7fp2k3dAozH/Z9fNO930WqxXjdusa8mA15DUOKCy8/NJfdsVVWXcYzYPzHOLv4J6IcXUrLP5jdiBwbCi/cy8eFtSBG0bWdNbV0cOHDnDWyz0VQTxubNyu+Li/YylAfCR38Gq/bQ+XL2/BosVtHCCvPGxc4HfiUTiPE0eEtd3GhkGp8d4nvQaiRH79hScepZ3h7k/xrOu0gfuTl5spd/sjrYFB55cXGxTurNVez4d+npGCztlY1+xY50hQRkH7424XbjuJN2XfPexxawnntfnBXQYxhtjAEG4zhjN/kHtZrM9TKJNZr/y0PdZx0nkiIAIiIALHj4AUFsePtWoSAREQgYgE7I5H98vDCw2avMtL2oDPj96Ve7ERHFPgpg3efoVzFyhUlONW0ICg4oOufYYYtzWbGr/89GMcu8RIMvn22sWOWbhz5+vrLdp03G2kJig6bHwLLwGs0XHsOc1ITvwMN21iF6Qzr/EocqKReR70c36kPAjR2Jk6a/qUCbGURdBBG3Daff4JJnQ2wleEqs5jSTEzjILJnd8qLL6fOnGcV1t4wUKoHC7AIcecQZbZ9W79K8fSN69z7Avei6+/3YrYJs5gryhRiEFCQN/6TVq2O9H4fWnz9uvHBA5HeJ4zX4HCuK3wqsO6D5gzY9qkaO0m8PVpZpu1O98bLdod8f1vQj6siFaO3+Pu6+WeilWqEsgUS6HeXQ+7iPrvevntGKuPw9fL/iS3auw2f71F247EjMBFE/6Y+R3XW17tYUfj5ijxK2y5bssUfHrPN3E+ENgsnn+YO8IsW4+1UGC3ejQWp5o+kMf2AwVTtafqvNyxdbM3cYVEP3DN4d4Rzzk22DMKH2f8D1undXnkFiyjjCCPkbUeNdbUi8CIusyG8LXRLHKi9c153O+6w1rGeQZL1PUs4nphhKbWgmJQr+6dvdoKHy+he5D1NMhYB+EVLu+hAwcOcIxg7NVq1Xl59vTJE3AT55Uf4RhzFGXoE8/Xe53d4R+2eOs1L+X2n3/sCXH3dx/BnWK4+yBtiXavDFpfrHM9aQ2J0FZcPXHfsvds1vkOnw8cjvVlg2cfq8K1l1SGEVJ73bPhe9it5PYfvZTjCOJJXvMMAeGhg4eOuu++1rT1h7OmTxrPPdq9tgS5NmKZa/GyoM4ixl0S35ONct29ZhF7g2Pjv/36qGDv/HbTbXfeDUc/St4gfcOSB9ePs4xrz3DWCjamgDFoOCrgNkHDsdTjmQQlzBvvtOlY4tY77mr7zpv17f2WeUF73HMjnnWdZxpcRUaLr0S9kdbAoPOL8lAaOe9lJ5p/+N3rXuDnGSnInIVxrGt2kDnhzBuUUZD+oPi01ka2Tp61UYK5XSddniXr1eRxPnPyLIDVm7O9PO+xGcPPswXnBbmXxfo8dfmVVx3Tdix72WgT67joPBEQAREQgdQjIIVF6rFXzSIgAiJwFAHjKmg9Lpiuy3U4KDEfXDDhpmZAz087ut3AGJno2eRhp6UXSutiyjjj+BlBVvfBIyfzElb38SrlreDDvD+fyrlm8/xR7lv4bb8xr7DlEkSXneZtm79ZH+UJwiaOeQlgebFlpx8v5/Z8Xv5xM9S0TafPnG39bOjoqW27ffEl7eJ3LEAQMsyZGV24Gm36PPx47eepd/rEMUkBSoN+TKzOkuyq9xIssJuMsgsVO7xjmA8v9u936TWoa//h4znmrC93/sJFsWIJ5+Mb6wrye7mLoiz8wp9uTA7IgxCr26BvJzZ5/+NuQfsUKf/aFcuXcJzA217uKrD+yGpcQpUp/0CVHp0+bO2ej5ybp2DhYoy7ezeurRdhDC/BO80W/WhtR0GChZAVGpAfV1RYLswyglH+x6ogWjl+jzuvF1yptWj/aW/c8+Cb3c6BU049JWlOW0GBs2yz2TzpemG4mn7Q6bPzjL+bDq2avs5vZ519btL1Es7CgkCpfvy/c91eYoSaVohTtETJ24gDMOqrwf1wr4P7qSRrrBlLNuD6jTptbJRwgmSvPvAbQsr3OvccaNzELLLWNlz3bgsPe75VSHzVv1d3L+ZYEPC7kaUe5Qedceb3W+88LEDkw3X1QsMm7840AW+5rpLb5YzfdccK6dw7emnfOx927YWVmW1zpPWCfAijECx67fykj6yZXj7ig6ynQcba73URKZ/RKycpLO43ftARCHVp1+rtcPm/mzxuNOt8DaNge9TMTWJSjP922DHCYs7Hmguhu5s7ikCUHVhnOOvhXhjuPki+aPfKoPXFOtdtW8K11bpH456NFUrXASPG585fqGiTenWecK6p3Le9rLFsu4YP+qKnO4g5ddu11H0NcgxBuBX28X+tuq81QpFOXmSaSxfMmcW6+N2KH37H5Yp1XegeI5SaBAe3AYRjnWfxsqBe1ke+cVvlbkeh4jeV5DcvxU5BYyXIsXD3sVj7RFwArvW5M8PHviIPyhX3PZL7E3FEuIZwU1i5xlPPcp/ub2IR2PbY5zmrgLO/23sT/wdd13keYGPG1s0bjnHZ5+YQaQ0MOr94Vug1bPyMZ15u2MTWw7WPkNy94cHvM1KQORvPmh3r/AjKKEh/3mzZrnPPr8Z9x3MC7cNimvhQWMM6Y0pxzG7EOf2MM5OeOXl27zdy6jzeRZx9Q1nBfPbzbMF5Qe5lsT5PnWQaT1227axV/UdPn098pVjHReeJgAiIgAikHoGjdoamXjNUswiIgAiIALvipk8aO/LOe+6v9FTdV98koF7l6k89i0Cv0/vvHBMrwMgud0ENv+G86NxY8o4yDz321HMNnq35EL6rd27fniQUbvp+x+7sgP333//9W6daxbLOnfOb1q9ZzbkPPPLYU3PNDmxnUMrNG9et5aWmzad9h+ImaMTgfr2mjBs5nDLZmcW38bRwTLDv0UY4cPf9lR9FoD7yq4FfIOSuYvrBy82wgX16OEea8ipUqfa4EcxMMLqagzfcXKo0gnD8TcczIxBsVa9dtx5lPPbMS6/eeOsdZYg38ZNRGhCYkgCS7Co75TRsQc7IjDARAREvcwN7duu0y1iSGLcfeZcunD/n3Y+690V4xm5g26bhQ/r1QmDQrN0nn3cycRwQHj327IuvFjZCkG4mqLbbLQ+WHnaHqle/rNDHKViw+SjLeGRad/vd5SsapcfmMvdWrIILlGcevq90PIzc5y43QQr5jb6P+2bYYPdxXPYgLEHo3qtLhw88+xHyUZ87X6EibYw1z0NlSuS3yjHyYxWy0AjV/bSbYK4oKNr3GPB1764ft8UCggCRKIt6Gbcz7JA178on+ynLT56d2w8rUYZOmL0M4TH11H2s8r0E4bbn22DTr7z1bhvjQWu5U8FEflxAMZcRlDWt99wTVujE9YLSw0sxiBKAeedHYTHnu6kTURw2NgIrxoG5jbXU5VdlzUb5XK/vde41ECHEqGGD+1nmxALxs0OWtYDxeuixWnUIqs5u+Hq1qj5gFTb0w+uapx7chiBAcQdht+yssBShm3M8vp86aRxKLOJ9GO9QZxtZ7Gn0izrbv9u4wedGyJKc40zdftcd4jE0fOeDj19/p83HXdq1fBuXFuUrPVqDcV69fMmiPQaW7Uuk9QI25BvUu5undQU7XxH8uNlwTpD1lOvL71j7uSai5bGCLnbDz5w6cSyWWeHOQajF9UJge4Tp7zdt+FKk8kd9PaQ/VjYIKXGRhDupyiboMOt0s9deqOU8l3sh9yjc5XCfwdrjW2Pd1KNj21bki3avJE+Q+mKd67Yt4dqK2yfm/UOP1a7z4KOP12ZdaGc2CYwZPuQod0asQ8zBZ155o2nXD1s1syxoF/c1d9DzaNcgx+d8N2Xi7WXLV3zyhfpvsP7Rxqr3lCzy1IuvNeIZpKZREqHE6GPiV/E/9yUCxNc06wSKY9bJUneVq1DugYeqoQBy3+ujzSX38XhZoDjPlb9gEdYWrzUJVzZsInC7XqIdBPzl2/msFLT9XvnZuMDvRgd8VHwKZ14ErM57jj3G/QmXS8OnLVyDGx8ULa0av/qC81zmxW133Xt/6049B9SvXe1Ba70Uz7pu41b5uT9FWgODzq//mWcN7qlPvfDqm8S+McYjV6G8I1YCllzOfvt9Rtq4bs0qv3M2njU71rkSlFGQa5D4N1zT3QeNnLzR+BflGQXlz2vGcsvdXt4L+O3Vpq3amcfln1AwT584duR3k8Yd5coT5Rr52Cjhp89B7mWxPk/xDMIayj2A+yqbrYzB3u/hnln9tFt5REAEREAEREAEREAEREAEDAGEepMWbdi5YMvv/5LYYYYpdzg4CMxtXr7Z3W+tHzCp7tTny1EzV//0B+XwsutVDi+401ds+61+k1ZHKQkQVk5esmkX5WIF4XRVxa47fkco7S4ToTZCZme7+n4zeXbpcvdXcuelrZ8NGTWFvNOWb/2VXctuF1GxTAz82NLv2et//svZjmh/j1+wdrv1A917+MTvyT9syvxVXu6XELA6y6O+J+q80tDdXvpDPnZFhusLL1XkKVuh8iNeeWA3a93O/eQZN2/1D/HuXvWqg5fX6Wb3LAJFr+MIsOdt/OWQdaXhlQdXGrRx7obdB+s1aZkUf8B+UCLN3/zbPyiz/I6pm3GPL8dMQ1iDcHfqsi2/NG/XpaffsqLl4+V26MTZy2DwQZfeg8Ndd7hom7Nh14FSZcpVcJbJmNC/eZt+/Ruhn/PYA4/WrAUXxtndDq5Ljt15b8XK0drIGH3Uc/A3lvHDNZ9+nnNeNa5bqJt2Ube1WOLYF99OmRNp7rnrfPGNZq3t9egOboryjrG1roec51KPm4nz+Odfjp0+du6qo6wr7HEEKc5rdeTMZRtxd8Jx+sv/0dgEOR5k3eF6cF7no2Yt34wizWlBRt2R1guUTMxdtws522aCi1PHg1Ufr+3uR5D1NOhYB2HmlZd7AvOda8YKNiOVadc5BN/R6kZYP2L6orWWPWsPsRxMSIXC7nMrGoU7x23er6cuWG3j5di8ke6V5AlSXzxzPVpb6zZs2hKeCKaxaPDixD2K4/1HTTtK8P3a2++1f+nN5u+FY/t8g8YtYGTvcc58uE2BG8cnL974c4Gih60MBoyevgC2/IZ1m/OcwsYacsaq7Xstd9rd0Cj3Ij2zRBt35/F4WGAFRbuqPvXcMYox1lHWMSxBvNrzdtvOPcbMWbnVuY4GaXe4vA2bf/AR6zTPVl55kmIomee/rybPW+k+zho5YcG6nyYuXL+DNZp7oDsPuy945pu1dsc+u5Pe5ol1XeeZBo7W4iUSh0hrYCzzi2uYtZ/6WXeffvn1Jk4XUc62+H1G8jtn41mzY50rsTDy2x/mlp1/PCfwrmCDirvby9zCGgPuzNfWnXr0Z2658/F8xlz1e50EuZfF+jxFG+s1freNXZP6jZw2j2fGWMdE54mACIiACIiACIiACIiACDgI4IaBh3V2k/kBg6CIuAnhXoL9lMFLoNdLBy+pTpc8zrKwoKhc/clnwpWPVQECDpQb0dqAX+1wwrxo54Y7bvtD3xCW4xscdxX0J0+BwsUwb2eXGX6S8UnOcacrJ3jyMuh27+Ssjxe+eys9UgNBrVUUebUnX+FiN9rAl17H6TtxLiK9+KGAQhAUqT2xsrLn4W4qXBm8sHoJutz5Yeo1F3kJRiDr9+XWlst4MY8IAOusCwEFcyzePsdyfri5ylz38pXMddTh80EjvOKbcA3xch1OeOBuH/zY/YnPbo7BZ9T3yzchzPIqnx3P7Er320/mFwoJr7mAELBd935fca34Lc/mO8f4NInkRxrrEMaZMXUqA1AW3nXfgw8Frc9Pfr/rDgKPW++8uzwCtHACMz/rRaS1ivmNIDWe9TToWPthFC0Pyji/c5e5xVoYrUx7HB6sJyiv3AJYdxnwZ366/bQ780W7VwapL1Ifos11P231wyjoPZN7SCTFEv3n+rP3MoS2CDcRRLMJwKtN9BVFNdaFbh/3fvqQXHncLJgvXA/h7jc8A/Cs5VU/91k/CrigbYchcUYincczSjzPcpTtNS9iXdcRVrNxxU9fo62Bscwvxs/v/cbvM1JyzFnaFW3N9sPMnScWRkH6w7NwpGdRZ3u4hsgfrh+szTaeT5C++n03iOV5yraDa9uPki1Iu5VXBERABERABERABERABERABERABDIMgUat2ndhlzrClqCdxp0alj0oPPBRHfR85RcBERABL6Ep1hp2l3JKKQxFPvEJsIMeC93kbGmSKyLNr4hIxSg5Z5zKEgEREAERSKsEFHQ7rY6c2i0CIiACIiACIpDmCZjdhoXx13zgr/37/XYGVzy4uGn6QcfufT79KMn11vLFC5NikOgjAiIgArESwHIL92VYJ9iAzssXH45vpE/GIsDueqwq16xctiS5eq75FZ2kGEVnpBwiIAIiIAIZg4AUFhljnNVLERABERABERCBBCOA14JceQsUJoCz36bh8qbPiImzbi19d/nnqlW8a+7M6ZM51wgV5/otQ/lEQAREwE0Al2z9R02fbzwUnlz13luL7t3z228EbCZYumhlPAK4/MGV1OrlS33fnyJR0vyKPofEKDoj5RABERABEcg4BKSwyDhjrZ6KgAiIgAiIgAgkEAGCLRMTYcGcmdP9NIs4CgT8PXTw0EEEirO/mzLRxJso9Nf+ffvWrV6xzE8ZyiMCIiACbgIENCbOzvSJY0c+/sBdN/+4dcumHHkKFFoh64oMO1lKlCpdls77vT9FAqX5FX0aiVF0RsohAiIgAiIgAiIgAiIgAiIgAiIgAiKQwgSat+vSEz/x4QLbO6svU/6BKnM37D7YsffQkQRAt8fafNp3aO+vJ8xM4aaqeBEQgXRKwMYTeK7+m81sFwkqPHnxxp9ffP3tVum02+pWBAKM/zczlqyfsGDdT+ECl/sFqPkVnZQYRWekHCIgAiIgAiIgAiIgAiIgAiIgAiIgAilM4LwLLrxo1tod+4ZNmb8qWlXZc+XNP2vdzv2fDRk15ZRTTj3VKVREoFS/Sat20crQcREQARFwE6hc/clnUJq+9Gbz95zHrsmeMze/lypTroKoZTwCpcrccx/j/1brDl3j6b3mV3R6YhSdkXKIgAiIgAiIgAiIgAiIgAiIgAiIgAgcBwK4f0Ag9PhzLzeIVl33wSMnT1/xw+8XX3r5Fc68ufIVKEwZd95bsXK0MnRcBERABJwECKrMuoKbOVzTOY/VqP1CPdaWc8+/4EJRy3gEPh34zUTGP2/BIsVj7b3mV3RyYhSdkXKIgAiIgAiIgAiIgAiIgAiIgAiIgAgcBwIXXHTJpVOWbt49ddmWX0zc7fMiVXnpFVmuQnDUqFX7Lu58dV5t1Bw3UdHKOA5dUhUiIAJpjMC9lR6pwdpStkLlR9xN/2zo6Kn9Rk6bl8a6pOYmA4GbTOwK5gWK8niK0/yKTk+MojNSDhEQAREQgYxLQEG3M+7Yq+ciIAIiIAIiIALHmUCmTCef3PKjbn1RMnzavnXz33/79ZdITbgq23XZOb5mxbLFznwnZcqU6b7K1WrOm/Xd1GhlHOcuqjoREIE0QCDrNdddf3htWXrU2nL1tdlzFCpW4pZJY74Zlga6oSYmI4FLLrsiy9ttO/f45++//273TqNX4yla8ys6PTGKzkg5REAEREAEMi4BKSwy7tir5yIgAiIgAiIgAslAgGC1Pb4cM+3q667PGak43D8QJLv4LbeVnjVt0vh+n33SIVr1+/7Yu5c8biuKh2vWfh7riy/79eoWrQwdFwEREAE3gX1//HF4bTn3aCuvF99o1hqB9fBBfT8XtbRPoPMXw8a8+1H3vmeZm0ik3iA87zpgxISLLrns8q7t32u+fPGCufH0XvMrOj0xis5IOURABERABERABERABERABERABERABGIgcPf9lR+dt/GXQwTGJngtO5SdxRB74pHHn35hzJyVW3G10fvrCTOjCY/s+VhkjJu3+geCc19xZdZsZ5oTH6759POz1//815AJs5ZiaRFDk3WKCIhABieQPWeefPM3//bP+5/0GoRClHUK13PJEWw5g6NNqO6/8W7bTozp+PlrfqxSo9ZzuCR0NvC6HLnzoqT6fs1Pf5LvzZbtOp9gPvF2QvMrOkExis5IOURABERABERABERABERABERABERABGIkQHBSrCwQ+JBmrd2xb/yCtdtnrNq+1/42c/VPf9Rt2LTlKaecemqQakrcesddnGvL4Xvykk27cuTJXzBIOcorAiIgAk4CtV9s8JZzXeHvAaOnL8hsNKMilX4I3FOxStVvZixZb8eaYOvcn1B8299QjJev/Ohjydlrza/oNMUoOiPlEAEREAERyJgE4t49kTGxqdciIAIiIAIiIAIicCyBXPkKFL7l9rLlrs2ZK+9ZxtfK/n1//rlj+4/bli6cO3vquFEj9piAE7Fwy5I127UPPlqz1mVZrsq6ZeO6tYN6f/bJz6bgWMrSOSIgAiJgCRS+4eZby1Z48OEzzzrnnCUL5szCzdyBv/bvF6H0RQBrvBtuLlUal4RXXn3Ndaeddvrpe/f8/vu2zRvXL5gzc/qMKRPG/H3o0KHk7rXmV3SiYhSdkXKIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIgAiIQIoRWLDl9xNTrHAVLAIiIAIiIAIiIAIiIAIiIAIikKYJnJCmW6/Gi4AIiIAIiIAIiIAIpAkCRlFxmmno1aG01nxvN2lfoSvP/jtNdECNFAEREAEREAEREAEREAEREAERSHECUlikOGJVIAIiIAIiIAIiIAIZm0BIWfGmofCUSReZ9IdJTUxaZNJ8/jeKi38zNiX1XgREQAREQAREQAREQAREQAREQAoLzQEREAEREAEREAEREIEUIRBy/3SZKXySSdldlfxi/p9q0kCTxpq0W0qLFBkGFSoCIiACIiACIiACIiACIiACaYaAFBZpZqjUUBEQAREQAREQARFIWwSMwuJs0+LuJlWJ0vKu5jgWGL+Z9I8UF2lrnNVaERABERABERABERABERABEUguAlJYJBdJlSMCIiACIiACIiACInCEgFFWZDL/PGJSHweW283fh0wqYFJHF67J5v+2Js02aZdiW2gyiYAIiIAIiIAIiIAIiIAIiEDGIyCFRcYbc/VYBERABERABERABFKUgFFWnGwqeMIkLCfsp7r5A/dPBNkmAHcFk1qZlM3VmBHm/y4mjTVKC5Qb+oiACIiACIiACIiACIiACIiACGQQAlJYZJCBVjdFQAREQAREQARE4HgQMMqKU0w9d5vUzaSLTVpnEpYW840C4h/bBpPvJPM3LqPOMAkrDKwvnB/cSI036bf07iLKsOCZHB4nhtKp5pvE/wdMQnGT2SSClfOBI+mgSX87uboY6l8REAEREAEREAEREAEREAERSFMEpLBIU8OlxoqACIiACIiACIhA4hIwgneE6p1NeizUyp/N9/MmfWWE6gjXj/mEAnNfZQ4Q66K0KwMuonAdtTm9COVDihqUOheadL5JP5h0uklXmFTEpEtMKmFScZPOMgklxTaTsFoZHvp/p/k+16S/TCJw+XqT9pq0PxxnL/b6TQREQAREQAREQAREQAREQAQSjYAUFok2ImqPCIiACIiACIiACKRBAkYQj0VAB5OeNsk+Y1Yyfw+LpmwICfEvNXkfMqmdo/u7zd/jTPrIJITye0xZ1sogTVAKWU9gRYLCIYtJd5iEggJFzpWhTqB4gB8f+ofiJ9JnozmIRYY9f575e5ZJX5u0yCSClx9UHJA0MUXUSBEQAREQAREQAREQAREQAQcBKSw0HURABERABERABEQghQlgRYDQPiS8/l96cnEUspDAtVMDk94IofzJfD9r0mjT1/1+8YZiX9xn8jc0CQsD52eO+ae/SRNMWmvSvkTk6LCgQDlBfA7cYj1nEkHI3X3yQrPC/JgrCrMt5rhVVrizouD51qQ/TfrKpN3RFEZ+x0f5EpNAi75cGkeUhPbvf80fpP+9Vb1YYjZcrRIBERABERABERABERABDwJSWGhaiIAIiIAIiIAIiECcBEKKCNz8IJRGQM9u+stDAsNzQn/jHgnh9VaTEDizQ36PSQSgxl0Su+wJSP1vIgrivRCFFAy3mmMoJyo78jxp/u5n+kGfAn1MmTC8wCSE9o+aVMMkLBLs50fzB+6jiHux2SRiPKSaEiiksGEsaSNWIqVMQjFRy9Vx3Drh9sn9+dX88J1Jv5u03STcPp1nEnOCvmFxwf8oKJaZxDwradLNJuFKC8WIkw/nMf/4TDOpt0lYYKwIojzyaKd+SiUCIYXEkdqdCghzjPc5EvFO+BDbxP6NwoJj/5hzjsSPSaVuqFoREAEREAEREAEREAER8EVACgtfmJRJBERABERABERABI4mYATVZ5pfUEogMEaAfJNJKCNQTBBPgN9QTNxjEkqJpaE8CJERHiJMfM+ke03Ka9IGk5aYhPXARpOIcbAjVBaukRBeJ+2aTu0d8yFFBUJ6FBPEmEDQfplJfG4xaWY8bQwpgGBGDIeqJr1m0kqTcpuEUoAPHLEkmGwSzFFkEMMhRQWzjgDZtI+xL2MSsSdqhtoV7gtXTQVMwvJhiEmDTcJ1E4oMYlKg3GF8bfv/cSquQooRK5jGfRTzD9dRzEHm2I0m2cDla8zf2R0Nocw2Jn1oEnMJd1FJu+/j+YSE5UcVYQTjcZcbT5vS47nhFBZbs2TeAAAgAElEQVQOZQXXIoo+FJ5JSk+TUFqguOIYvyVZOml80uMMUZ9EQAREQAREQAREIH0RkMIifY2neiMCIiACIiACIpCCBEJCY4TEF5n0qknsekdQeHeoWoTPv5iEsJAd8wiKUWQ4PyghsLRYZdKnJpU3yQqabb7x5o/bQuej9CD4NDEKEOBjsYHwEcUGihErjEShcSg5BNGu9ib9GxLU0/fCJtU1qYJJ7Pa3H9qCcgE3UJ4Btr3KjfRbqE76nMekfCbB3CmI53TcT80waaZJxLlA+I/AHsE8bPj8HZRLaKw5F4EvCgIUJQTExpoB5YBtE9/hPgiOiSvRzSSCY6NkYJyIxRE3oxAfnucZB8Ymh0koMFAeEfcDCx4Sv/FBIdbVpCkmrYq1DS4XRNRvXQ9JWRFhMiTnoZCygnEnHTKJuc63VXgxLqxNrEXMYeYbx6W0SM6BUFkiIAIiIAIiIAIiIALJTkAKi2RHqgJFQAREQAREQATSI4GQVQFueJ4yCVc8uEJCmYADeXbZIxRcHPrG4uB7k3DnQxyDa0LnsIsehQZCeJQWuDQiCDOfXSbhCokPO+9RTNgPu/NxC0S99oPFAcJIBNII61GAUCc7+BFOIshHsYEQ2QrucZ3k2wIh5J6JfmHtQQDtaiblNImYFc4PFhAI5X8PqhhwleP5b0h5ADPcRPFdzySrJKJvtNH5QVk0ySRcIaHEWGcSvGGPCyZrsQI/eJAYGxKcYY/jfxRSd5pU1KRzPRqH8sGptIE74zHSpEEmYQXCeKBI8s3dox5fP4U4IaSmreVMwurjNo+TUeg0NQnF2M9BxsyhrLDKiaT3Ce3c9zVEyZbJjANznmDuzGHWmSRlhMfHqbiwawEuoqRcSrbRUEEiIAIiIAIiIAIiIALJSUAKi+SkqbJEQAREQAREQATSJYGQsoJ4CsRqON8kFArWZRO71RGITzYJYTgCYwSIdgc9gkGEiU5f87gTYtf71SbhOgpB+WqTCDiN0oJYByg52Nk/yiSEz9E+WDgQZBkBO23A5RDCcsqjDJQjtIW2WwsQrBEQpNMeBKC0g2NYEpQwCfdOCORRFFhLEVxbcQ5Cf+rsYtIkI/Smrpg+DtdCnkJU67M/FNCaduKK6SGTiBWBtQvtDPdBEYRlAyz50EfGiXJQYKCcQAmywCQE+A+ahNWE3+dkykKhhLUMlh7wTRr/IIqACO2P6VBozjKPUOwQEB3FmfvT2vzQwyRcmeFOS0LsmGgf35PM9cI1ynXJvP7DXB/7IrXAkR/rIK5dFJmHzHlHFJnHtweqTQREQAREQAREQAREQATCE/D7IiaGIiACIiACIpCiBP7991/3PSlJcHbCCbpVpSh4FR6VgBH8IhjEsgB3RAi9CXz8mUkLTUIwzW5+XA7FtIM+JIS3QXKt+xYEiygN7M7psuZv4iTkN4ld/VhaXOdqPBYVnGM/P5g/8GGPQN/9oc2bTJpvEkJPzkN5gYUIFgIoKIitYeNF2PMnmD9QFgwIJVxg/RFr322hIYVFWGG5M8gw54RcIdE3xgPFEUofFCxwQXnhtgCxVTkDEntgOeonFBsoeSiTMUcxgYKGeBlYt0w0CasWFqm/DIOk4N+J9glZXaD8wkIGBQ8KGeenk/nnk1D/fjL9CLdTP9G6liHbE1I+sE6gaON7tx/FgzkPJSaKSetCCiUHSgspqTLkTFKnRUAEREAEREAERCBxCfDgqo8IiIAIiIAIpDgBo5DwqsPuOLfHrFsXG3g2KcBwijdOFYhAGAKhXerETCCoMbvQx5qE+yV21O+LV1BPtaYMGyjX2QqsFbAMsML5XubPfibZwLoI6tkxj/CR8xHYYxWAeym7k97GLbBCepQUVpDPNzEhSM4PygjyU65TWYEyY7pJCLexJtkaVLDtDhzsqPSEoELTkCUACoIDZoxQIuCaa6hJKC9wh0TfUTTQz0dMIu6GDURM1fQHV1FYVhDI2+tDP3HthFspFBckhPkokbBGiDsGRZh6k/Vn5qhhRF86mMS4DjMJF14opZhPz4cS1jmtTF4UWTtlbZGsw5CchdnA6yjsmIN+rSTIhxLOBuhG2XEk/khyNlBliYAIiIAIiIAIiIAIiEA8BLRtNR56OlcEREAERMA3AQ+FhVVWIDzhb6cfeoRoCE0RSCYpLWRp4Ru1MiYTgdDOdBQB15uEgPe70Pfu5FBUJEczQ220gngEkAjr2UVN7AWE8bgEwoUVu7FxeVTAJKxFEOYj8HR+sKxAoEn8DSwnrGsjrCqIB4H7JCwJYrIkSU6FRSR2ISbWYgU28MAtVlaTWFuwRCER04IYAChmiFtBEHME+nzDgfXHBioOHLQ7UhtT85jhg0UNSi3mR3eTUFzYz7uhsSf2xsqgSqnU7FdGqDtkicQ9Ewss5jRu2X53WyCFYxGyzmDcUXgyx3ENddCcH9M1nRGYq48iIAIiIAIiIAIiIALHn4AsLI4/c9UoAiIgAiLwn294BC/WrQvCQVxU2F2fCBn5O0lpYT4IVI6xtpAiQ9MpBQkg6CemBC6VEAziBiphlBX026E8sFYaWA7w2RJym8TfXEdcZ1xv40wi1gJ9I6Es5BiWA1hgcN39aBJujyiT64+A0Sll6ZTsO7xDTJwCWCwiSJsdCh64oICxn39TsI+OalL/T9PPvYYDcUhQ1lQ0CYUccUiWmLTcpIImMd67TT4UO/9kFDapPzpRW2CvV8YOpYVVzEU9kQwoJozSwgaK51rnupcLMF/0lEkEREAEREAEREAEROB4EZDC4niRVj0iIAIiIAKWgLWs4Jv7ELt9rW9thC9WYYFw1f5tXdpYV1GiKQIpSsAIapmT5U1CqIeAr6NJs2K1LkjRxoYp3CFkdrucwpJim1VoHC9hdJhd4CmlCPGk4hq/41p3asyBcHWGxvyPkKsoFFQVTEJwjSD8stDf1vot2ZVKicQijbXFzlnGyrqGCjo+WFVQDudxb5XFfRqbBGquCIiACIiACIiACKR3AlJYpPcRVv9EQAREILEJICjBqgLhCb7mEZbxQcDKrnZ8+LP7G6GK9dXNt2JbJPa4punWhQT5xIPIG5qTuMcZllZiFviFf7wUFX7bk1by/VXrSEuPCHpP7Z42Y+2E4qfsMXMed2EoiFHQWWs2rGwyrFIngecj44PCgjg3fAKNEfFiQlYWjLdcQSXwQKtpIiACIiACIiACIpBRCUhhkVFHXv0WAREQgdQngJCFnesI/VBW4I8b39q4pWHHL77k8cdvgwTjmgQBDQnf23wCCWpSv8tqQRohwM5y5iMukzKbRLBpXArpIwKWAOsW8yRpp7pRYiD8tcrUYygZhUZCf0LKKxTFWF3MMd/OGCAJ3fYM2DjmHGPlvBcGwhByDcU5SVaNRoFBHIsj91Mbb8ZvbIxAlSuzCIiACIiACIiACIiACEQhIIWFpogIiIAIiEBqEbACP5QUl5hEUGCEw/jl3mwSygzcRaG44PdfTUJIY/1tc9wzrkVqdSjR6zVxQI5x/WFigEjpc+zA4RLnTpNQWCC8XS9rhESf3anSPuu2jjWLv61CNU1fUw7lRapAVaVRCdj7YFJ8mai5w2QIKS3kDipWgDpPBERABERABERABEQgxQgECtSWYq1QwSIgAiIgAhmJgBXmISjBBRSKCoQuWFIQ/DWrSSgx+KCsQBB4jUn5TcJNFELk8+wxhPAmZSR+nn2FQSgl8QilE833STaZE9mogIstvkkc07OAg2goKPMj5qecJhGAuG/IbU6Gn2MpAcDs5D7B7uZOifJTuEyuHZRb2U26OvRtLcJSuGoVnxEJhKwgrEtE3CnG+0HpjwJEHxEQAREQAREQAREQARFIGAISUiTMUKghIiACIpChCNjA2wT/tC6hcP9Ewh0UvyNQv9QkFBp8spmE0oLfsLxA8J7h72NWSRFiYYOWo+SBz6km4ZOebxvAHJYcx2olSXlhyiA5FR1W4ZGhJmWos/BCAM28HG3S1owI4Xj0GWXF8agnheqwWlKUrsyZLKGEAoPrSx8RSCkC1iVU3LGcHAqQlGqryhUBERCBdEXg/AsvuviUU07luTruT448+QvGXUiCF3BSpkyZzjzrbPsul+CtVfNEQAQSiUCGF/Qk0mCoLSIgAiKQgQggqGRnJy4tiEdxhUkI+vABjyDduosiD7tIUWTwsIsSgxgXCGouNgkLDKv8SNf4HFYTR5QJIRdPVhFhhVfwwEUNbBCkwo1d31im2KDmCFQ5Bld+52+UFxla0BoKtm0Z4d5nn6wrUu6yQlgaSilXScqWzHq1x6R1JuGybq9JF5qEhZhTQZiyrVDpGYpASMmAVQT3x+QImi0TxQw1g9RZERCBWAkgeP9q8ryVT9Wt/2asZdjzKld/8pkBo6cvOPGkk9L1s3f1Ws+/MmHB2u0oeuJlpvNFQAQyFgHFsMhY463eioAIiECiEEDIgmAdoR5/rzfp8pCwjwdaBOm4hrrRJASCKDPIT+Bt3EbxQTiIwgOh4cGQW6hjBC8mRkOi9Dm522E7Zq0pEGDBAuUD7KwgC4XFbpNQDFkXW7BGMA9/gklzLuXZYOYZ2UXIdYbDLpNWmrQxuQdN5aUrAriywxoM64qrHdcUCtixJrF2cS1JIJyuhj1hOsPcinvzmTPYtu2Zgm0nzBirISIgAglEoPANN5U8+5xzzyt8w823xtOsMzJnPvO5+o2aH/hr//5//v47XT9z5ytU9IZMmU4++c8/9vLepo8IiIAI+CYQ90Ou75qUUQREQAREQASOJoA5NUJzBOUI9paY9FtIAIPbJ1xAcfxakxC6I/Szbo4Iys0DPop3K2zPKHytogcW1pICKwnifKCowJ0RzJwJpQb8LjAJYSp5UV5gRUA8EBRCxAfBuoW86VbLE2WSwJS5xkvVZJNQ9OgjApEIsGaxDvFMfZVJXJM3mETQdq43FIgZ9XrSzEkhAg4lQ3JYWKRQK1WsCIiACKQvAoWK31SSHuUpUKRYPJYRVZ+s8xIWB3v37MFqPF1/sufKm3/d6hXL9u/bxzuHPiIgAiLgm4AsLHyjUkYREAEREIFkJGCF7kmBn01CaM437lTYtXyJSeRBGYHAD8uKX0xCkLzBpByhvFgE7DQJywLOI6XnD0yscBReuJ7hNxQWV5qE4gdOW0xC+YC1Cu6gUADxN5y2mcRLA3+jxLBjwN+wxmoF7ul6x1eYSQLPoiEOv8gdVHq+lJKtb6xBWOPgEoprjmuIa7OMSQiTx5jENSori2RDroIg4GUZITIiIAIiIAIpR6BQsRK3UPrpZ5yROXvOPPlWLVu8MGhtWGg89uyLr3KesTrguT3dfuCUJWu2a0cM6dcr3XZSHRMBEUgxAlJYpBhaFSwCIiACIhCBAII8BOIIztmZjAsoBO3zTUK4jvCPexSKix0mIRS0LqOwvMAaAFcsKDJIuDWysS3SlaA95OrKKnhsfAqrWLCxKawvfRQ+KC8Wm4Ryp5BJKHfgi1IIZQUKHr7hZ/3JWkUP+RgP+BM7JKPt3sWiB3dQfDOn9BGBaARQRLA+ca1w7WC5xNpFKm4S69q8v2odWZ+OKu/U7tGK13EREAEREAEREIHUJnDqaaefnrtAoaLbtmzacMWVWbPlL1y8RCwKi5rPvvSaCYXB8/b/9u75PV1bWFyfO1+BE81n2cL5c1J7/FS/CIhA2iMgl1Bpb8zUYhEQARFILwSsRQTC9jNNQnnxvUk/m/SjSQjV15pEPmtZgKICC4DZJi03CeEgbljY2YwrFoSE6c39CvdqXBXZPuJKC+UDzFDO4MII4Tq7tDgGA44hSEV5QbIKD3ztI1yFKdYElLvdJF6YOA+enEs5/2fvPMDsKso+Puf2rdnsptdN74VA6EjvIoI0RToiyqfgZ+NTFEVAQVEEpQhIEaRJkyI9SCghIQlppCebXnY323dvPed7fyd3lrt377bUzWZmn3nu3XNPmXmnnfn/37JfBQ2WgNvUF5daEDovSwZoNslIoD0S0LF01svJSyXrgMjEQ4EwZAwy1kwyEjASMBIwEjASMBLYByVALAa/PxB44clHHyTuxMQpU4mz16FUUFjU44LLrv7e2tUrl9fX1dWKgUWXJizGjJ80BQF9Pn/Opx0SlDnZSMBIwEhAJGAIC9MNjASMBIwEjAT2hgQA07VGMtrsgPEa3CP2wqmSj5Y8OblW4eJojWTIDLR0sADAuoBPAHYAfMB2gHbcsexzCUuKlGzJd49kTSJAxlBPiAfICawnkBsaWvjJR3bnSj5G8njJgKQQOZA+mKvjRgtLFTKWKpi0cz9igXAv7WaK74CtyLArkj+t9QvqDKFDX1LiDgoizSQjgWYSyGAVwXzGWINI5XOhZCyUIC907J2MBKBYXiiySUYCRgJGAkYCRgJGAp1XAtod1KyP3p+2cvmSzyceePBhHS0t1hUE3H7k3jtvDwaDIYlD3aVdQo2eMHlKLBaNLl+8CMtvk4wEjASMBDokAeMSqkPiMicbCRgJGAkYCexCCQDkAY7jmgiLCjT+x0kmKDQEBoQEwaAXS8ZNFOA8IPsxktFYRisJzWaAQMBmAiTzPxYE3Hdf9Bmfah2ilQp0UHHqCHGBlQlWFcgHWWEtQaBtHXuBWBaQPtp6gt85D/dPkBj4218pmSDnBAfGsgVrAogPzoUQoRzIMSakiet/37K6muGK1KppQrbFSRl0KbdizWpqDuy0BNJIC0dIBwguCFTmKuYirHQYNIxbfuM4Yw0Lnn1xbtppmZkbGAkYCRgJGAkYCeyrEphy6BFfisdjsSUL589d9NnsmWeef9HlxKOorqpsl0Vu96IePc+/5KprtmzasP7Nl597+pe33/1AV7ewGDth8oErlixeGI1G2FOYZCRgJGAk0CEJGAuLDonLnGwkYCRgJGAksAslgIUFGZKBBCGBFQUxKXD3NE8yZAYg+lzJAMqcqwNwa4sKgHsIeM4DHGRt25fXN+0HX1ueUG/IHD4hIiZInigZ4kKTF9QdIgINb6wktMsntLwBUSGEIDB0kG7kBXmBCyRIITS8OBegnu9sLLBWUUJU7A9kBVXVbsnod/Qxk4wEOioByD7cQjF2RkoeI5k5jnGG1RMxZYg/Y5KRgJGAkYCRgJGAkcA+IgGvz+fbHrNiwWfRSDg8f86sGfJ+bI2deADKQu1KWFcQhPqRe/50m1duyEVCWHRZC4tAMBQaOmL02EXzZpv4Fe3qIeYkIwEjgXQJGAsL0yeMBIwEjASMBPa2BCAhiKMAQI/mMe6LCB6NBQDWAoDsJNxB8fuHkvEby28A9Lg4guxAixmwn7UNwN21DNjblevA8zXRAjEBqImVCZYUEAm4KYKYwWURBAMa3ADsR0mGZEA2BCPHGqVYMoQF/mKRA9dhUYEGGFYpBJVGNviVRVaQRFXJ+yIvAFeupxxesbAAcN0fSAtkMTspI6MJJoLY0+nmxxv3tJq008HgtQu5FsfzDd+cuqeLm+l5eiwypsZKPlAy85eOLwOZSFyeVYypzlBgUwYjASMBIwEjASMBI4HWJTB63MQDcOU0f/bMjzlz4dxPP+Fz/OSDDp4xfdpbbckP64rzLv7Wd0u3bNr4/JOPPdhdYllwTUNDPYoOXTKNHj/xAIieRfNMwO0u2cCmUkYCe0AChrDYA0I2jzASMBIwEjAScDX1M4nBTgLiuEohA7oD1mMNgDUBmsoA9F9OHgM8/4pkgHwAdTSXscIYLZk4F8RrgPjQlhmdRvTEp8iQtFB0zAjWZYgK6o8FCWQF4C3WEJAVfFJvCAz+Rz7vSEYuaHS7GyBJyBDw9Njk+VyHWyisLSB2cKmFixqIIggjngmYynO5jsx52nKlS4OryYDbgMpYolRL/AoNlCfFaT72hAQgHYS00LEe6Hv0b8YB44T+qINb6z6608W6c95Z3FuTmzpui7b+4v70fef6lQ+nP4tyMW7cuDIyIXFNouq1AsoJcajLzhhmrDEmIRqZ45irtGXZTtfB3KBzSsB5W5a9EwwxtSdaJ4XsTH3RaFy3OgmhuSdEYZ5hJGAksBskMOXgw1EQUvOShMXKZYsXETR73OQp7dKW0NYVd/32l9djoRHKymKvosJyk91Q3E5xS9xBURDcZ3WKAplCGAkYCexzEjCExT7XZKbARgJGAkYCXU4Crga/ZABziAZe4gHeAfwA+dB21xYF/M/vgJoAgVhZYDnAcQB7bUGgg0d3ZqA9layg/BqYRR7Ek4CUAdgk8DjEDFYkEDMcJ0E+bJQM8AkhgUxwZ4TW1yTJED7Ik0QgYKwHtDsaZKc1vyGK+M59OJ9P7aprf4rlQF+hr+0S8/zQ85W0B32Y+wJiayuBZJM0/QifTfPuuSTlo/9pckCPEz0WmxVkT5VPgEVbwEcdQyUUkyL63e7ojnsINfonhBJ9U/fVDo/zJFHBezCWSprg1JZMxJngmHYTFvvdsMsSSdKCccoYxLKLOUePFQLar+t2WuVmIS3oQ9yDeQtyUMehYRxzPpt33SdcWQu43VrSc0WL9RRg3KS9LAFpQx1PiZLQtzxyjHbW7cd3yGn6MW2pCeHU+SEzs72ft28KIZGplbV8NfmIjHWMLI61OK/t5S5jHm8kYCQgEhClEeSgx6+WCeNYj93UebHZHClKJrtdjsSv4CHzZs/4iE9b0sLPPp05blLbhIW2rti8cf265//56ANcHxLfUHw21HddC4txkw6cGhYTEgKU7/YGMg8wEjAS6JISMIRFl2xWUykjASMBI4F9SgJsPgAg2bEAwGMJAGGBJQGgH6Akx3tLBnQHxD9eMtcBxAMc4kbK1Y6XrEH2zhwlWoPFbMgAQEGrIRM4Tj2HS4a0IEYFICcbG7S0+eR8LEnelAzQxblcj1so5IG8CKZN4l6AaABkyAjZAaJr7XVcQWnQdnnyGuTOca7rMBCcvMc+9SGbXVs2zNS5Sr7vcJ2TJIDW0qethqbIknbBHRfadB1+hgDsqTJNBej0vfRnRldo1016ofF6KSdlpJ3pF4D09Cnau0QyZJZrVbC3GvHm7BGqpx21PMqxY5Yn0seOxI6PljndnBjl1uCudqGWXv82iy2y5FrICIgHyL2FkhkbEJ3cH5BkvGQslKASmH8CZ/d8pP6V8q/3jNpBxhXXnyiZeQfy8BjJyyS/ecAxczbMfW8KbqGmS8b1GsQG5Crtr8ceRGFLljx6XtCWHvxPYm7T82XykPnYExJohVBivDGOaCvGFBaBtDNjij60Ntk/+J3+RVwT1jcILqzk6FtcD0FG/+E83Qf3RNX29WdokFOvV4wV2kETxdQvKoSHy3oKIbrX5rV9XdCm/EYCOyuBJDGRehvGL++kZMYt7024fGUcsxfgvZiYYqzRvKOhoMTayXfGMtfrdXFni9fi9cSqOGDqYUdu3bxxw+YN65nT3bRA4lgcfMTRx/Xq068/v7V0g4u//f0fEbvijzf//Ec6+LS2sBCPUF3WwgIyZ/HCz+bYicT+pPy02/qhubGRwP4oAUNY7I+tbupsJGAkYCTQuSSggQVe2tkI4GYFELVYMiAO4A/fAXsACnslP6kFIAQAK0QFGjyAQNp9DL9nBG87QfUpF2swmzNAU+qr/fZTJ8gH6soGTpMOAKAAW4DgaG6XSNaunt6V72z4COwLgcEmD5+6bBK4N5s/5Iuc+A2Sh3vwO/cEcEW+PFsHLNdg6X4B8OwMUSEyU0myAlkDWCJPwMhTJNOWyJRNNzLHAkaTFh2RbapFDo/kfw1ke7PqI8r2enyRoD83FI4mJNdJ4JHoiKXrElM/Way+c6VSDw+61Hq91ymh6Ym6vmFPqF/C8nIPTPYB1SnfU5JLJEOu0Ff2qGZyilVKj1JPYJgQFhRwS41Ep6wM9tn85ejWml52hDprC4sOlS9pVcH1jDnGCnOHtk46Tr6fKhmgGUsm2vBgyesdZT2UcHxZxaHlZYODK2pKwiOy445fmC3raPkdspAxxOccyfmrsoe+ce2EP3/+5wXXMifRxjyL8UVcHhKuJT72jldbJOs+wHzAsxnzkCGUgU+XSJPMXDFfMufxv3Yp1ZE+lHy8+dgFEtDWFLQXbr4gmOkDxC6h76Dye4TkRZIhIIgpBNiGli5rGO1Hn8Mah3WLvvhism1xKca8wfxMXzdtnLnBUskKTWAyhrRLRH1VI1gGcWFIi13Q+80tjAQ6IIE0okK/uzAPYoHIuysKOSMk8x7Cesn8iMUrxyH8+Z/r+I35kPcoFJp4P14k909XWHJLt6ssL4aNHDOumwSdeOPl555Orfb8OdvjWYyffODB776+8QutkJSTCiRWxfmXXHXNhnVrVr/45GMP6Z+CEpCa713VwiInNzdv8LARoz546J47O9BVzKlGAkYCRgJNJGAIC9MhjASMBIwEjAQ6iwQAZgAbAHMBa3iZXyqZTQ0bFjY2/EZGG1q7NKL8xZLZ6HAOpEeqW5/OpNmT6rJCa7cDSmotM8gZgK4JkjmOxi1xJiZKZkNGvArIBkiLY5IyACRHaxc/ugBfALIasMGqgvpjqcF9AT35zj04DzANywpkTEZ2gGvahQ3Btg1YJgJpR2LTTRsUSy6RfIbk8yUvkUw7IG/A8cclT5OMNh4gpav5m2ZBoR+nSQrAON7ZtGVEP8txegpJ4fHadt9owN/Tl0g0xCy1wZuwc6XB+njjiXXdqurCubUNJVV5eblVqqBsS06veL/IpkH9Gzb0qvQX9N4WKJwUt3yApgCuJID0uyUTeJ0xRrnj4g5qt/eBJFlBH6Qs9OfetrIg6eIJZQ3Z5AnFHg/2f+d/G1bRxxvL00HwEXAZAIR2wmXaXMnExDlZCzz9U0iJAQnHe+O2WM/Y6vDIjdviPetiTgBQWicdUJv/IX7I9a/2Pm3F+OoFzvkbntmUH69mHuO5/5XcXUb7ZKE4Nlk9m5BCxfIbcxrzmx6n3JP/Oc4cwDzIOGYuwMqKOQ/ygvHq9gJbrygAACAASURBVCOTdqsEGI+aqGB+Zi6lTRg3jG/m4sMlA6rpdFryC+tbS/suCArWvg8l0y8hO2ckr6ONIQ9NXJ2mTavbQisl0P+1ZRJn6rlVExn6fIDPzvROsFs7rLm5kUAnkgBjkDUeC2Csz/i+UjLEP4nfeS9i3ed37aIUKzS+Y22Mi1TmUd6leF/mHryrkHlXfk0ya7JrJaqJkp0lLg5Ixq/4bNYM5ujGNF8sLPhnO2HxckbCQseuuP+G3/46Ho/xfu0m4St4H1G4TEq9Z0vffT6/P/X69lzT3nP6Dxw8pLBnr95rVi5fWl1VCbHeZiKYtsTmc1qynsAdlEfSorkmfkWbwjQnGAkYCbQoAUNYmM5hJGAkYCRgJLBXJZAMxs17r/ZJz6YDAAeNZMA6zMK1mwz+R2uZjQ3gEMcB/rHKADxik8KGR/uwjst9sebe7YBrO4SYqhGvgWeASAAVtHMhEchs1ABs0S4rkQx4DAAGScFGQgfiRrsM0Iy6AZJB1qyQ/Irk0yWjyYv2PEAY9yhO/o5s2RACurJ5ogyAYZRPu9LgntrCQr6apCUgwHq6MDQQhvwB/7FwYUNOvyXRnjrOypHynXyP5Mck4+aAzaqjXTYRqJeL/tzTDQZN38j3x+J04dyY13dMViQat2y7X9zr5T7F4VBggPTwsoTXW1u0rWZVTV5WrjduF4uFRaBHaeXrca9n3epBfftssAaF60NZ/nGVCwpH1C9b+l73Y476oOjIKXGvDyBdJ/rLI5Zy7hegnn60QciKxg32rugFLchPE3bICtdJgBiXS0ZD3U3SIRvqLe/V4i7qX/Iv4IUL0Ov76RgbrRA/Os4NlgsXSv5ye+sTtUNqa6yvX4iKwTWJZi7DGD/p6e7SQM/oDWNuniWWLJu+t/ovc6VVT5J8hEAt3ayAjPcsNckKuWOceQuABaAaYAYCgjkQ4oZ57QDJaJ5SbsBrrDQukAxw8oxkZOWXfsNvLQbyNjEuWm/tdsQQYU2BSGLOZZ4eJxkSiX7IXIplFW3VUmptzwXpwf1pVz0XnyTfsdh4Q/KzUj7mfdZEfm9GTu2n7cu84cYKScmMc2QEscf4Yn7V7u/4P94ZrSwy9D+t3MBarN1dtUhK7qft38pwMz/tTQmkWVS47zGSmTP/RzLvt8xnKETQv/kfUv9VyayHKM6USGYt1C4q+eQ9FrKeeRGygjWT9xcIXd4JUETgvQsyn/dcrt8hF5zpsptyyPaA20JYfJD6W+W28rK1q1cubymOhbauKFmxbMmrzz+NskpjCopPKP5paGjdJdRxp5xx1tU//NmvR4weN2GVxIK45qKzT011S8U9cEt10hlnn3/7L3/yfe1yimd/+7rrf5mbl9/tgbtuv5lyptfL7w8EfvvXvz95/KlfOZvfYrFo9MG7/nDL3+783U3p5+r/R46dMOmHv7jljoMOO+oYCJQ/3XzDj5965G9/ST9fy2TB3FlYw7hpxJjxE8+64OIrLCEy/vWPh+4jcHlLzzHHjQSMBIwEkIAhLEw/MBIwEjASMBLoTBLQxAQbEDYa+PqGyMAVCqAO4CkEBZ+Ac9odFGbhbFy0+x3Wt93u17Y9ghPChNO0prx24aNd2QCu4J4GLTE0xgBX0BQDWAEIBRhjU0ZdIWhOkMxmTbscAWCmngCeWruUTRsAJ/dFk59nsLljs0g5cFvD5pD7s2HiNzaIFFTLzJAVIox2JG35QJsALtOGuBHSZAW34DesLQChdfqufKHNAJk3nO1/0X7ibVf+tGGwzJfvP7h+SWCjp8hTofJGCPnQLRSNOKWF3b8V93mH+xKqPhIMDHEdKWxPhXJcGtcBMLUSXo8KZ+UrITK+K9BmdEPP3o5/tb8it7qq16bsPvbi0LiyrcGeqiBWmVvnpdhNk9+OHe9RdlFWomFd7hMLli6cNoH+52ostiST4IMt/dLmcfokhaC/QlgA1KJx6QakTEn01UclMw4ge5Bfe7TOaSPuz/wA8Yf2ejpZAaFEW0AKNEnCd6rKeKFaGx6mNkcHKiEv9Fhuq2L3RzzB++8fdvXjF5Q9HeoRL/eKOUx/K08Nlpxl9VNjrByXVGQ+YzxeKpl+w9wGoQjxlSmdmTzI2NdzBSQP/QughjnRpF0nAfoPfY+MnBmj9NNzJWvriZ19ml4X6A/pibm8RDLr3+uSAflYJzrkDm1nC9hJr9fWLpbP5wnI7OSJJ+wcj8cdoo5tO4x77Rtfk5yshw1CWiQ6aJ21UyJogRDTpESqtUgqAQM5poO2A/iipMC7AfMx7a+tS3aqbOZiI4FdKYEUsoLxyfjjvYj1irWb+Yx+PS/Zt3nXf1Iy1gklyT7tKnEkM0VL7edYKWqCkvHN/Xhv1eOcPQPzKL+xL8AN57tSpoqdcft5wMGHHVVXW1uzbPFC9iJN0vzZMz8+5uTTz3Q1o5Iv/PqEy777g58Su+LeP956Y7olQlB8QnFeaxYWl37nup9c+7ObbuMZTz18/91nX3jpVd/+wf/d+OsfXXNFaiEuu+Z/rz/0qGNPfPYfD927dNH8z7oVdC98+Lk3phcPH+m+04yddMBBXzvuYPYATdIFl171P5AVWIesWLJowTnfvOLq7wg5MmP6u2/xzPTzDz/mhFP+9NCTL24rLd3yxN/v/fNRx5502rU/+81tr73wzBPplhnjxOpkW1np1o3r19KuCrdYP/7V7+70eL1eZHXqmed8/StHTR7RXouO9LKY/40EjAT2DwkYwmL/aGdTSyMBIwEjgX1BAmxQACB1QD1cv0BaaLNw6sCmHcCR4NtYDrCOoTXEMa4HVAL85xo2NdrX/d60sNCgCuWnfACxHAP8YnNFGSFa0NClLgCPaOjreB0QCnqThiUGRAPnomEPgPGyZABeNiMAstwTMBdAg+dhRq/BDeSkNXiREZtFnsf5bAq1OyjjXkaE0UbSFjP0QbQCsQYg00Y64dILoJGUasnA/5cKwZBfYFU9XuvkLn4/fmTDwf6ZPSt8uYFST7chgUR8gtj/J3J84UNtnzV4W07+sKjPR59Q8pmxaHXZISu3oUEQVVtVifJeXf8sAdiDASEfVMNIX5/Py4ep12u+5hFCok/Qjjqlvp4ZwfeoJzBc3Bj5JlXNP/68jc/E5uVPqpxUPY8+wtjcle5UGAf0ZzQs2bzjnunYNuSOP2RcOTEHtEVKaiAQ0ggQgxgVX8twf+YV3ecB/F3NR9vxqNpEN7U6PErNrTlM1SS4TfuTWKl8uzaQU/bMgRe8e+WWhz7I6VZ/ppUrYzuobCtLLKK8LsiChuFXJetGhcBoiaxIf/jv5QBzwG8kM+4Bgj6SDKjZlmzaX5H980w9vrUbMfon8zKWVN+WDAi3OxPWVxAjENaAeczbzC1/S35He5gxuSvH4+6sz07dW8iFJtcL4eD+H/B7PVkhf8J2VJYdd4IebwIwLE+QQxWN2/XKcXhPEO7CYW1jjNGu2kplb7wXpJIUEFWs5cwDzIN67eZ9gLLiXo5+pt2JAfICmKaa+THWqdveqMtOtam5uGtJIIWooI8z7rAKJl8nGQKBd07WWqwf/i0ZRRksokuFTGjNkrPRtVNSYlqhhjmQ2ECawMDCmDmSeZo1lN8ZY8WSh0j5VshzONah1G/AoOLeffsP+Oi/77yRyf3RvNmffPTlc75+cfGwkaNXr1hK3dxEIG4IgSUL581965UXnk1/qLawiETCyKVZOuak08+ErHjlX08+duMPv3OZLalnn779x0084KDUkwH/cUlVI8j/iqWfs26oX91xz997SZlvuPZbF5129gXfPPzo408eWDx0+LqSVcioMZ1x7jcuWbNqxbIfXfXNr0G2/Oelfz3541/ddmfZls1YsjRJQ0eMHnvH3554bumiBZ9998KvnlwrD3z/rf+8/MAzr077xhXfufa+P/72V6kXTJwy9dAFcz91rSu+cu6Fl15/8x/+8rrc/7Zf/vj7p5113oU85+SvnHPBs/948N4ONYg52UjASGC/koAhLPar5jaVNRIwEjAS6PQS0Fr+aDyjRQhAC+AOaMMmBW0pQDnAIzZEIIhs6GdKZlPPdQB4rG8QA2zmM24GdrUk0hSr9O01YKqtH7CYQJOcDRbuREiAE4BgbOQgMdhskQCjAMvQ/MYNFvXFfy/nIAM2erjtgXRgkwIZAdgJoLFKMnEwIG+QGxrbkCFsCompQLmQJWSFDuqqyQoDfCQbIPWjBVdG9DE0/M6T/OMMl2myIsNPqrcA2t/JUg09glbkhS2eHuu2+LofVO7Ji1m26l1kV38p5vUWfZLdF9Cy3al2u5cBQa+EDhHAvSLeQ8WrstV8Z4qaXoPxgqgXS+8rDJZaBbEKQb5Qemyeqn35xQvzx91wxdqaqbmJ2pUS6+JVnxMvkTMBSHFNw9iyxbJiR/sLYwD5FUvGKgV3Woe1s6J/kPNwLUFfd8d3BldQ9HHuDwiIJjygfiqZlPooCJA/SYb0g1gqF/mNjDrBcZJnF/m3FgtZocdl43VZnnrVN7iuNmxnrRcrjE31iVxQVcZmY2pQWf/zcd6hY47v/l7teO+iIyyfjaun1NQUiW2nAFJOgyz7s+TpknEpRX8keLqObdHxO+6/V2gwGQCZ+Zh5mT6h3X7RP+mnzLU7khg7f5TMujYpmTPdhzk93cKINe0nkgGtWfcg8yGnAP1iosHfqgVUV3QZJESFJxjwBXKCvqxYPNFDBT05iYQnEI0miiT+TZ7Psctt2/KKYHI8jtomrAUuZVCEYJ3ENZSzB60s9LsA7y60PxMv30+UzFzIWnyoZJgYvhP/iHcFgFfWflzBAf4ywfNuBMnLmg5AWiHtD4nBnJxxPu6K7S91NamTSCDNqoK5inWN2FCQbq6ihSTW639Ifk8yaxXvnO1SjmkjBoUtz+c+vEvzXss7M+ssChbsCYol8+48Qc5jrYe4YP5sVzog6Q5q7icfscY2S/OSlggA9KmExVXX/fSXAQlU8dff/+aGdMsLbqJjWEQjEcZtkyRenAp+cdtdf8Na4qaffO9bkBWckCXmGqLH0sSytP+g4qG4fcLlVCIejx9/2plfg+z40bcvOued1156DosGCIuevfv2Sycs+g0sHrLos09n6vLhuuqab551Snp5uMetdz/4BC6jfnDF178KWcE5cz758H2IirdffRFXnY2pT/8Bg3jegrkP/HX4qLHjf/67O++DrPjZ9664kGfN+/QT1i7Vd8BA9ncmGQkYCRgJtCgBQ1iYzmEkYCRgJGAk0JkkoDfbqa6JACQBSNmM4DqFDT6gPccA4gF30IpmgwIgCdjE5p3j2pXN3qijBigAGwAxIS3IemNFmTiOGxeIBc4jUS9ACXzTU2dkwm9YT0BycF+ANDYM1BnAEoAD8AI5cC9AjLck42IGzTZMu7kv3yFC2CBxH2SktbGNRvZ2+bcnITv6Ge0H+AW4SD+lfflfJ7TZ0Ij+TOiDMwUEvyb95hudvuf6E+PHHWJ/8sKkxNxD/Z5Ed583MWlNsLd3k59m7niCrMhJRFSdeERZ1TBarUqMVovqwA2+SBJEWnX3laupwelqbd1wFYhH1Tpf071jWaBH94cGXX7B7z6/XkwCPIOkJ6J1BwAAeAYptily5XZrnraIiwyED3Kir9LvsEQBdE9PgA+ZhAAYQmEpQyaQjvZhDHEeFhvErGiJrOCZ10sGTCHTllGRT+2HVScOKg4tiwpZgUZ9E8Kim2+bGpU9XyUcf27Q0+AVsqJifXjo38rivX4g5zZaroRVqNsaZ9CkhZ5xw3p6SwW52ao8juiDxwRMCbjjcVcknqfdCUFUQmZSF0ChvTkH7oq67al7IEMAZG3FxrxKH+ITOcL2MYiYi7VrwkxlAwh7J3kO9wRk5hjjhLn+ecmAzfRtAsRCakKIQIIwfzCXa2uOTPd/InmQe+HuA7/vENqAWDxnv7C4GFncw6qpi1g+r7dAPEDli0v07nHbGeLYKlsM0IrE5CLf8vvWiIuobZal8rwez9ZozE7EE4mgEBd6/aN9dpRwzdQ2GY8JmaDXfhQWsMKDrNCa3rgLpM1Y3yHJLmrhxlxLSnUFg3LGLySjsAC5QT/lvYH3ALOet7uFzIm7SALamoHboYSAJQB9nfHGO+gdknFj2C6SYgfLxL15/2d+1EoLzL28u0BgUKZxQlzgGnWtEBdtBryefNChbiwtwPlMZVopVg24i5oghMVLzzz+MOdgzfDV8y+6nCDdH7z7JvN8syQeoVyXUEJYNFOqIlB3YY+eva67/PyvQBJwHkGuh48eO2HG9Gm82zem0eMnubGTPnj3jdeISfHDX9x6xxv//tdTkBUcJ1h3S7KsrqzY1qf/wDatBb/2jcuuGjVu4uTbb/zJteWlWxrdm0Kk3P+n3/46/f4TDpjqvi8t+mz2rJv+dN8jG9aUrPr1j6+5UhMjUkx3v6OJj5bKZ44bCRgJGAkYwsL0ASMBIwEjASOBziYBbWWhA+mx+UDrGS1ENheQFmze2XBo0BMtak1iACQD1mm3SHujftqdCOssGWCSTzYe1EUHDwcAY5MH0IDWLObtbGLQcAJwQBsMIApZsKmgbmz4ALgAjtH+BdAFpND+79kcopXPpgJQjPsDrONaimsgQZAb5QF4a7eWm5xr0heb4GIRBoAhAc/xz+xuPiVBFgFIPiL5A5+KzzvD/9qSOYnJ67c6PfsmHN+UqPJzbWNaYw8euzIxpKjSKui9Ppiv1kp8CSE4WpV1UDyc4PZkYKxU9YpXStTluMqxw2qDv4cq9XRX/qilPomPU4saprikRaZUZ+eqPlnrlCOIX8ATURM2z1OvZeGV6YuUF69VW4O9Vf/wxosCdmNMZyx7dMBnSJk6IS60m5V4W+RF8u4AbMiO8QCoC6HWxDpB/p8hGTD2RxnKf4kcQ1salwOpG34dswIgGBAQrWUstFpKXO8G45XMOIqvDQ/3vVj2TWtrtN+olQ1jcrfFeqFV3ySNyl6gCv1lqsi3VQ0OrRghlhiDNtcN+eDdii+v3Wj3a8L8iJXFsKX2COWLx9WJvndUgVVpWQHXv357EvE66FuMb+YVZNZaYk7AWgTXWQQIRX4tal63pwBd+ZxkkHvmSMBi+gzzbIlkAJWjJF8pWWsItyYKyHPmYoAy1h8sIbgHbUfcCeZdbfVCf4VgZm0D0ANg5vna2o7+Rp9lXWspoTFMZgzQvpyL9RxWBK25V2mtDvvEbwI2WlU1YZcEEG8o3cRNS2EsoYoCPtUzXB8vclQiW4K6ZluW1+sTk4tYLJEts2k/n9fKFjdvcUvZW4XQoL0qxMoitjusLKRfaTc1kF46TtXX5TtzHGsz2ufHJP/fUblDpt2XcjHAKAQWVhr0OfpXe+L87OjzzXVGAloCjEcUEADPeeGAOGdeItC0VgbgPbYZWdGG9US7JJzhHtrijPeKxTJnoNxA+dg7sPayXxggx+fJtRB/LabJUw89gkDWCz+bjSV3swRoj5XCxAMPbrQQ/f71v/otBMPdt/36Zy3dGOsLfkt3CYWrqPMu+dZ3p7/zxqvapRLn4VYJN1O4iEq956hxE1gH1KyPpk876+uXXEmw7Ttu+vkP9TniGcolJKoqtrEHaJI++WDa21+VINiDhgwbkSkoNydDglzxvR/+DOuMZx578J72NAjkDXKB5Bg1dsLki888/rDUWB1YhXCflp7ZnmeYc4wEjAT2DwkYwmL/aGdTSyMBIwEjgX1RAmxsAO0B19n0A9YBxuDzHXCfl30+Ae8B8dmg8xIMKARgAwAEMNQgWj1uPLw9JARNVgBWQTBoABVglv85jt9qNnhoc6MBDmBFPSAwuB6Ag7oAfAJCURcdbFxvuqg79UMOAOTcD3ACGXEu5A4bMQAtiAoIHM7XFhWuWwzJyNjeg/KRx+3TifbUG/Nz5DtBkNkU6/SSfEHDek6uVfv+z4O3VVwXuFv9NHzLtiX2qLnL7eHx1XZxcboEHo5c1rtBFOGGeOdKY9NcmVP3RI3qEa9WwyIbVdTjV/VWUOUmGlS2KA1n2xEVsmMqz0moGdFDVdAXVw0x7c2m6f3yfZVqat774kWlQR2Y94HyC2FRHhJcFmcKKWlF7nD1au/T5Bm16oCquVgH8CtBq8mAswDjAGT0Q3eMCnlBBWKtEBf0VcA2+iJ9lxgO6WQFcsTPNWP/KslYqqSm0+UfXDQAPJIZ39ryBaJCj4ftfrCaJ8i8RyQzBhhvjMva6ya9EOv775XeingR4HPRlmh/3Elp7Wb3LoX+UpHZhyrHW60KxNLCa8WJdxG0cuzjvh5/rPyV2rMTSxMjeb6bpM3V7ZEfqov8/1R5Vo06wfeuDNCMmDL9hvp+KBlXP4zRNyQjT8oH4IDcLpd8Q8ZabT+I5RUWK2hY0j7zBECtE7cwu1OztZXidL6fkkRF6twM0UNmTqYv0e6XtrPkaJgSU4VYQnyiicuczn3oX1rjnf5JBrDm2SRtjaPXM8A0iGqAaADu1sg2rsfFFOPwLsmQFu9JxsKmS7Y1ZEV5ZX0wEokHxGqim89n9Y8pZ6jlVUUSbHto3GcXiBcosaVwEuJEpdDr9wUisYRwGHaO8LvE414jDcL+l/cEFAe0S8Rkc+z8R5KsYP5gnQe8RQGB+YDvzHes57sj0WfJWPEwd9IPmUf2C6ub3SHQ/fGeKe6deF9lHomlEwIp5yAi5kxAcxQ3dF9nHXta8kOSozsT8HpXtIE8n3eNdVJuSD1IFW31PEyOlcvvGedLXC0NGzlm3NxZH38AadFSWYhjccX3fvzzHLlArCDGn3D6V8/5+P1332zJKoP76KDb6RYWx558+ldxCfXUw/fdrZ9HsGtiQLz87D8fnfXR+9NSyzFq7MTJBLaurCgvu+yaH1z/2P1//kPplk0oQblp8NARo7BsWLdmNQoZTdILTz32EITFOd+8/Nt//M3PMymGqONOOeMsYnjwOy6n2tMeEyYfdMiGtSWrLrrqf/73GQkEvmjenO1Bh5Jp5JjxrkvcZZ8vgNg3yUjASMBIoEUJGMLCdA4jASMBI4FOIoFkDAQNaFAqDWSk+qZuBroL0NxJarBLi6HBR26qrSrQMAYoBlIFhEczlf8BeAD0SiQDAoEEsrHgdzQMtRXBniAsUtsPgFFr7gIyUlbQYzJgKeeyDgNm8Z0NEwRFqhYuWmHUYaxkABA0fbknAAQaupA3aIqh+YVbHTaYEBwcAxSDvACU4Rl6o4GMGoORG6JCpNH+RDsBItO3MDfQbADtBLBIewbEOuJzcctUnq9qKs7xPe8Cl7eEbhy51enx5WWJkbWfOFOX3BG+bnSN05RM+DB+uBroLHCDPXutLzAmnxAQRYlq1TeyTXV3aqTxvSpLXDj1dbuRPFR+x8LCK4hcRHDt9RImYV2sWC2LjFCb4gybpmlAsESNyF6khmd9rrqLlUCOFy5LOprEu5iYO1PNr8Wbw/a0OHe0m4fUr1aja5asyEmI/6gvEiDFI5IhDP8qGSAOiwUAVLTFM7lboP8yNujTkA5YSmRKBGKECOJ8APj0xLgGKAEU1P6wNegLkQT4DKmSKXHfJyUzfnCnwpxSAVnByUJW0DCAL8SDwJd8kzQguDpc5N8SCgnZA1lBor26+SosK6e+x+3OT9SZ1S82e+5Ce6w61P7EddXVLVpVoeqdRdJj1lshmbf8rmWO3rzzHW1U+hNzG0Qj8wNzGHJ9Knku7osgLlqKqUCAcYhcwCPahXvu9ylJVtBXmFPRPqVP4yqEvoYsiUfT1h6JhieWCu0DOAwAhjYx8y5zuGvVIiRR6rqT+r0JiCxlYj5hINK+3IPfmb+xqKE/65gWJfK9OK0RGYd/lwxArZ/tkoZp5+3z/24qrfFYHsufcJxcRzmyXgphEbcnizuoHh5l5zVEE6FoLFEvXtdsjxfLMe+IrIDfcWx7Yyxh14o7KDG6cKRtHUhI152kWFlYu8rKIun+iUkXbWs+6V9YedFf6FvpsUl2R5ucTb0kQ1zRjxqSMS7iaf1xdzzb3LNrSID5kb7LnMT7duN8lRZcm7UFpQDWWpRveL+EPMUKE4WZTuWSUIiJcik/igEo/DA+t7/8tJCIS4G2U0vxK/Rl8+fMmiFu6TxYY3z7B/93I8f/evtNrSkVqJYsLA47+viTysu2bpnxwXtvQ1x867qf/uLCK7573ccS9Jt4FulFxcKCmBAnffms84hx8Y+/3Y3rrcY0bNSYcRAa0QzBvedL/I05Mz+afra4fHrwrt/fInG7m2nLfOW8Cy+FrHn5X/98tD1dG8uSMRMmTcEyg/vd8/vf4LauSRohhEVDfX3d+gwkSnueYc4xEjAS2H8k0NbL+P4jCVNTIwEjASOBvS8BwFBe9vXczKcGlrW2sAY8uqT2ZFoTaNdQmnDgZ4B4Nk6AOmyoQGzZdACMcj6APcQAcuQ35Kc1WfdUC9OOlAVgGwAX7W3KSj0gVwAs+A2QVwcJZ9NHeXHfUpy8jk0ifnc5n+vQlARg1f5o0eRlQwj4y7WcA3jL/8gD4AqNbOqPzLTLHrcPyR5sf+hDVHVXJmRLWzEe2czT10gA28h3sbiAKiuyypeIFv3K20M/711obWNjfLRXxSf0ssoOER8lap3TR/Xzr1NLo2D2XyS/FVObowNUlrdOhawGaThbjVq/Vpzq16hIwq+6l1aroqzaDdm5EY8/Gt/gy7VXez12vmU71WJEtDDiDY5Yb/cP3xe9qs9W1XPqtPjRzVzZDPKuVednPaEG+EtUJJBQcVE5xviIuBe9/BvVhJxZQlwUKnGL1KRsQXEHVePLC2cn6lcKIZOu9c24/J1kSDTICtfySSwtcBcVTVpaaIIOsgct4+9JxuVOpgTaT5/F/RvAL3Mh7o2OTBWXfMf/OxYIet5knDE+mAfSyQrGE+31NmWSDMAMIMwzGC8uICOxNrgX5ed35plmqY9n81M+0eDOVpGJEa93qnbfBXlh4FX1xAAAIABJREFUBWwVz46o78bvUffUf7fJtQsS41WZt6jy/ZLD3j2h9J1PgrnReitHFTpZaomnm4DNQRc8YXymgjw2IKMAjjpBtqApyXxAn0PmAAktkRZoTQKYXiX3cC2BjKWF20eKJbN2QPogS75fJhm3UG0lXPfdLJn5FWAYUpg+BLnsksM7CAzT9lxPv4S0YJ5BW/42yZArxG+6uJXCYcVHveg/rB30DW3p0VadOv3vQix4tpbX+nNzglkySvJEyWNQNObkSJyKUDiCGyhpA8eS+cLJE0EGhPYNiJVFKOC3InbCg3nF5nDcDnm9djQhw1QqzHzO+gpp0WLMByEz2iWbJFnBnMsFuPViXuQ5TSf61u8Gacl6DmtMv6Jv8p5AP9UEK25mIFUhI1uywLlAfuN9AEUG7vewZIj1PaG40S55mZM6nwRSyAitINPoB5LSpvyuyV3efYgBxXrJOs176cuSSyS3OKb2Zs2T1h6MqZZNWZMFnHTQIa4LxtYsJfh9gRAWfF77s5tuGzF63IT33nz1pXSrgvQ6B0NB1yVULM1yY8ohR3xp4dzZM7/1/Z/cgIUCwbnv/9Pvfv3g3b+/RdzfNSG6uxV0L8RN1NLPF3x20VXf+99H7r3zduJp6GdBHuDuqaU4Gpx33x233vi3p1959/xLrrrmgbtuZ11rTFiMHHzk0cd/Mv29tyu3lWd8H0qvlxikTMStFcfvlXtLfG7WxSaJc1YsWbRABxPfm/3BPNtIwEigc0vAEBadu31M6YwEjAT2AwkkLSsAydgAaL/HfPLCp933uJtqyfplNdU0uStvQLVbKNYrXsLZeAMI4PoCeQDqsEECoASgR1MaEILrOJ/NFrLc02Yo2tJCl4v/0XakTLirAbRlQwggQV0ANcigxIC5gBO4hEILFCCMzSDtDADM/5AT3AfNWkgLyA8dnJxNGH2JPsIxZKf7EURFV+4vUtXdlmhDNpjIno0b7USsEBJjdZG4+bmjr2ezR1xABb7uf+aofKsaixmA88OEEFhlyx1yrFo13LtUTbJmq7JET1VtF6iYs52DahAIfGHtQW78ivG+z9RxC2arnMoGIRb80ZzukTe6Z9Uu9dfHN3vj4vAkZK33OTagZKH08GCDlbXyncSxzpvxEw78yD70Oxvsflj1NEvjPYvUhPhydYA1Rzl1CfVa/hfWFGIh4May6NewrhlhMb3oyPoe0bL6E0vfKstKNLQEkgFeENsC+bwgmU38e0JcbFSvFUS6nVZJv0RmAKstkRVokzOu2eTSl5nzcJHzX8mphAV1w7XDtixPfVCIHk+fwHrtaopypCfICoD+vyTvzRiDIKwTy4pUNwfa6gkw8DzJTYiS7lblc96od3ZRrMYZHV+dOzt7WCOaSbs5Xlstze6nJsfEoCGNsIjLUHwgeoV9Ru4r1YfUzNwWKC2vdyrURrGwmO1kqwrx7hVrB5nA+GVcM7fRJ7Go+q1kwGxca2VKyO1WyQQEDwuwurUdz2nhVvvu4aSrHmSGOwosKiCmIJQZKwRvyThm5DjzNmswfQHrFuZygGXagd8aY4TsIFGRKlRtUamBQldDXjJ9lPkfyyDKTnunJ8gWXERhOcA45Nz0GC8ZLuv8h7CCkFJadQ3RLI/PU5gb9BfIIu8PR6OF4XC8mxhU5HgtbyhhJ3rKifkeSxhflUiI5YU/nrBiYm3hEceQeT5LDU14PBC9YnDhxpFBkSC8sxYWSasd+ghzPmT2JMlu4Nk2EuQX7zAoN+AKjnrSt74kGRdSaySXSIZwZV6EhMKtDe8PvEc0N+Xa/kDmQkgTMqQs19+PJc/+OPbbagTzexMJ0Hd4L+XFRL9Pp5IVvFPzfoo7TKwkOYd5kbUTazP6a7tcB3V2uU+YcvChkAS4fGqtrGJIsG3NqhXLICtwv3TPH275ZVt10xYW8Vi80RKuqGfvPgMkvgP5yGNPPPX1fz/31H133HKjGEhANjZLI8dOYJ5REAv95KKnH/0blq6NaVDxsBFYOrTmegkXUxAu51921f88fM+fbovHY43lmXLI4UcRtPuT6dO+UJloo2LjJ28PuE3Mi+f++XC6K0/VvahHT+o57Y1XcftpkpGAkYCRQKsSMISF6SBGAkYCRgJ7XwIaTNdkhXZrwiYAQATwgY0Dmf8BwQG6ATRiScJD12KfdRnVgmsr3v0Bg5AJ2sHUmxd0gEzAG2QGOcH/aMgiMzQKOR8QWWtO70mQnvZkw0dbQaLQTpQHMAPigfYD5KKslBswigCFgGUQMhAQnE+ZqRvns1kBcADE5b5oUwNYcH9kgGw4zv2os9ZmB+xysyEqRAo7l7TmPRrOAFIXpd5OYhN8fIH/2c3DPKuOOMP3WraQFX3EQsJ1DYL1gthE9K/3hNRafy+1NlAQ6eWsCvZJrFUN4SwVE+sJ0qboQGlwjzo5/pKaOnOJ8kgkWV9NvFYU8b/vybf+6y+PhTzVdp01QJVbEYm6Xei2rTtv/Dj828S/YmdBcG0Wl0O1cp9mlkVDPCWLr/L/fcwwwe1722UqEI2p42o+U59mj1TV3mzlEwuPuJAnUYeu2TS93ev4hqATmXFg5exl/RMbjmlDlIAduC4AzCCOAr6s502snh+anz/xm/L9hBauL5Hj9GXGPOCctgLSIC5jIx1UvlBcWj2Q562i0BAVuPPBNUV6goAAGGQcQWxCXmxJIyv0NYwhxi2ATJPU29oyaaKzuOG88FtDtvrzj+gt1ihbfOCG2xOkBZxgfqBCnRt6Jvxs+DxXi1Kn9ap/oXdbPK9mU+7Q7jXla+T07cIWssJ3XYfiDmjZUJdnJTOnoIGN5UomH/mQGVgEvCf53wJculqYuwBgTxdRxv/TfJ67a96e9GueElybsYslBcQZwH9bLnrelXNukQwQzfrzumT6J/LXGddPuyvRDwH/6L+MCYAzQCCeiOsVV5M1JbH20CGpI8FuWTNWdYEYJq4FajgSD8ls2jMWSRQJCSFxKpweMcfO9zhOFNIiGk8E4nFb+b1eeTeSED/ipE28Zvol3kVQ3iXCjsfKlc8xHjlgO4l1cg5t6hNCBBlnfE9It7BIsXbSYqdsrNPMe4xnZN4eC0bmo9/TPpIhJ7iOxYCyEJ+H8UybM+8xXsmAibzjQLZAln4smX6sLS91mVI/UW6gP+AKZynlN6RFJjGZY0kJ8J6KUgGELoSZk+YGivdP1nZIXvok8xFkLu+yvMM29v1dEVB7b7UKrqDGTz7wYKwXUq0WWirPwrmffjJ46PCRb73ywrPLFy9k7m01BQJB5gyVShD07tvPtZR89bmn/vGX3990w+YNYmLbSpJ4GewdFOTGEw/d+2fcLKWejjso/l+8YN6c1u7zjwf+8sfb7330maOOP/n0aW+80kiCjps0xVXI+HTG9Pfaqo/+ffwBB7paMFhrZIp5oUmWJQtbL1N7n2fOMxIwEujaEjCERdduX1M7IwEjgU4kgTRiQZdMa+IDMmDir93NsFEAuCOzEWUjjCYo4AXHuI6NgbbM4H5NXP50oqrvbFHY/LBJ1xru1BvQEnAWkB7QlnOQETLU/t6RG/Lh/z2VXFBFMqAFmz7dPrQZmznKqQEJyo12NBtDXEew0UAjHTCMTYJud4AJQAu0zLVLIoBHtHwBXUnUEZBVu8bimO4PxqpiB1pfXAOlXkU7oqEPEK6D8wIgcow2CY3wrLCFEBh6vG9aqJdn61YhK2iTQbayKiKeQPcqb06wypOjPg8NVqW+bsHCRJkalb1AVQngXZ/4It60BHlWK7eOU6tz187t37Dhib7rltKm0+y51hbLayfsKpXw/6J5ENXQ85do4uoTAc3RqD26aQXsbXVO9tNr7EHOFO/cn2U50aBXbjMysl4irnvUykBftSbQW2IxSNBuLzxY0+T1x2u7+8o+/bDoiFVnb3z+BJ8TP1fO+Hay7zUB5VOuZIx+L+IJ9nq19+kPhj2h8VK2swTSZ37LlBjbQyQvkAz5pgFExg+baDTjAUkak9xv9KDQyv5CtoyT+06S/zORFY/IBWgvY8HEHAoAWC9kRRP3CtLmjN/u0nZHiWzOiCUxQLlnXO7tvjMf6/vv8G/6nxyea9cL0GCpEZENqtKbqyJWU7xwWaifSuSG62VkNpPNzKypw4bmr4qcX/P0DAlmTrs1dJCsSBUBdWA+QAPSrZdkAPZM6Qo5SLuhHfuY5I0CXmLVsScJXcrF83a51VsGIFnLgPUVYoK+dbJkLHOIMdBaor9g1fOqZABl5mrt+om5lfLvMrm1QXjYUje9DlIG7SrqPfmO/3iINT5TE/PSJZKZryBd/iv3qJDnNOnzbcigM/2MvHMkfnY3Kxrv7fV5uod83hxx8RSMR+MBMZfwb3cTZWULi8H3HIl1IUS9zJder3CziXwZaJZYXCSk5fr6LKtUftwm72XajRzzAjJusU1b6V+UjXc35ikIxEslt9a/AHmxrGC9J/4O63hJUti8J/C+Qzlo51SXPJSPZ/HJewJKG7dLxtKS9Yb3BuJXZEooekyRzHsDVlbhvTDuWyiaOdwZJJBCSrBuM8dBjDUGb072Pay4UEY4RjJ7EuZIYi6x9jRamlGffZmsoPyQD8SQmD3jw/fb0z4E5j7xy189994/3npje873i+kDGlmpbpHEwxOWn+o/Lz37ZFtkBedh0cHngMFDhz39yP1YjzZJBAznQFvkwHti7VArvpu+dMIpX04lLAYNGe5aq25Yu4b33XYlAm5zrzdeeg6rm2Zp5OhxbsDtxQs+a5VEadfDzElGAkYCXV4ChrDo8k1sKmgkYCTQySWgNeGZj9G20VYVvPjznayj5rIZZgPLRhYNWn4DvGDDzafWrGl1093J5ZGpeNQ31bwcNFXHhUBOAH7ID/c4eoMP2ox8uBbrgvZoO+4K0WirCAAHgENABA3OUU4AWdoJ39KUmTal3FjR4NaJPoAmL21Ku1Nu6ssnx6g3GxoASoAMwCfAD+0yRD9LlwOyYlfUa3+/B0KEVcCqBc1sdxOoU0hFtk7xfjbmQv9T3m5WZVTiWAwVgDvbtqwJDSo4u9yT37/GmzWqzM4Pl/nys9HCJ07FyOyFKuF41foIOOoX6TnPhU6Fp0/lN6r+OW9SbOn6aI5v06DD1ze6gQud1qw5KB99gz4zSZ59VYYGu3+bU7j1n7EL3hJ3VbOljBfKOfUBJ37FsMhGCdyNw6KEWi2GGf2Da1S2t7YJkVJhFw2eXnzYAW8VnvR53/CmlUeVT2d84boE0Az3NFg2NEuQIXW+nJO2BbrnH1oxY8O6rIEVDd6sTIQF7mvQAGYTi0up1DHLdzQN35TchLCQup4p+UOJ/4EbgibtklIYwBTcWDHG0BitFbIiEzDpybHqCuR+J9Y72RcLcVEtlir5kBXi7itxbfAvXrGeUUXWNje+SL6QFkMim1VI4nu8nQcW+EUSrFQFvA2F+d7KWHWioAmbIVYmo0fVLF00tvrz8sMqPqZPtZnaAWgDlAKsEESc+QT3TxAT6Ym14xeSIUCZW2oEvEzsBfASrV1N2ANu7dQc3QKYzJyL7JlvAeEgKtBgdd1otJKIw8IaQp9jvuYe9CHm9VSrnzbbbTecoAl62o6yYXFBgPhMCU1XMm4UZ1J+kVP1XmjrXSIGn89jeSU8vc/n9QoJkZ9wVA8Jrt1HxmeeI7EqxMWTeGy3EgGfNy4N75Hfg3KswbETlkxrWX6xs5D1sEa8Q3kEJOwlhlDECtGWaDsTeFtbd9E/mIMvbaXCN8hv9HssdXgfcMegZE0kpc5LmYKma2sz3i9KJFMHyA/mVNxFQV5kGvcU6VHJD0jGMmdt0upmXyWwdkmfMjdpJgHeQSH2ed9krdQKP8yB9LFfJ3+n37Ke4npulczfe1IxaI80m7YuaCt+hS7MS08//vCM9999a8O69oH7xJcQp3VNXGflC2PB/WIS5bo9lRyeJCz+/ezjj2QKmD1M2AHIgy2bNjBPtJhi8sDP5835VN9Pn4j7JgJuZ7p3ppvhmqp4+MjRb7783NNcl+kcAm7jZmvlsiVYkJlkJGAkYCTQqgQMYWE6iJGAkYCRQOeQAJtQ5mQ2zwCjaOuhEQrwBAivrQkAUbAi0MA0wDWbXY5pX9daA2+nAKDOIRY3ODRFsUURSVsMIJMSyWyoUkkBAHwNLnGRtmiw5Fqsu3eZNmwrsnEJkmSbIX82eK7GVLKsaOTrwNtsDDVwhgsP2pD2hcTgWurDJoOMBiYbRvoCG0VIDs7hfECN1E3PnqhnKyLokj8he+SKJQxgEG3imu5nWQ3VR3o/qjzR944lwbZF597JEjA7GFW+9WErIDu2wMTPg4O8q7L6SiRe8buUTJAWud5qleejOzdNApJbn2UfYB3sm1Va5fl47eA/bI6ECL2bOdHXuS+IOUGoj085jQ2hC+LLPRdIXvxJYmqJuK8CaMCCISDlWJtjh/9vVGR9qEe8Wo22NqgyXz81KmuBmlvbVEm4KlF4Xn63imU/OeyWFR+/8iXIBfot42wW95J8bYa6qGpffvcaX/6pq7OHKCErMtUCebK5BXgDJE73f61JS2JO8LzUm/hF3qdGnWAwYIUn6ADYKQ+B/IBYQVuUOldnIitwGbQgcWRogT1O3RK5vv8qZwgya3St1MezxXuu73kJhh6WQRh3g5T7RFm7IFGrRH6C+HuWfpw9dkDYE2B8i6VKwiV+BoRK4p/XTW5CWIQS4fDmUJ9g3ONjftCkZubWbf9R5gPtyuoJ+U7bQyKdmuEWrDW46bpUMtYsuAxivmlx7uiIy6MkEdFel0/0X79cw7wZ34VuovS4gKiCqIAIg2y8uhWR0k+QG4MSuaABXyKZvqk18NvfIrvvTL3O8ATKd69kAt3i7grt3nQS7GtyjLphabE4aWnRKdcJcc2USWruS4CwDXFZx+OiklwficU98YRTKBRENOD3VssaXy9qCaGcoM8rJ9oSvEK4WNfXni/g99RbysP4qBDCo0TetDZGokLUWVa5hLOnbXfGWkaTblh4Euga90zpCSKB9R3CFVdPvKcwz7F+u66o2hpfLRBy+j0BLXgINQiQWyXDgGNNhfVmekI7nvcO5uoSue+WfZXAylA3c2gnJIBFhMzDWC/Tp9lb8C5KYj6BiGMeZU3ESof+ixUaCgusyV0ujZt04FQsILCcaE/lcO3UXrKC+3mFsUiNX8Gx+rrtAbMJtN3WM9nUaAuKZx598J5M5+MSatWyJbw3NUlcV7Z18yZib+gfhMf1SBWakKTSESxiWLjkSvwLcoVjuH76bNYM+kBjEpLnIMo14/1pb7VU/hEScJuYHJFwQ5fsN221m/ndSMBIoGMSMIRFx+RlzjYSMBIwEtjVEtCgARtrAHgAaTaxgNkAXwDcbEox++U7G10ALjYLfKJVDRDBZllr3gO2AFxpn8ydEpjYAUFqAoYXeuSAfCB3kBl1ZiPFyzfAFy/d2s/4Djxqpy9B5rQpbcLGA2CSMlFeys3/tDEgGptCNoSUF2KCa6gL56MFDdBKAhAGmGAzSf33dh13Wkid9QZp7qDoX1i9HC+C72Upe74A5Flij+ASFr2trSvEHVSDxK5A6/5EAcxDcce7WsIUFG3xdy8r9+YHl2cPOFA6RDNTF8D14XUrSkerRZ4lapwmtlyxlAV6HPO7EdcPvHXkz5apv7bkQck9FZITMIzEPEBZddLjAV/p1KNEMtr0cQGqQAaZP8JSjmoB348pTFSfyVmH2bNVaXYPtbJhjBLrgMabRZxg/xxPzWHh7Kx3JID2iqrXCogHwX1JAKWAcf+U3BgEI2F51dZgL7Ugb7yaXtQ8zrY8u8LrJB6LWz76OuVjfKeTrYwn5jSIOgAS1w0CSeJXbKqMF07ZFusRkKDb6VJmLoXqwfoAAFrHdGmsE19EFt56J6t3oVUxcbJ3/gAhKgC5m6SjvB+4ZEUvq1RlSzxfTYx4pA0lVwkdOkfcbIXDKgBBJLF9JY6Ft1Lcfs1XK+rH1Auh0khWVfoLCqb1OPa0qRWzPj6wcs4sr4CwNz8+Lb1/NJm30/3op5cv5X9tdYWbDuqOdn1T84/tJzMvQVrcLPl+ybid21WBUtsLAGttcc53+4wAZjtLWmg5sp4yFrAwoP64dWqNrEAW9F8sEQDr6IOAwIAqAMqdcR2lrSGwsQhhHAIqtmSxc5P8BnmFK7Dnpc+XdtI6be+dzZPj8VjxeELMmsSzk3QWv99n1Usoii1iZdFNMLIeXqEqoomEEwsnHIJtW8oKCEGRwMoinohBeOSKm6g8YlxI7AvtOjK1D7b07JaO09dYq1kLeD9rEtco5SJco5RIZoytlsy8pONrteuZ7bCw4v2B+ZF4Nox5gq3jKgziIj0xJiBXXkiWozlr3q5SmZO6kgRk7uVdAktF3lF5Z2AtxjoNJQ3mlmMl09+ZSyFImS+7LOg8ZsLkA1evWLq4cls5Sg+7PAHsp1tYrF29EnJTYekw/Z03cEfopv4DBw+58Mprrvvwvbde/3DaW//hWJ/+AwZl5+Tkzp898+NVy5uTEpAKg4YMG4G7p/TCP/Tc6++vWLJowbfOO/1YSJmph3/p2AMPOeJLD/31jt+mnkvg7EOOOvaEA6YeduSnH2+PY8F9b7/v0WeOOOaEUw4b2Scn1aXV2IkHuIStPjf9uRAfQ0eOHvvpR9On7XKBmhsaCRgJdEkJGMKiSzarqZSRgJHAPiQBNrw65gEanACPANlsPgEb2RwASKD1ySZXazhhccGmget1gGnOhchgQwywDRBOUO6uFHAZEAlQDTIg1dyY44CnbLwB4gAjXM3JPWRZkd7lAEG0Wyh+A4xjzaXsaJNDQgBg0l5oQQI0cA6akZSdtgPcoM3pH9SFulFPTci4rr/2Uv3S69tV/9da2vQp2bg7fnEZtFwg6sm1jk+cpNdvO8n3duVxvvcGD7VWA2L7xZgnVhHNHbjIN7jbpmDR6Ors7IGZyIpeWyoafLFEzI74XyjwluON6fJ0IYo7Jdx7fCQESkta+JSPsjEfACh8Q3Iq8I2rGIBMDfTXhc8Wj0ecdILrHgZgln7FXLPJ59ib8hP1V/f1lKphntWq0F/ahLAgvsa47LkHehP2AZf2+MvG4IMuceaC3JEr3T6LBjH1OE8yfXmCuMXCskQNrWe6ap7O2Pzyw+KO6rNPCw6am5VoaJh38SEZLcNEBjwHkI+5sJGwiDmBQpF7MGzLcGpGCbma5wSl5bpYeswKqT9ji3HYJ6G8Ry21R/brZlVVJJQHS5om6UDvXBnQPiXWKSLQRi8qaBHOE6JqZZ7dUDUwuvX16lDW5ULSHM3Ffk9EDQyuzBqe/bn6vI6p+4skBE32krxxA97qferbAxJhbsicpq3jUjXouagjYLm2RoGkAZDk3sRtOD9jA2wPxotbD65jDm0x+HAL1zc5rN08dcDFE+3NXMn86FoyYW2xE5YWzKOshZB3EE9jJOPipDGQaFo9APt5NkARAB1y0LFA9gX3irqvoEXLPEBbMv4yJUymALN5PwD0yuRyqD3NvNvOaYGYc8TyQiwqbAlb4RGLCk9YWIiwxLGok9gV+WIlERYri4ZYImGJayiPaApbXsvx+D1WPV9tW+XJQJcA3Eq4C6enkBXLJUdlsCG7HbWeoc9AMhM3AvAfF3uZEvMiwC6u2rDwauLnfxcLkvpoF5E8h0DeELWN82XK866U725MNJkH50Fi7+KymNvtQQk8dFkTZQC9r+BTYz2uBdsVD09vbS1BgQGSl76Acg17EWJWsH4yn9K37pTMmsr7aZd1J8bGgeDQr73wNNaKuy2JZ6QmMixZuXwpAbIv+fb3f7R5w7q1YoRQf/RJp33ltLPOu7C+rq72xaf/8XddmCHDR7G2qWceeyCjdQUxOCAXMhEu/33rtX9/5dwLL73/qZffEcOJ2CFHHH38RjF7ePxvf/ljamX//a9/PnrORVdc/es/3vvwX2+/6QaCj1989fd/NOXgw4964M+3/SaVrOA6CAtcUGFBkUlog4cMH0mw8QapzG4TqrmxkYCRQJeSgCEsulRzmsoYCRgJ7KMS0OA2L3Bo6QE6sEGAeOA7oKUOQAvwyAsugAMatABraFTynTkdc26yC9BJ5t64U+pKgZepvwZp0O6i3m49JWu3HXxvr5bv7ug2PJ+yQTZpjWdU1WkXCAtIJspMewPsskEEPNV+qQHudIB1gAc2io3tmbyWcncEyNwd9exy90yzrqAPsYkvEFAc0POYLNUwU0iLRK24DDrQO2eTWFYERnmWRQJWtNSOWxvicW/fjf6iKVtyu3er9wf7+KMJrxATkYasIJt/N/lj8diIpeselmO9Nmf3+WhTTn+f34kdErP86TEYAJ1bAxXpMxAVxHWgf6VD9oDx+Lh/RDJuoJpsjpMa1lEBrLBaKJM6FoScyON94uXn5yfC/k3RZri9zCOJcYfmTD95vPr8o3vfFhDwC81z+jxz2BuSAX/xLf/TKl/B4dOLvqQeHXhJs74ytXKWOm/jsxcH7Gjxz5fdWtcnsrkq90q1TYiQTKQFfR0ZNqlD1A4Gs7z1uG9ScYm16/dEtfUDYD1zIxqiAPGNCfdP8o8GtgG1h8RU4OBKJ7/Qp2LnrbOb13u8Z5EwPIEqkRHjEg3U70hmjo7JKKwNOtGNErS8h2N5AChdwkK7/ZqQO6sZYUEBJJ5HwUsDL+x2sB3mfjp+EW2q5wLqqkmMjrr4Q16sG5BIzDmQU99t1gjb+w/asvi1x68+QMPOgqoeIR2cVNKijQCs8aRLKOpNfXdk7tbgHG7KCBRKXVkbcJOERnmmRB+hr+p+i5wg7zqd1nAbGvYO8QiSbc04J39Z8qgMlUZbGk1pgnC7AZ73FUsLsYyIi5WEagjHfR6v5Qs43sqgBNROOE6R5Jh0AIlu4RG3UU5IgDRHyXdxDdUgv4nFk4qKNcY6j+WUe5RnRdhJrJZTtAu1NsdWmktfuhBBAAAgAElEQVQm+imkGGAuhLC2cMvUxxhb9CuUD3Z2XLXQjZsc1u+TvCNC0r0imffIt9MuxhKDtYF3yiBxbOSzyftEW26q2lMYc84elYCe78bKU2l/SAbWKd4nmRP+JMTGGvmMphMXSaKZtZI+ynrJusC40HMnawmukVjfXbdFXTn17tt/ANYLM6a37NpoZ+sPaB+NiFFmWvrDr6//wV8ee+61W+9+yCVLIAmee+KRvz141+9vKS/dAlHkpqys7GzcVb3+78zBrXv07kN7qsUL5zULbv2HX13/gwGDiodiWQHB8NoLzzzBc9NjVSyYM2vGY/ff9YeLhUC55a4HH+d+kCh3/fbG6x++50+3pZed+BXlpVt5b82YxOuUGzOoYjdZrexsm5jrjQSMBDqfBAxh0fnaxJTISMBIYP+SgAbeAbl4cdUvemwe2WTqmAyHyncAJzYbnMsGGE1j/TsgExsLNtCAEAB7fHIfXhCx+hVl5z0Sx2FPtGCq5isy1IEzUwG+vQXma/KEMmpXCwCSaO0CbgBA0z6QGXznPP7X59NubBq1Wy/qlh6nAhnvrfrtifbda88QC4TGZyfJi6Jcq3aAaOD3lgDZniGeNX23Oj0KRMs+YjuetWM9i9f2szb1thrsyuq6rMKqSE64plvWwOrC7EGRQMDfvaImnPB6qxqyXM1mlVddv6RHWdWyhuxgTlZ9ZHn/LeXzq0cU9pBzcEWTSlgwpjWhBaFAf0hNGqCl77igUwtCA4QGlKW/ZewzAkzZ+LWX35+Rm364xBl5T1YicccQ36rDlkTBPr5IM6qPV8cUTj9kQnzVsOXB/gJsbADAV0IycG9ymVhbAM7llweKImWBoute6vOVU3ALlZomVs9Xv1h6s+oWr+oxoGH92fK50m+DOarFcj3gSjx5T/cyaRe74MVNpXHHPyvu+Bq1mYOeBhn8CQle7lMV8R6qyL9F/DG5ysKPSmZOxJppqWQXlExaVfD+S3sAbAPMnCtE1EleZQfui+HivWma7J2n1jkD1DBr1eKY8s8MqggAkLbo2irXVfaNbQtHLH/MVhZjFe11N3ZESMrXzVuh+gbWKQig7Wg8bqRkQgj1Htm/Pnzoxqw+9YJ44naCw7Qj5aO8tLn7XTTMNWHZrHzbD6Do3SxxDw1wcG9ALFxApSe0aol9ol18LZHvO6p9z3OY59oEgdMKoedNl3QDQGvJyiKDP3+ugQSG/C2WTKwK3PQAJENgtJSQB2ODsUc/aVeg01butzd/0oQhlha4AKFud7RQoOvkOJYlAJBY+e1oW+/J+rpKANGYzMQea4vH4+VdqH/CFvMksWqT95uY5VFhec1RQmyIigae2mxbmIoqCcIdjMUTXnkLQnujWrxGwWc0SGae0oAhVhzN6pPB4oO+xvjHMlIrIUAYZ0rMA1g4MLfulOXSDgia50GoMhb5PELyrySfmOwXDyXrAajNuczj+0I/2AFR7BeX6JhouAH7arJNJ6bV/AT5HzeBd0tmD5GaNAnHvABjz3wMeastfiEqms0VbRDR+6zgCVL9vUvOOV27X9odFbnnDzf/QuYx7VKz8REE+T710LGDCfodrq+vW7zwszkN8plehnf+8+/nyS2VbeYH771z1rEHjdmwprm1g3AUlVecc+rRBNWGpEiNT5F+vz/dfMOPX/nXk4+NHDdhcm11dRXl4/pMz/2/ay7/emsBulcs/XzhBaccecDa1Stc11cmGQkYCRgJtCUBQ1i0JSHzu5GAkYCRwO6XgAYRmZMhI9gEsyGGsNAugACU2EQAZgNO6iCuAHtsODHfRquXTzYYZMByNKEAcnjZbUi6h+ookLT7JbBjT0BuWhNXW1Rwpz0NDGQqvS4bBIp2m0Pbac1uNN8Bx/hNB00HnKRdydq/dqP7py5ENu1Ya++dq0I+FR8qYPZRtSp3iFhR1K+0h/audXKDQlgsOtz78aeTnXnb/JFoVjTuy9+aKOi11VtgJeo9S4WswCJDVXTPY/yRVTASrZMesKU+J7Qouy48QywtVgTjkZI6T06luH8i9gPueXRCExot8fmSCXLp+tJPEwNa+fQlgOZ0cIJTAae5r+smRLuDyiRKtKwFCIbUiPZNlBdvdvrfV2ytmbJEjW1ChNQlctXqRPG4bf7ZP+ulwj98debBi08/eGYTqwchGuJC9lQPq1u58viyd59YkTP8SLkvc1NjOn/D02pk3bKIWGEE8yXYt8+OA6QBGmMVgebveiEuYqnWFmNz5oTXhEesrI4XbBBrB4gGASC9CldVGyODVDffNm1igosENOvfkQwKWU+gbWJVyHfIQ8YhhMVVkgdIGQ6Py08VMvVK+zYTT0hwUCEpNvS1Nq8WcoSNNqDOSsmuixetoX7nvADjGXlh1XAqxIRP+IsCX7nqJwG4txMWovjNSRKwuyrY64hNTnxzodwzVzS/BVHNQxNcGpl2LhJAFXdf2mqMMrcaGLtZwbcfoG0gwmlbwGzIb7TvUxO/nSaZ5yI35iCA1h0BMPWalW7t00LxmhzWpFdHr+V85I7fLe5BO9DnWkqQ/5BYxH96TzJr6o7Itj112tPnME8QvwCiCpnQ3pkA9Ufk+A2SH0rGs+jU7l2EOIBQoIzi1klFxdCiVIiJ4u2midY28Tonc7IE15YfLI/T3++1JNC2lXCUE/f7OK5icn6tXLw5FneiMrb0eHKtHrh/OxuK6xjCnA8J8NOU65hnGUsAvcQMgTCDWGEc7Q35Ih7GI/MI5WJehKTSY5txDpPMPAaxx+eOjPl2is6ctqslkHQFRZ/kPeAayfiGgrgl0fZamYf/eSf5ieRBct23xMpCB9XmN9ZnCHzuw9pK/2b+YL1jDeUdpMkY6apkBcJAw+uDd998bVe3V+r91qxaoePTNXtMlZggfPTe2yib7HCiDiUrlqF80GKqKC9DkarNtFziXZDbOnHlssUo0rWali6az/uTSUYCRgJGAu2SgCEs2iUmc5KRgJGAkcDOS4CNdIbEO6UGt/mZkwCr0bRm06EtMHBLw+YDgJKNJWALm2HtYuAM+Y51BZtiHbwZ8IaNs/ZR7+7tXU1Ey9rnSIuW5JeUERsMLT8+2ws+7HzDJu+QoXxuGaRcAGEarOBTkxIabOZ32kYTTTpmha5DqjXJLiuvuVHrEhDAnXboGbIiR0ZU6LCoE8DSYpME284OWQ1rD/HOevUUz5ubPFvia+rqAtFwt2DPbU5e79UD+k4IB13gujH5JOJr3Of159SG19geK+xJJD6I+73vlvUsiJ1x9cxE6PkAIBH+5QEFXCA+mSAttcuz9AJrcJf+gQWGq9GfkgCoHpPsWitgodBWmyctLeq32L22fBI/pLrS6f5fueak9OvWOAPVB9njTzohPOssiU+x5s55Z9VCCOjzRHbMY1krc4ZNKskuPlRiOjQhKzhvTrcpamTt8uABVXOVBN0GyMf13QOSSyQTe4IgyJshLeTTvvd7Z1krGj7KGZq11C/xIColu3IS4kJVxburj6qOVyOyFzHwmRsBXQClCRyqyQrkSDkgf9G+L5YMOH8o7qTEJZQSQkJ8fyG2pkliVCwc7130ksS3+NSv4rhXANgDGLZT3emIDGyRBZqHAB085zqPTLX5vgo1ILhazas5QvlFA9wnpcyROodkSrd8OQN9qn6014n6BQX1Cdq6SXzuhz2WCkiA9xIBWJkbkCdEi54bmrVlG+5bCLJOn2T+uVUymt9/Takl6wvpdMmACcS8gEClX3XUt70GdLlfR6/VRXLXxHQriwyWFannUwf6BHFbWorhoM8HCHpfMkFN6Se4RWpzfKTIqzN/RXY6VhIugT6VzHvApRkKDaEJoDVNZEu/bVEGnck9ELEoYhI4WzpapbiGKrfEgs2OO3FvQAVlgOTKcSsWw6CUly4rLm7i1/l8jCuxrojbK23HRlMcEs+1DpPUXjLBndckozzCGDknTaZMHryXMbaIWaGtJqt2d/9qpX1cyxtpX9oZ8gRrC9xZMZegHMO8yDsl4LV2PZmhq5hDnU0CKWQFbmAho76WUkbWp39IBkBmPcQ9ELFWIKjox8yTrO860SeYP1kbsfZjXsTV7BYhJnZ0Hu9sIjPlMRIwEjASMBLYxyRgCIt9rMFMcY0EjAS6pAQ0YcHGEnAOggGwiIxbBzYPbDhwEYM1BUQEoDcAJyAUx9hwshklCCQbUsBvwDjmeYAINKXYaLsbaAHR91Yw6t3WgEnCYI8TFe2sEHKnLbT5d6rVhbYO0VqYAAmNwJGxrGinhHfhaUnA3TvEU9K73smemiX+ngQ83jzUs7q2p1W2scQevP54z7TVo8LLsqObrEFb83oeXervXl2TleXbVpjPxp/sJguzJq/XG2qIfiLBqt+1HGue7fV+KgRG7IyvNVom6IDqrtuotMTY1xZVqT8BOgC0cQ2WGV+SnEp+EuiVMa+tkNolIQD4f/2nqGKT3WdmvcomvkMzwmJtZJg6XFyi5yXqr4xbnmdz7PBKAcTiKeA9fRgAeZiQFU19QSVLUevLK8tO1PXITdQKi9oEJ8XVyo2SIVoI7olsIAh8hb7S/hE7a9KUvI8CqUGsG2ywfNiNAdU9/Zvmi0sogBaAWpdIkbLpsQcBBLHL3PkDLRBxMqNqnFy1zB6h3o83V8yvU7nPfhA/4pkx3iVbj/B+7LZVS37/5XlxIS2Yi5+TjGXN1TTAgMBasVVZrDaER8jTHJUlREaODPMeHmk/x3eI1+PEREW8m2iEDxbuFe34etv2RCRi8DpxYxMW7XDAVUjOmGiDdxhcT1rQQGazjjD/vCv5uAyd4udJubOOAFoh+2b+7TNcpw9RXXKqZm8rp2//KYO2bnvmcv0sxgj9jL7TEllBPRgTWCM9JRkyC4C2xbZss9Cd9wT6B+8AWAEBXP5e8rmStw+UpgliEEsuyA3au7MT5FhHbJZg2tsJfkcCaltqq+1RfvHzlCfuoarEbdQ26TxhsbDoKdNvd4l74ZeJuEbG1Sb5v1yicm+2VUIHwLY7YF3B+g2oizUSIDHzY2oC7CXxPnaIZABhyKL2EiIZmmfXHJLxn5B5kHdKiAvWBchbSBuO6cDjmsDZNQ81d9kTEuDdHhJakxVvyXc097GywtUdY5rMXMk88O1kfxwjhMeHYmWhyQj6KQQ1PiBZt+gL9O+DhTjGfRSEFnsJHVtNW++483RXtrbYE41onmEkYCRgJGAkkFkChrAwPcNIwEjASGDvS0BrSmtNezaQaEWhxccxNpZ6U8HGFyAQf+OANGxINDgI+II/E/y2s6kmo0nIPXB5oWMiAFpEk5r/MBftAYb2vpT20RIk5YshjQ6srf1Fa+sZaqZJitRj+2iNd0+xkxY06TfXZkupn6myJNh8h8Hd5EO84iqoT0QFuzU4oTyJXSCIV15+nqotq0wUrKuvCAX828L5DdFQz60F3YtlhJbIk7bkV9WVR0KB7GjAF5TB5WGABSOxN7pV1d4thMXiyu65NQUVtZUrh/dPLRfgG6b5AAIQkKkJkIxxzztbqrsO+gpERrHks5IXMMY1ScGYbwIqtLdlzjn1xcSwF2+tkADU64NWpCLiBJvEAVheP15tiAxRq7wrB02JLr0lbPl/LPfeAiCWBPJpD+Yp5p4xzRvNSfSIln7SO7JlvMStGIybpJTkus+ShCsrAsPeW58dWijus2yJBzFErCly8rxVI/oF17puoFKTxLBYKxYXq8RiY1auqt98XM1cde3bLllLWSCRzpZ8vmRiHDQmLCwqnO5qXqK5V60iq3xpqd3D/8fotepY339rjzz54/aAj7QTrjTEYkZgU/kL4hrKU61KhZwJyZSbJ7hwN2mebI8a7PX6rGDQU5Wt7KCog8u87i0RmWyV71YsbmVFo3HaFRAKwiIhrnHqd5C0IFYJgD1rxaPJT0B+wNXUBKFDsGBAWRL9sr2uYujX9Dtva3Eo0p7X5r8txK2g/6MlXiyZda+RhMpwQyxjsCxBCQBCC633rrz2aUsLQGnkhF97wMz0xPxyv2TmHwhCCA5IuU4nmxS3UBJ/wk4IaSFRtWVYWba4flIVXrHk8vusAnG6li2kRq6TcOodj9UghEWVxK2oEtJiudhcbJLrKuQ6QPpmZEULVjzMZ8wjKIRA4B4tubnvuO2Sxdc/cy/uU5BjKpGbQfx77lDSyoN6R6SelI167ej6uOcKbp7UmgSY/1ItK9g7MJ4hKVjQiiVPk8y6NUQy6zFWiMwJfYW0oP3ra0sW1OQWT2CdwUoI4g1XcqxhkyTj+oznoETAGNBECHsUiJEKmeuZR3QMIOZ/1gvux3HeXbT1dyP5bUgOkYpJRgJGAkYCRgKtSsAQFqaDGAkYCRgJdA4JaNKCTwBXQAPIBl7u0Wxi80FCQxjCgfMAr9gssGlgg8FmgQ0omqZsOlxwK/k/mxM0qAAeOcbGg894V7S26BxN2qwUqZqryF6D7JzYlQKi7wnxa81qDbgwZnSwXx3Y3B1T9O/keOkoOZe3we4/RtwBeQqsyjIhLIZucvoG+zkbK75a81LPgys+yfZtjUVqCgvDFYV5vupuOVPkOTNzahsWSYyKAfKwgYJLh33x+HO+WPwPtblZy+tys1z3Rlcd9p90kEi7cMkECuNihLroemn5Ul/ITOYKnVItLAAfAaZT+1m722aD3Q+yYU7AiqCJnwqIuPcgNsOi0GA1yN502oBYKXE20CaeIRnyhXIAlBLLATKjSZJ4FQt7RstmdYtXfyDkwjHyI+5VMiXcXL0ooGN44NqtZfFin2d8zqfHrgkPd2NBpKZcb014RcOYqhxvTUmvwMalP43cHx0QK4OkwC83VhUA8xAWTcgKIaWk42xvjtfiJ6scqy5W5+Q0WrRIQO0Xy53CCnlc5O/RS2TcXttCUb84nOIaapZyrL+LVc3led4aNSy0TMUivVVDoqcqtBLiKspShR6v8ltiWeGxhmb5/flij5MQTfCQPK9XOEo08cRg22sJyO6pjSdstMIBTuNCWkR3kLTA4oQ+A4hFxSEr0gkLKkN8D8BXAK51co3rWqylyqe5pNHrWZuy2sET6NPsYXBzclDy+zdauReu0XCPAlHBeqoDLe/g4/eZy7SlBe0BUQVpwzyVKSE/vS4xd2DZ2enA7BTSAksLAUQdf8J2rS2EF455hKygrjJenV4y8zOfrkvYNu9DK+Rzg9fjqYlE4xzvCCGj/frzbgUhTGoyjySP0c9wZwcgzPtYuLOSYrvbRdU+M0L2/YLSj1PnM+Y45nesI4gHBeEwWjJ7B1xCwfK/I/mu5DHWkzXL/n599ZSbXn1PvjPmIeMYM6zrWORgUcT7B5Z5xMGAHMZSjzmDzDoxKvk71+HakjmEPQxrhnEpJUIwyUjASMBIwEig4xIwhEXHZWauMBIwEjAS2KUS0K6MUmIwsDFgAzJXMpsRtIOLJQNWoWWLBjIbZ631yuabY2wktOk3mlFsVthoo1UFycFGBKsLNP/cuK/J+xut/l3aoplvlsFlVUcAkz1Qwk7/CE1SUFD6L4QcxxgrOi4Ix+n3gO3aZ7/e0ItnHQdiqD0gHPcRdsHnk+DabuBj2/F4s1R9ff+GjZuHb1u+qW/pxk2xOm9/u9DKquye1zsS9Ac8tt1dgLKQuHsaKq6gqoSwmB/3+WbF/D5c/LjkCmB2BklrqxCALkDY1HS4/AMgkBogk981EUGAap0gJbXbF0iA1N861MAS80Jia1RuTji+pwXQP1WsEJhLvnhQvKfqHVivKjz5oSHO5hvEo/w4j3JiAmx/OqRmi3ez0xuNzKslA5Q0SRJg/P4Z3Q957aubXijtFdlKLAFc1wCMH5tyomuRJDE/bhOZZg9cs+WeLX0Ks+LZtQfm+ypVD/9msfIY3Hh6bSIvVG9nT/ZbsXu718caBvjKIGeZJyE9mAOZH3Gn1yQJYSHK1h7fVqenI1YWyLSJ+60ypygsdUdjmv7UkTEbcxLBWaLVTf/8ul/ZWX19W1Q8e6laWddD9ZA38FDQpwRtlRKIRCxV5/d7CrJCAfEKJYfj9oi4YyfiCac02yu1kq8NYbVOSIs1cj9kg6VFR4IFN9Y76R4KSwP6FYG4aSPInNRULP+gkf93yfRLQC5NoqeLsfF/0Zp1RNt2dxMW7F9Yy9AgZrxTdqxC0hMgPaQZpBv1BIRH4709c0CLdeyMP0AYtWAdQFsAntPef5GMz7PLM9QBWd6UPA9y79+SIR07naxSSAvA0YZYPOEXqwksBrwyx/NeJMPaiotlRYMM6GphAOu9lqdGqMBqiWeRkOvbay2kiTHmDtYE1hUIZObk9MT88DvJuM9xrWW7Yj/rjH1/Py8T6xXjVSesK3j/550i3WUZ59BPITQYA6zRkAscs2Xurpe5mzWBxPsV7z7MrxCdzP0oSOg9Bs8skczaSsw91nD2J9rSm/0FYwXLLZ7FnE1Z22OhmCyC+TASMBIwEjAS+H/23gPOsuOu862Tbuq+nWampyf3SBpFy5JlZEtYtuWAI2axCTYYYxtM2F1Y9j3Y9wDzHvCeAcPyFu/iJS3BZk0y4ABeg41tZBxkW8jKWZoZTQ6du28+4f2+t2+17vR0T0/oGbVmqj6f6nv73HPqVP0rnFO/3z9c6hJwhMWlPgJc+50EnATWmgSsOw023QBd1mKC72yC0WJiY85LPxsSAD5AOUDKUWWuI9ijdR3FpgFgh/X+PmU2+Gw6cDvDJgUABy30hoBct5FYa6PhEqrPKVw+dVsIABox7iHoANCZE2T+x1UBv1mijvENgM/mHNCOTTOu0E4nfgv3RDt/RPENShPZ4GzONPemiVc8EG9pvL76qacnR4oN07s+fuKqrTfVinlt3rOZnrnGdDMftUECP0n/p2JVPCAtX9wnUJfGMmQFp1M/QAEspm5f1O3fp//xuY+Ge3dCFiD23UEXsLYiQZAw1wEIzgVwbKj9e0VYANifAH5g5aB4EearRQWVzirhtfW93xNlydceS6/c3TQR6xG+sK2rqu5636O4FnNfG7xl+h+HX1d/wfS97aC/yl9RRhPUEjZhEvhhMxeV4ig0tVL+Fyo9BXVwYoai4yJLwFlOTFnmZ0fr24ZfUvjgFbKI+ZbItJAlayZapkumhsn9/e70sr/6YPPfCvI171l8ksgK2k2/NETinDZh0bGymA5qhUcy3/xB5qc/Facl05DHJ1lUmH4vNi053s/lfKNmlvoLWZILg0oxF/Qq0PbWlmfKJREaAlrlESsqVmrNdVGUPDUzW2uItGj36Rn43j+p7R2f9qz/zI+f7MgJ4Kk7MZd+RvljyvTpx5UR/CmfFQK+EkgLyIvl5H4Oxxn3gGWMe8AyNN1ft0x5EBWQLgB4EH4E1z4fdTqH5qzepacIvIxVDUDjp5RZiyDzuucm44A1FEsk5grkIe8SgJesI2tOZh3Som2xRr/K2sKO5TbBrCpPQQV6vsElVKtBlO4O0beUxJcge3iWANoiFwg91tr/0JHN4iIAaX9QmWcQ3wFpz2XdXb1B4Uq62CXA/MQNVPfajVXhUok5/Wll3C0Sr4I1YVpxLFivzT3Qlc/M9bbrMGWu2aPMOxFrL2sI6wfvFswPLLasBThzj3Ih1CErIO/svOM9bc2tIxf74HDtcxJwEnASeK5LwBEWz/UedPV3EnASuBglwAs+mwE2ymzI+c4mgA00WqQATJhq8z+m2YCT+OZGk5hNAVqRHAdUYuOMH1mAJzSgIDP4nY0GpAUbi7ZLGWJaCMl1ptsX44h67rXJWlNYgsK68GAusFlmMwwZNx94dZ6EY4zzHW1Y/gdkB8RirAM4MRfaQCtxsJeztLABt3UabhEAASa9NHtAsRZaTS+Xlzb8/lJpZsvUxp5NR3YO7Dw2PHitrClqyrP1Qm59GviJvn9an3eLrECrmflZF4B9Asir+3T3CnMe4AFygwQoDECMBqTV8u3e7HMMGQBM/ER3QZ3vrB0EnT7XgK/Ui1ge3W6n2re4a+ZlZmfhsTZ5cF9xp9nSGjNDycwL8qbxpVF/36DifPQJ7LdBaLur+I/6BwCk8f5dP5v93BPvp92fU6b/fkT5vcq3KlC5qfTkTb2YN4pfYQ5unQ+ngCsoxbIwOwpPmp3Fx8yeGnzEfFI9e+ey3t/Yl277oIKlT/d70wAuy5IVuIOqZcXfeHXl06GuY/3sThDDP6f8JWXW0JNksOj8k/6Np68xIxMPeI18bvf4uuJkKagO7pSFBUM4SDabgTAzvZAS+cBvmfjKKApyKZVStXzf1KMgbISlLMznApldREk+H4b1emtLlrXGRWqMy8ICbfGzBkY7lhZtMk2ZYNUAX0slLBggCRifzCvG4invK7LirOu1TB3smoDFIcQWz793KC8Hzv2WfvsfnX4DUJtbiqyQDLsJ0W6XalRjYc5Jzit195r+vdPXrAcQhKxLxIchEDfJKjDYNozqC+sK6xAuZrhuzYGNHcIO92iMNQgpxbbIbMwf1VfO1Z4ZhcyV01XKYEwwvlh0GF+40YHUOykeT0dgWFYgM54/WMI2L2ZibE0P9EuvcqzfBN3+QGe8WgnwzmQtGzjG/Piy8n9X/qZIihPc4q0QT8JazTGbeI8i2/WYvYi1SuRdi2cJBDFzbWH2uXgVl97AdC12EnAScBJYDQk4wmI1pOjKcBJwEnASWH0J8LLPZgNQloTWHoAZfmFBOu9WRsMcQJDNA5sEADaAHBungmNsIAAoABz4H+ANrVRrrk25FvCtnIHLnNVv8QUoUVqUgBm7BCYgE1xobNQHwVfrHQ1LgF4AMUgdEvJ8Am3kC1A9d4tnJGC1+SxhYTe+9A+/AZ6iic94ZsMOak2QSDblaMLyfgP5hpY/1wC2Qdjt7RyvY9GxDGnBPSmbsj6h3MylzThIkyuLfnVfTzSzp682s30qLAxMrOsbVuyBilxBzYmkuF+unwZUu6dkw8EmnjEEQXh8MVmxTEdDQACQQVadQNEAACAASURBVHBgFWUTbm2oezeZiAyYw7QTC6vFCYsFXDicMci+qCDkRn0AOk7y2a4A2G2Lh8mgbKaDkulPqj8g4H9GMR9Yawjyu1TCJR2y4Zys/w1TzK2p6U8P0I+AfR+S/P6xXsy9Wx00KgsL841brl0gLCgwkCgUp8JsDvdX95irTnBVpV4NZ7L+wafSy758Q3D/bXLptUw1zMG6yf/NHzff1atg6lfIkqRb5lyDhQ1jgfWWsXBGa0DjPcY7+vGP+41cLt63ffPDXpL/7ER/7Q1BmCtvLB02heYms74YmJIsLPImTYt+2J+LgjiVg6pcLghi3bpm4n55Mbt6tiKnNlmWj+N0WMG5H/D8aKZSba4KIdABshlbjDEII8BXZGp99Vv54QaHgMOMbYhxAN1VJ7hPEfSYZxlr88uUX6mMC6PlyIq/0m9/pMwzlOdi5VeO3GXe95ET4rlYooJ2MI+Qp43h0Hbf1slrDqhfbkCvdLxjVcOz7yPKgIzIkz4lWVdythgsWHAhhVu3+9QvNjbNkrc5hXXHStU65987pF0q4sKORwumLrgmOwNrJMYC4x+SmzWMZwvEN8+SpRLkj3W5hWxrjqw45y51BZy+BFinsHpgLXyTMgobrJU8T3l+4XKR5xcW1lhMPbSYrDidWy1BOHS7/bPPxkslNtDpiMyd4yTgJOAk4CSwChJwhMUqCNEV4STgJOAksMoSYCPAxtsGBwUwtBqEAOyjnQwgibruy5WxqABEsgkiAvCTjJY2Gs1swHEZw6YC9zIANYAUADpcC4CBy5zlgNxVbub5K07gCm1BhpA3yAywFaKmrWWv35EFoBfA9ID+t8SQNYFHixh3IhBCt+p35IgMrYUKwGooYOJ0fWGfv8Y+x0vuit1iW8K4tICTDazLxhtygk/mB2OYPkT+9AXgJYAzY51zAPmtz2Ssk+hHyqV/+Wy7SlrGPRTXo/VPXxMvYF0tLG7Op/WN/d7UNS/2vzQ8PZrbeXSk/+pGITeQ+r6Ihmxv5vljAtq5715l/L8zx+aWcwMl90LdPZfJ4oK20EbGXrdPagiJFyrjXoG20n7aQPuxCoCQ6U4f1T+Azmg5nrEbhkWWH22Nc60I47JsGNMnmtgL6eHqTea6nnuMiBzz9dLVphg/aHZnO1+qmBDHZF3BfFucsPpgvYFAPSHl/9C0Dvz8wNzQxCygyg9MDfTuVy4d3rxueP/2EzkZTzWCKBlOWBpPTncnL3jtd0affKvcQhWWISz+Xlf9P8fSjev+JbltWG1DrkslSDBcdTEWTgu4hqjQuW23ZRtnH9kW+7kXDVYOe897ytx4YMM15S++4iWm1xszWaoh7OVMPktMQdYkYRTWQnm+io3fFwSBgm9niaKixK3YK4ZhukPLcn8Y+Ed9338y8L3amGKxzFYYzueeOqQFheF6jLmFH/Sl0i/pIM8crGRIgGLncw1ckKXuw9hjnrOWs66/ZJk6AtAxxiAuv3G4dc3sH4//6eK+s4Qox5nvkIUcQwZ82jWGttGXK1qULFOXNXdYfd3U8wzwkucirr5wmfXrnXYuri/WScicdw362lpkrgpZttrC6SIlTmuuLro//WyJCsBfQF/6n1hA1k3d4irfqwOssZyHMgnvF2dz79UWhSvvEpCAiAfbypk/evdLf0X//JmytbrknYH5ynvrbytjLTWna9bk3L0Euss10UnAScBJwEngLCTgCIuzEJq7xEnAScBJ4AJIgE2vNalmEwx5AbkAaMn/1yuzhhNIFLLCBuHmd7T8ABcAJAB2CDoKEIo7KTQF2bhw3Gqi8xuAHeUD5FYFltVOMzjxBRDFyrcQAAPIBBkDCkwbukkKgGNreQKgDNALCMkxQG6Airs6d2GTZ4FvysQ/LxqUyBegjM0g92mTF7ovmuKAFWhh73ealSv31RJnIH/SYqKCOUB/InM0gQHyAYfQfAdYom8gFiCT0H5FsxCgHw1+XMAwfwBXceNB3zFfKINEn9G/WFoQiLsbZOI65huxC9YLzL5JRMTLFEg72RKKl8i38vvWb3xhXPA3+2n2Vbl96hVZQTBnyA1iHexWboMDp4hZ0anGCR/MQ4BEysCXvNV4Zowxb6m/BVMh2AASn/GH9ExRuC9hblOPBasA+ahua5SfYVwB5AL4yxz4mvK3d9d4f/0yMxWvk2ujcXNcxiUHwmEz0+i9fqt3aO+BNkd0UsJiBbKCMk8A9j5w35u9v5FW/+Dk7OyOvUc+emDrcGVyqPxexbFYqhxz04OPmKvrB0sKrj372wP/EcB5IT2e7towk/UlyibnNTWwFjAaAHnWw0xWFdO/13xP81+TF+6QdcVJ1iOdwgBqWRurpxO/okNWAHSyXtAHNwdZ/NZic2ZXzSsNKbCJWTczY8KhOSHjY6YnlzeDuVDkRRL6WVxI01w95/vBPF2X1eV7X2xFUPYCT55usv1yE3W81crCVhz3DZQLk6tFWHSJjucG7gVxf4M7paWE/xc6/h3KzBEYIwjB80VaQCYwv5mL9PFLlXnGvW3JQWHMT+n4XuX+OMvffzy+bPrOyjvpfOYO483OIS5nDaF8Ev1FW+lvjrHeME7pS65rSXvfxktY8tbPMZdRkFLIEV/2tJV14r8sI1PIK8j79ymzrrKG8rwDDL2YwHmeKzxDcE3HOwLtRGN9ObKC9nMOz5t/VmYuEGj7YpLJMkPCHT4fEhDpQLE2dgrvsRCo9hnOOrYwtrrIinZV9D/j8UmVwRrGOyzPH87n3WHPUlYVOpf1jXEPkeGsI85Hp7oynQScBJwEnATOSQKOsDgn8bmLnQScBJwEzqsE7OYEty5Wiw8Qko0FgAEADpsNgETAI8CEz3c2KQCZaF4D9uCLH9/jfOcakEQ25WyGyGzIARDZvLDRYePdEpDbWgTkntfGnmPhuC+hHf9OGbgPMAqZIAOICT4haUZNkKuZpIl1RduiRBlA8sbO/fkOgMNmD9AC8Ap5cS6/QVYAIHM/iCJAZvrpd5TZGPK/S0tIYImg2hZ8t6Co1XRmTNJfHEeekBKA81gMMEYZu4x/fsNtCS5qLKFEXwD20+dcQx/xrgP4T/8AfAL2A0Yyzq0mdXuudeJXQJJAgLxaWfMr25v36rViWO3f3L/nkJerz7VywaMaZXEStF0/AXYD6EM0oHl+NmQFtweQYB4yp7vds9BeiDbkRVusqzgAiqUAZdoCaUE7Z+682beub9qfBNc8FWmB5UeXlQVlYa11l6wr9uoTt0DUZyHNJn2mkRUU6CI2DxV2mFqzaOJGONp9Tuc75Cpuh/CJH3cTAJAVOsacvXlysPxiWVYcC1vJrMiKEyw6bJlDEzOmXK+awaN107eucgJZwTnHs/XBh1rvCHb4+xTcelqCaFsi3KOM9QlyaezLtiV/3nprYSrrVyQJj3VjcaJPGXO0f0V3UCIrrOUO68YblF+hPCZXYS/21WX5Vt30ViZN72zVNAZCuYKaM/35qslH/VqOMpl9tfpl2pZkJtdME4Vr9/1SMZ/ToBCbIQ9RSZwOZuJZNB4blVo8oPkE4Lzaif5mbhBcGyLiB5RxE7U4YUH008q4JmSdPSbyloDWZ629u8gVlLWsYKyxNkNaMha+W3kpyx3qh2UOwHrbEuBIfOX4Z2b+D3OkdTVrBmOLMvluXV0R54b5xDOAOc+aw2/0O7+x5tPvrD+c1w0cniSQZ/sA85o2ng4h2QHVWT9mJXfeL+hP2vdtyieQkp128bwkQzhiSYCcAepXx8TnWRReR9mBZw99z7qJsgPvTBA1du1cXEPeuVB6uEMZKwvmYuLIimexIy+eW1vLZ/uuwvOKd3fWJBRrWJerIhtOWGu7CAzWcBu7jndeFHYWrK91HWOaMnlP4j2Hd41jOv5ZldGez/pOHayFKmsmawPransNXEyWXDyidy1xEnAScBJwElhrEnCExVrrEVcfJwEngUtWAiIHlmo7vsvtxsQGGGbtZoPMpgKNQABMQBbIBsA7fgM0YzNiN+L8D6AP+MZGm43J48qAMtZvPoAu5wGYAgj7S2ifr6n+EdhAewGWX6cM2GBdASEbax1Bm2ZNzzUF45d6zeBLN5ugp2lyUsZvyg1PVL7STH3pmJn+VyGJT4922k5nsEGkfOvbHFlZoocy2ThaAPmX9H2f6gNg/TkBF8jZpZMlYAe51XRmA8yG2Lp6YjwDmCI/iCIIOruBZ9PNMUA1rIjoa4gKC0Ja8B5SicR8gGTCRQzzg036aKd8LDEoD7CVINyafm0rC8pgPtC/nD8QeMn0SG7/veVw+vr1+SO9fi6eFozFuOAcxh7zknsAbmNlcaaWFZ3qLridWeziiXH3m8rvVQYkhKih3ciSoOCL06/7Jqvl5XPop2u7zeHjm9ty2bShbDXMCaBpwdfsNABOgE3WCvoE0gGSaCH9/djbzU9u/SUTyZJhjzxGeVm/+deEqfdMkpVKPTDpnyguA4TFCXE1OmQFfQggjYrpdvXGE61ciDXESenaB/e0G943O2c2CL9/08CnzV3pi8xnfYbFM+kTre8w3x1+3Gz2DmmSxr+nfqQN9Ok9R7PhA6+pfMqfyIYYdxy3mvbdRQDKtmOQKC8JxHcsKiwQzpgaVQYAYq0F+NX9iKIt0cunU7k6bUaf3m3Gdm6TG6gxBQ9fbyJfPIWsSMLMLwR+1q/CxgPPb4SyrAh9P6k3Y4K41+M07ZVLqHIu8g+JyGj09QTJu77tqrMmCJaSbecY4wSQnr4GtH0r4l7i/P9PxyCACNQNcXGv1j/m5GpomVsCC3LCEoIAbEuRFcxtrEGYFxDN37in+papT8/8HFWmv8n0iSX6WMP5PoABi+Y+45o2M6cBqxmLfGdeY6HFb1zP/9aqYM1q0WNJdRpzeqE79ayK1W/IECKC9etvlXEhw/NvcSKmA9HHbZwnwFBLPC9x+to91CEqrBsoyArWVEs0QlgslxjvX1Rmbtj4Nqsx5teusFzNLqQErDtY3oN4p8WK583KKCG9S5l3FshZ3CvyLEXxYlIkg1WegZyF4GVss2axlrffuzoWFbxj4U4PZQ72AVzHXgG3Ulh48kzh3cYm1j4bJ29F4r7rOvfVScBJwEnAScBJ4Jwl4AiLcxahK8BJwEnASeC8SwBwhE0Emws2MVYz1PqCB2wA1GQTgvsbjqOJxWYGkAdQASCJa7s1ytm4WIsNADs2SmxwAGwhL9qWHWuJtBDIAJgLKEUGrGWjxcYM+aDtDlJqXf9Mmp6rN5vBV2YmGt5kcutD4wu7qj3ZMMVdJeMX4zaJ0TqemtIVnum5ttfM/Gtkxv9BDuW1R4srAFfWdc289nQ4NG7S+gaTVgHCkRXAJHKDBAIIA6R8g+oJ2AewAQD0NEG99XlJpo5lhSUTbF8x3pCvBXvZZAOKAvpazT7cngFiQzwAkvMdsAy3XSRAR8b995xCsFgdAa4BQEIqQHigTc18oL8AKymHucXcsNqJ6r/seapcKKD7ZfWsWN7gH0lK/lxP4MWjnTpBDGK59EnlPcoAA7NyA3W2YKadm4CkixPjmnkPsMZ5aE4u6cZIDoa2FH3z9Ru9RrB900Cx1oi9RqOVRkK7B/sKXO9LfZ/2ttstgDNdAeC08XO470la/fW0aB6q3GR2lR4yRxpbTRos5lvakL1iScQlxZOIGibnW+uKDllBu+h3AEPWq3+jDEh+kvWIgps3s9D/5q59+28ZimdNtCFRPmLeFX/EHGsOS128bBRse0F2v1b7T43RcM/hkcrR+wd6pu/sKYgx8M3B0dnHaTsyRGvUugljnbRkF2XcoYw1yKnmrgW3GWOvUmY84maHNRSgvJ1EOJgobZhyZWK8Pj2xu3826U0HzDUttaEpwiLwc5oINNeLotAvBl5AlO1mmqWtIMj0u1/OZ2ZG/RbreKOvtyCrC99X3/nqu/NBWlAmaxyV+k/KgLNLpe/VQWRJkGvmMoBXQ+sfQG6b6D1DrXPKQIaMB55PDCYsLH5jmftzmLnHeAZwf/iR+qshK6y1i11X+ASYo2xJzuuVfsAGdQvzQeCc1+iQlloTMsm4bZFBuxjvzGuehazzdt8EcHe28/wUTTn7nzpBcc+2ToxxnlmAocyLn1f+b8vUhvX4/1RmPf4tZcBMnpPnyy3Y2QtliSs7RAXjjLG1rtNe2gI4zDw+FVnxnzu/82znfQp5ORB3VXvo0i2sy3KB9Qz3Tqw/rFGMM9Yu3l94l+F9wCoR8Nxi3f3nzrm83xB7iTWMtZF1q0dlMa6xkLTWFYx15izlce73KbNms3bz7sWaZ62GWTvdOL90h6ZruZOAk4CTwLMmAUdYPGuidzd2EnAScBI4PQl0LC+wtOACtMLZULDZZgNh3VawCUH7GnCHzQqbEM5hU/JyZbSFITYA0kaVLQnChgTgk/MA7yzgwUbeEhzc82yBkNNr5ApnCWQAgIKcoG24+8FcHrAZjVjqCvECOYAcqqZw2Vaz7lV503O9yIfBfpEVqak+5huvLzT9LxHKudE38VhTWs9N03vzOlO4fKOIiNRsfHvOXPbLRVN/IjaTd8YKiiv5xiXjFVNT2D5r4vGyaR4dM6XLpEqe22aSatNM3VFX+OaCmfnaOhNPAXoAklOPlymjUf6o6o8LiYfPxWXKqgjyPBayjMsn7kjfkRlDALxskq1GM2MUDT4++Y33EkggYkKg5QcpxfgEJOM8S1ZQLmN/pfQOnQDg+FVlgDWAUMYNYKzVuKYc65+eOgDYockdymqgPhQe79mUO5DbUXhysi+cmpK2PK6F9iozX9DAxwUU19fPgaygHZawYKwARgDe2wSggEUPQAaypA24JjshBSY7WDDZ1dcEzftfm6sN5nNBvdZotcqlvBcEXu9ctZmGoS8S0viFfBgI9EbesYDvWjdpsSggOPdI5CaKtQILopPiB+xvXK44FhOmkpbN/tbJeJ+IilTume6vm8KBHd6+1hvnXUDRDuYJc+YtHRkyl2nrkqlUb3y4P195rH+o8jV9/5FwV9YTSBRX+E+abw//wfxO80dPuO4hc23+xxsf3PLr0z//tgPTW556aeXLR7c8st9/7bd8pviZ4ddCkFGPb1GmD7vd2+Dmxa5/J2iQd1w/ITeIFtYfSGKAHhtvBaCdGBBdKXtavVsNk1YrCPs+UfCGRqt+epUXNPwkE9br5U0IaZFFfmpi2VsE6iLRPJ6JFIA7llOvOVlcTCqQxax+2BOFimrheycROsvJ7SyP83yhz9G4516A1KNLlMX8wXUUmbHLXPvrzrW4imKeWFLlVM8RSEwbWwlzGcY/z63vP0X9qRtjkvnyDZEV8b/M/aglQ+16wrpBX8lqRY+AzEv0p0cV2SC5KvtZKlGnaSp5ey0d19esKPHzHYIUay5AQRLgIeOkbZl1saRO0HVASdqJ/CB0X6uMJvdSiXOYbK9X/kXlL6ifIf5wC/asviucqk86ZAXjlTHB2sN7BOAsc/Z2ZdwILpdw+wgxxzyHyFxwkXOxjAPXjrUlgU5cibrIBogylGF4/71Vmfd43mt4B3iFMu9LrJOs17yLMK55jvJs5b2ZT8Y26zDv84x5Pnmn4F3IKkMwL1iDmcOUzXv1hOqx4FJqbUnI1cZJwEnAScBJ4GKXgCMsLvYedu1zEnASuNgkwIbDAptsvK0PbjQEIR3QIr9B2WqEAgQDLpAhNADpIC4A4dicADJwLZsfgPbRTjmAu5zDph5tX3zmXDAgQsAC2u/UxW6gqDcazGysaBN1g7gBWLYuhGhHzax704DJD+ZN7w1Fk1s3YOLq4ybq22j6XlAy+a1FE5TUjrAqb98CtDJhvM26yW1XuYk2evj7T2SBsfOg6X3xkNzF583M3UdMftOASXVetmVGCrjb2wRIPOuZZNIzI99fNK3pG83ArZ6ZvjPR+X0iNh5XJF3agBk/1iBYv3xe7UITlQ0iYMdegTvU/WJKbdcDndQNSvMdoA9AGvCT8UmfotlrrS4AA3HthUYgLmYgoNAIRFb0NZvwM03ckwxRwfiwPurZjHNfqxUsJfjMK358mjkFhNlTzmbueXn+M3NbB5668fHmdTs25fY/JesKiBPrMo0yrOsagILV0EBEHoBhtHdx+gUdQOuZ9gAUkvcpA0Y01ZivRyY73OenUy8ptMY2RVmf5/k9wmEbkzM102qpelkWqdW5nmLOS9LUl9XFrLTNa4Vc2Ox2E7WUkG+9K6VOn1b+pU5eOK2a9Mi9UU3mWHlT9J8J4xKpK1taol4ffsb/ifzv9iieRLAj2Dvy6fhb5ibC8qbU+Fg0MBb4hOlgjp+UFDT7PkH4U1EuuWdn79Hpcq5xRajIE6SccJdR/2nzPP8h87bor0Va/NgJ1z8YPC/6ZPNNLwnj1nsuO/LUA7lc/XMbmsent9X2b6mEPd5kNPjjwqsZGwsWEfrOWglQ3Zr+NPik1s/3tNdaa1HBeGIs48IKwIhGszYxXpdKW4WGfy4Lch+P111z32BwzXo/TVpeGLzTePVSkPVoXY981UPdFNc9LyIQvMilIFQ8i1mNsicD39unNs+IsKir72pxnHbPtWVue86HrcYtgbiZl5DfEBPLJQA1SEbmL0TjHcqQQfNE8vwcoeOoO2UzB5ErGYANMM7Gsnm3vhOzYrmESxTIijYZOZFsMyIszFi8k+u5H/egXAC4IZE/Mv8xg34kwDn1S6nJdiiouWg7T8HOTUECPyiLlgMiNHapgkVdrXU607OvTUjhYgXXKzwj289PBdk+4+dhJ87EUu05IzdOp5DJufxEe1hrcW1nSXdc3jHnGfdLJeYt1i9/ofy7yqmecbw7WOWHC0ZgLIqBsriudizQDghx1homNqQ4igW43FkufUU/kP9UGQCXseUsK85lpLlrz0gCIgzGRFp8RBex1mHVxnOHd0meW5AXfLK2svZahSbedXif4T0Bq02es6yxEBiMYcjJLyuzDnOM91LeuRjbzGFIijbRTDBwF7fijLrMnewk4CTgJOAksEoScITFKgnSFeMk4CTgJHABJQCwYIEfPtlgsElh48J3tL4B1NhssGGByEAjm9/Y5LQBHGXKYRNjXWVYkIdPLDSsmwdAJeGFWXK+SQuBDjyXXqkM2AWYYC1JqC/gLAQFxwDPMI/fqwwhcL0Jy0+YzT86JEuIHrl4Ck3jkIiGHTlTKq9TzArhpuvV1qhpogIbtVFl2qV25gAxBE5G3BtZSY7F0ETrcTH1lNxI9cl91A5T358YP1ynOBhSfo4bxu/NmaRfBEjBM+H0VpOr9pmwMGf6XnTETH7lGlO5t25a4D4LMUbQWIWgAFADmD6k9tJXX8CPOCc+xxOgUHdGrsgYmfJJmwGKkDMbY8Yn4wwQFEAQlyScy5jmHPylY1EBMHy2iT4ESOZegKjMB8YQ8wUy7ATSonMTv5jVDgx7R67d1tqfNWZLgz1xvdAwinsSeRVdAWFBnSApIC3Y6MfnaF1h20fbGSMADPiY7k6AtwRDRjYQO7fbHzWgcoGXvVQC//DmIH56m2n253OhyIpsYy70h1sKHjFTabSiyJ/L56OG4iLU6/X4cJJmc709ud6klGuKxIAI4f5LEi+yusDKgnXEkhYLdXuqdk07TgPBt/fXn7GwgKwgDQSTpj839sNZrvWip+WJJ/X8PQqQs1WQOwAK1gy49WozA4tTkKX7RuKJQ9ubx45vaY2X+7zqq4Ncypyn/9qpV91yRfCkmWgsWYR5vLgreMn4V7+n6ee+ZzI3ULtt/CsviNKW/8lN33mjSAIsthaSyKqD/fH03e/a9+HZd+7/sF076W+Aa/6nzjSMtZO11Mb0OBX5+Jdelv56GuSb5Zl9PSW/NFOLyvc3suO7G+nE9fJzFRSzAWHoYUW+s4ysYSQacUpZVtN3rdNezvd1v6wdDQPbijgf+atBkC0l8sXHuA8g/eeVWXtxP0KACNbkpRJzGm1fFj/mGesAzyPmmnWjY+NG2HUccI3rGPN7lSHhSBwDOFsMmFMu5PwXlQGRswdrrxdh8SpLzndbX4mXMFtlW3GFBmmUJtnlmK/IvdagLFU0YDKFEPGqrSQJdXy95F0IPFOTnKdEZLBuEOeCZyHrCMR++x7v+8hd2ZmSFh23TUvJ7IzJj6VFf85HqQfrABYWyJB+h4TDumY513uApVgUfYcyrhF5vn5dGaLqPj3jZvV8u1BjdSkB8Exi/NB/kN68WzDnUSZgnGGVulyChPkVZeY8az1j0QK5a6XPTlF999NFJAEbS+rX1Kb/qsz8xDKIuck7Ce/HKMawlvK/ff/iO2MeEpF19w5l1jPGMdairMn/3DnWbQ23IDpHVlxEo8g1xUnAScBJ4DkmAUdYPMc6zFXXScBJwEmgIwFLWnS72gAUYBPCpgNQhQ06wANEBZrkNggxQAKm4ABtbNoBXLnOag6iScrzASCC79ZdznkVvoAN/NazCcPVxN8rs8nif+qLJicuQthwUSfAMmumXhVZ8aS57FdfZebu2yvComx6rusxQX7CFK9smKBvtwmiF3faxGaOcpGNlRPtAzAHgGSTx/0AKCGAdpri5QAwmclv/qZJk10mmThsansj05ocUDQAERgDPcYb7zf5oWkTb/BM762bTc+upqnui82RDz9sqo/jmx+ghPLpN/qBewKAoDU/rLajiYq7iedcwjJBlbaZ/moTXMp204wsGVtsjDnG77gkoC/oRyyC0AwEDOZ/wE2ICjbj55os6I8lEWOIcQ/wTPloaDMO6HMLqFHPLT3JXGNdz7Hy8Wz9t/a1ZrZtMgd6RuJD+VKt/qV6TwTZAsgOYTElomI1fbczPpjTxMbAnVV3Ql6AgtyXMdVOCB5MW7SZUNm4+pp8ze/LmReJXBTYm13pBzJ6SE0oPzezcaw4CF5rumn8mUYrluFCJrdnJpmZbYjEwATDZPsOT6enAGKpH+sF5BJamQvpydoJ/y4cHwrGTUto+/25Xa8o5KdfQlPZfwAAIABJREFU0Z9UALIPRllcTDx/RITBv1vUzoV/Bc9nN9R3P3pF42B+Qzz9OpEJb1VAcfqIelhN/TZZMuo9bXKHGsf/Ln3zhl9a93+bR6JrTM2fj6dxx7rbzb19N5p6kDfXzD76n+/pv9F8boPMmyL4hhPTVZXHx/ws2XH97ANXba4fYhxbkhfXUcgdN0UwIz+lzLpi0wKBsqhIxhxk2TFPJiKyaDlmhkY3lMJa0Gy17paxRH8zm1HcikKEb6LI8+LIKzUU06JC8HSdjzPAZhwnrFfjYRA0Qs+v5mQVs5rxK7T+nCq1tEYBiLEuM59ZE4k1gt/zpdIbOwd/sPMJ0A/RgaUGgDjzHHdajHWAOFguxvftSxS2mKxAKxiiAndFzOu21eGX5n6EdYXpYEF3yA7ISdbbYZ00FPpeiSwiqCwLuN40DYrEBfHlhCvKshHig2jeyGeU4liIrRDT0RSLNK4Sj6tQa4XIPDnf7riWEesFO2yJS+SJxQVBuJH1fzhFDSARyWhnMz54t2j74seyUOPrQrqVaS+LnfFAXzEG+B8lB549uPoC3F0u8Wxmjf+cMu9BEGTdAdcdWXHBhqK70SIJMDd5DyYRqw5ymOcS5Bvv+1hfWCURxilrLdcQd+UO5b/sGs8tkRFuLLsh5iTgJOAk4CSwZiXgCIs12zWuYk4CTgJOAidKoBPLYrFY2t6adJDNtHW5ATAAOARa1wZrlAGHrGY/mx1ABQAYQB2AMP5nU2M35nwHgKOs86r9LzADDcd5K4n5jRYbKLTuARcAPgAHAR1w0cJzC+1IwBOAy4pZ99qSGXzdLabv1h5TvmmLXEHp/OBp07f1ZhEKtANwAuBkrzKaktb3NG0DJAMQA4xDVtaFCOdj4cE5yOip9v384IDxN8i6YmDIxEe/YRrHAMSvNvltAr6jIdM/ImuLovojrZv+20siO9ab2bsfN0f/co9p7Kc82kKZgOe0kbYCek5LDlggEKAboGRNp068CuuSBpnxnf5gzEHM0E7ICcYk/UiyMRj4nU00x9Hwg1DDbQHXAP4vjXyfm0QY89wPsJzxjPwB/hkL9H/1bw+2LOkyU8gaYW88N1hN+0YJKrA12LcnLNUmZGfUJ/j4qPyjQWoxZ1aTrKCFgK/Ih1gAaI4/Y64w3/53KTO3IXjaicGmBnzjslz6hedH8eRGL14X+sGwrCs2i8dY5/l+VXhsKM4glNVFphsUa7Vmn3wPESZh6Eh99ogGYQM1/v6efGPThjL9sRy4yHi1ROaK/aQYIOaa3m+aJF8zh0plWUIQWjpbNxHI6ukUSQRELAsMc0Xz4PTG1uS2wWTu8jBLuoHrk9whldLaAQXWvveG2v3ptx//1E3f3PoCO+7ad5qKBswf7PhR8+bDnzCfGX6NOZpnSZxPW+oHzcHCFnPl3BPH3rH/T28YbE3Grzz+hbkoa7H+4KaINQRXMtT7J5QBfxb6oFNMt0spDgEe/bHyndxeuR73bqru/76Pssjke7JerXXxXePxoz3NLBlupI1NkUxHmmkjzmetad/3jwoxr0vgkRbueuYHceZlR4LAjAVByPpkyepTiXI1f2MtPaBsnxto5TIWiDexUmJdx/UOhCbyJLE2QOSw7i9tGnNiqaz5H1PGsoLrAJUpwwJufNpnFUQkZMUtGnJNPTtF9Pgjsp4YFuETafDk4xj3aEwHo1juaV7n9GjIVVVIS9c09MDpV6SQLXoqbpG5i/iMjPYyBu3zFnms2rNR7qIs2bKkLE9hnbGS7M/ld2TKGom8WY+Q+TuVUR5YLkH0cw7zgfnCtXfr+YbVGDLjPQS58d2uuekKhNnptMGWRR8xznjv4b2BzBhlrWa8YDGy2HptcfkQspDGPJOZxzw3bOylk+qyCnU/nfa5cy5hCSxj5WDJWZ5T++W6CVeGzC/ICzv2eX9lzbZ7BN7rx11cikt4MLmmOwk4CTgJPIck4AiL51Bnuao6CTgJOAksJYGOmyaIi25NKbs5AYhns8KmG3CJTTegPQASm3dLBLDJB7CHFADcBUBi42MD4AKQnRJQOZPeEXgBmEGgXQANMnUDDEPbnnoBJAEWUA+ADbTuSbY9aOuXFWtinxn9uVtNaZd8jhcUtbYst0xt105YTHA99adt1J978IkMaAugBuWhyQ8YSeLeqF2jVQ34DqjN9QAcnM99J2WxUTDBVsXK2JqY1sxe7QWfL3fnLdM42DBeb2B6rysrUHdoksqYGXnrqOl/8WXm0IdTM/lPT4vL4N7UjTZyv1FltIbRcR6TbLB8ASD5mICQ7kDAnSquiQ+rwWqtKfhEXmyOGXvI07oog6ghIUfrigAtQHzhY+3AWKB/yYCSq5kYz4D+9COBeRlPuCtpb/CVLUGQfdeWKFOFAOdq4/mh9fL/dWSuWd5db/Uc2eofuLNg6ttEVkwXas3HaiVZ72gcrZIbqMXttcEw8Q1PsE1k2p2YIwtJHTGjuBVfGfLi8UGTlLI4vryWphvy+bAokDaSFcWAH3hJFIRzlWojr/NbcZJFcgsFqTHTitPd6jwCEsf1KCBeTfiBj903pQDdrSUsLehb5ima9jaWxrL9dWv/F8zLB/6XEGUFzvAaRhYVMq1Y2cPXZY3DY6PNoyMDSWXdcDy5LspW9Chz2Auy8aGhya/vG9v2+MDk1DHFqHj7/uI2CEmTTxtCoPNmNiybP9222HBFC4zHUifTq9kHhrHWeOn4l18ot1AvnMez2xrmrCfdaTFZwW+AuZYF+U19JxYJ8xxyg/W3uvtHv9gGyJXnfC+aLYYb7wuS/T0tz391Nc3qpSyoBHK+l8joRZYWXFslZoWA8zT0smqaekfETzOWq6tpXbFsB578Ax3BHMb1D3OVZwtavlgssX7NC3L5ZMkKzmBthqy1rrRYl7tdOdlSuAduTyB+WNuRpfWxvtSdmC/0QzvWkdIGje29Iir2qW+3y2inZHw/DbQ6x2nmx0kqUXupCKJE1kixxn8rykWJDI4yWbz0iqScSNK4rHmzUw9YiBDqiwx8uYU6q1gWK8horf1Mn0Oi8ok7ONZ+rBTfpLycVRG/k5g3kHaQFcxF5AeRyDsGlmqsdTxv6x3Cnvlh54id9Nyv23qGNcges5ZWjDv6mzH1jHVkx/WijuFCz1r9nEq+EIt/pgwpZuct46/pSIlTic399mxLQGQF8wtiHWKYucD7FnOJ58XfKaPowDOFtXFG50NarBrh+my3393fScBJwEnASeDilIAjLC7OfnWtchJwErg0JWBdpNhPNvVs+gG/ARdZ8621BRtzwHI2+AAGZDY3VjvRao8CFFBe2+3GaohVwASgMfEc3qAMEAJQhTYs4Ada+WSOW3ch3BawmQ0ZbQL86DXD3/WY2fmLbzCFHQMiB54QiQBQAeAFgIbWLmAIwBbaZmzUrCk95QBWo0n+/E6bLPCCPGgnoBefAO9WNsgLywDIHjaEuLx4UAG9cfdUMWkcGa+n17T27DPhJtUz7jPDb15vhDOaws68KV0+Z1o/c5XZ95sHzeQXmiIzbBBowC/Ksn7eIY6oIwFMPyOghL5aE0lgHsAQ/WIBI8YUx5AL7bH9ZwEk6m19KPNJ36MFCEkEWUEm0ReAWZY4Wq322vgE3JexD9iISzHAqDboqGzJI/qbfn1RNSsN3Wdu7lkfHXvihuyexvbSk8P9M5P5fKMx1yhEj4uwqJ8nsoJ2I1+Ik/+ljBXDsm5Y5lm3LBnyk3oxjXdcFiWVgh9sFABbKOTDuqwoymnm5YW8thTAOchasfzxm0Yu9MpJ4vfXW+mY/Pdzv2YQKlpEmlXEZhDwue3LWoBs0k1aKI5FqjgW+LX/n8q41GJsLucWyFxZesAUg6pJslDI8dLLRzmtmVm/zSu0k6wpTCltjMgFlBnQd8iKduSGpROxFFgrAF5KQTH9/PbK00+MVvZ+4y2HP/bAh7e963+rBYVhkRWWeF2ylCP5EXPbxFfM+uaYkWWN6W9Nd5Tv26cvJiuWqwvjCmCI9YHvWBRBYrDWxPk/VL/+IVPAJNKmZy15Wh66JnzPDBeC8qbZRI690ol8Pginq2lpKucXDylYxZxiLzBmU30/rmjwVbkwsuDxcvU438cZL8xX2rdH+fPKkKx/qMz6+/8qsyaeTrLxLTh3KbKC48xVEmsKZBn3tu55uu9hSWjrMgzXZaz/Wle8nIgKX7aIrVSxQSKxRfK+xROhoc+CFgGN/VRkkd+S2ZGfxDo3NZo3WY84tv0d60Z0ApA96wX3X1ULFxFQq/J8PR2hL3XOCoB8pmcRz1MsDxjTrKt8QgKs5Lrvh3TOK5VxRQMxjysmnvf/XRlLNZ59EF70LX3N2oMsWFvoS57bPI/JjJG9yvQ1z3v6mHOtNSTznPpQLv2EFSNE2kp11CmG2ADElGKcYeEGIce9V7WfuZFLTgKrKYEOWcF7KsHjeQ+z78689/+58v9QZn7ZtbEusmJFLYDVrKMry0nAScBJwEnASeBsJOAIi7ORmrvGScBJwElg7UrAgh6WYLAaiJACaAqyYQEIwL0DADlALpt8ADTO4X8L4LJxty4czrnFAjxA63DFQ6wKSATuBRHxCmU2VoAYAEGAEopB0TNtirt6TX5javoVT7iwpWHiWawqyqZ0Tdnkt18lkoLrAJ4BLAA0AKCxhuCT+0FE7FUG4ABsok38hpYn30FK+bRy4rNbS5j/kZkFyGxcBs4ho9HGs3RGAbmPK4+Y6LoN0t0tqETPpHM14w0qxoVgycLOkkkfq5ud791mBl9WMfs/UDf1gxb8ou18B8DH9QhtwE3SdZIbsS32C1Cinc9KElBnLSksqYVckK2NpcBYAkCyMVPQ4qMtHOc8+pQ+oL85jhagTbTri8powS4HWp5LuyGwLNBmLW2sBRGAVzu975G25Qv1FXLop7MaTj25GYVkr076STLrpem0UPeHD29eP3MeyQpbHRvjBPAXmfzbpQRAhQte9snrovje0TBZ3xOY4cAPqkmSBsobFLW5R0isJyBW41HeyowXyTm/tMblHyoIkpwis2SBFxXy0RZpkzdrzfioSI5ExAUa0HYNaQMbIipsFTjOP/QlY5OxQd/frrzwXnnbwGdNyZ8DJ9ZEIVTG0nisJSteWH3CrEs0jcSobIinjonIqMgN1M5TkBUA5sxLNKLtPJ0JrjaVb1Rurnxt8BYRPtmIAm0vGyPDNqiY1MwvP/qLbUsMshwznel4Q4sVd0V3KLdduylDNCRtomLplNaTMck2DpvpWFhPt43PZKWCAnA/uS4KJsWc7S77CqdgZF/hmYrEckz9yPyyBM2Z1nE1z7frJW2jnZ9TZg1mTXy7MoT0L5/jDQHEITf/SBlLOOYq49IGPV6qeEumAN4xRp/AHZTIh3WZjChUvYrvZy3JsqxewQ2UAm6bgjg6ZMz/syL45qe/J5dRnjegi7bq+HHFvcBco6m1EEC9HdfpTINun6M8nu3L6XNkDxlHPzDOsUQgtgvE4anSqH782UUnvE3/f0GZeYNbyJuUIesh+CBEIA9QKGBuoaTA2gwBwZoDaco1kIn0OZY71IX3Cs4hYVl3OgkLqt9X/oiyfdZ3x6w4nTLcOU4CF1wCIip4BeAdlrljrSvsOxRjmDUUK9P9HWuK1XZhecHb7G7oJOAk4CTgJHBpScARFpdWf7vWOgk4CVw6EugG4C1YD9AF6ANBAdDHpp/fOJf/rba8dc3BMavNmnRcT52VBAW6A2DjBgggHuDBAoxokHO/islt3mLywwfNhjePmXh6vclt6DW+3I2XrhkyvlzwpNEjZujKEZMfASCzMTkABtGepJ7WBN66gmKzxmbOxsDgd7T4ITZoN3IAbGWD1w3ALSYskBvnQFZwXtv6oSMzuzm02p8AHpEJQsoVoDqw0bTqs9LfjUw8lYqA6ZdLqNj0vqBuLn9/qCDhR8yhP5HlxThAC5YwXIdMKIc6jiq/U/kbkuGXRFrQpguWOkQF96NeNlYFYCDfbVBbCAfqimY5mq2ASJASkAP0BZ/UG0ATggMw02pgA4Ah1xcoo9VKmQBRq5U+qoLuVwYEA2RjrNn+t1ZEbUD5/7q2iPUAm3w0ESdlFbCpbgrTxZ7p/U/VrqxeXbpvujjRmBRZcaE0bpl/zFdIix3KWJ/gZojxd4vybgn9b/uC7Hhfzk9HA7kkS5JEoHZd/m2EdyumdpLMVOutfBT6ZWmODyVZWhSJ0WrWYvVLJqMKPyd6QvErsnEd74vjlL4cEHi7UW50Wvo/lpXFUsBs2ypDmTXkdzsy+9/12SYH1kVH/2A4OrxLxhtRkCUKTp9ZFzEn9WtfUjU7m0fMtXWmMpMnEWnQHBZZUV2CrIAk2avMmAGIob6MO+QEsEnwes3R92eFj/3s0yIe/kiq8gfl8unn9Zt1TbZQh9smvtyU66jjz5t5aL2IivxI/YjplVVHLjslYcE9uTdAJ58QwcwJAkpDBNs1MxVZsZzWfHu9qaVHg0Z6pN7KqmOzcto1HQ/1J1El2pgf2DOX+jPl0JdlRbu60+oTrAXagP2zrY2/qBNpC4Q31haMTdaxTykzRljXmG8A0Kczr5l/lPFeZdYDEvJm/tq15FSWCNYikM/LJDNcd83JumdIMbR3aRwOpa2sHHup6uRpDVNwbbHJnacgpkaEOFcMC/kPM9mkbNyM4lfIo5p8RhkF6p4nZGgXa8d5s4iQBQ7tnu/5zn2epRgWnSqc8EG7GePEeEAeX1FmbEI4E9tidKmLljmG5QXZJtxE2kT5NtaEtbiE/MaV4FIJxYczSVh7kHhmQZowvng+IPzz2r9nUkl3rpPAKSTAOy1kXVu5pTNueR4Rc41P1tLvVobM2+sk6STgJOAk4CTgJPBck4AjLJ5rPebq6yTgJOAksIwElgvKrdNxZWE1q9iIW1NwQADcHrDpASDnf7RHSYClZK5byv3GafeDgHZiGfyUsvXvbgN9o5W934QDV5t1bxgw5RuapnF0VP+LrNg4LisE3Xk8MNGOIya/eZPUW68StkRZVtvfanbzLLOWIxAS8xYP88QIAB8gB+3CigEkknMBXABe0BalTOtuijJtsoARZQLCWVLCap5bYgOgwwJlVjPdAh6piQo1ERbym765IQCsYYLeginfrJgbwZDpkTVG8bIxc/D37zOz91EHZAJgDvCDNjV1pw/YkN4kWf6WAFnAoQuZut8VkAWkA2PCuvCylio2kDb1xS0B57Bx5jhgO64/sLBB9siMvviSMuA7Fi/klRLgElq4p0oQWtyTgN64GIGwoK8BtAG2uQ992K2pbsFHAFPknkvVpePxxsOfqLz9qXI43fqxod2NyaFy9oH78LrwTBKBsVKdT+t3uVvqtmLgGupkNdh/Rt/RoGQcAvAh38/nvOxTgWf6ZlKTa8StehgptLav4MFxWqo3mnHg+2UdybXStBBIZVw8Wpikgu81qzyxaiIpcrKs2NFsJjUN9kO+782kSXZAc60uKwvWhbbrG0iL950I0FI35hha0JB29OV/UX5MJAMq6uijP1wOpnBj1C/q5DW6gDmiGOb+t+eEE/clFbOrccjDqkIERdsCA/dPCjhtRFbwf7cbJ+YEmvaAo8wRiAuOWY36tsb7PFkxnyTP2Hxsaq++/rHyXSrvV0VeUOblkgCxKuqVoOfu1x37zENfHrptdz6t195w9B/Gcq3md+u87k6mjA8psx5AxGHRwThkLHM/mBbGNGspcsD90ynBbAgHgdLx/vqntTSnBXkl2tdMC9UJxUsPzCGvlkR7jzaHe8uBOd4Xtvuc9cTG37lQhJkVZftzJZdBtFvrE3JgrWVsWAKD9YGx9G5l5i5jCi1462qLeBhYy3Adllas08xVZIhMrWWFXXcX6tVdp/ehH/+MVRDry3wMC+ZKlo3IFdSGLBFRIYnrWdnSWBePp6gVXlqTezSNyzRWQPjUC/1MwbkV60UR0L30QBwnAW6iVM6QKmTdyjHmz5v/d8iJDmmBDE4gLk7olGf3H/suQV/hIo6FkPlFjB00vlmzziV1B8Z+xmfcuZQ4fy0k668qQwIjX8Bc5rN9zzlvRNS5V92V4CQwLwFZV/A+irXy7cptRYPOGP6MPv9Eg/jbtHC8Q59eknlv/Om3vP5P7ji2jueTfcftVtLJ7v7yR9y4d4PLScBJwEnASWDNScARFmuuS1yFnAScBJwEVl8C1joCdEylA3yxaQFwAGACDGgDfp1jgEsAPgC6dlNzxpXqBNb+Vl0I8MBGifIgC8gAP3Wz6R1yxLGjT8GrZYVQD03/LWOmdEVk/JLqE06avtsAJgnMCnCFhjR15nrAKAAG2kId2azhNgRNZ7shA+gD7EEb24JL1p2H1bIHSLdas1xnQTFreUK7bfn8jiaxJTcskARIw3fqRbLuJLgnx0oiWhSo2x/XnQDsZEGi9mfVObm5kquo7+mTu6gbzNPvv99M/gua74AnaCQD3KElZ/sMGf6Q5Irm6VfPd0DujnVFG2Rut2FejsjdBnSkPyBWLGgNSQChgWY0v0FEUHdIHDbUgHyMLfqJY7crrxQIFZcwxCOx6VRkBW5D9ipDVADoQzzQF8iTe9P3WHowZhiLduzg6kUa+W2XR4x7ymAcHVJM3kNjrZEW+QK4gepq5sJXxh7jCPCXOUAbmBP/yP8bgvTQS6La4RtyWW++5U3I/dOgDCca+VwQz1VbkBMFX25sGo1mVSB9wUs8RUrwADDk/qkVatBGsrKQ3/75+aE+H5Hrm6MiMuZEWNh3ROS0FEhuSR9kxvgHuP9rERW9s/FAVVYW9Zzf6FHZeR37ukiJ6lUNOAbzyY3x5IA02S/f3jr+HpETApWzgKABFKLv9BEgNWSi9SXPnAPYJm4G9SG3q2xzcWZKhM9JIrQBg+9VHX5YMugReXJzKalWepJKUkjr5c31Q0ffuf/DMi+ZMSONIzlZhHxSpeDiCDkjb8YypCZj9xPKzD/WFsY9CTnYbFYiK2wNCZr9wfvfrnUum5HRS9RIp7xKfCg32fJnqmlN1hWmpmE58aI+z1pVIZ7WGrOuOEHgHcKIPmlonbLa6jYY8l/rOGQTzxxiffAMoJ+/3ikESznm7FeVWS84j35uk7+nEfTYEnyMZcphXd+i8XyVfoBcHQ9EeKuwhki+aeV8Kg5PPSeOLiPYvPjkLOfJJ5Qf+EkYGlkf+TViumgujGmQjusUyGLW5BNiu5wghLP8p0NQdF9tAcRu0uIsS1/5MpGS3SfZZ5s9JvnDly6Z6J8x9TdzApmzvtO/zJXfUbZxolauxPk7g3WDNZNxxVzmGYGFBc826htrfD0rROD5a7Ir+WKVgMgK3rPeo0x8lqIWiDnRsPdqAB+YbEYfuePouuM7e6ufvaqvcrOMLzeIiP3hwVyrVAjSP68nPu9G1gUs1ok8X2ZfeNsPtMl25SWJCxEaF6s4XbucBJwEnAScBNawBBxhsYY7x1XNScBJwElgtSXQIS7ieSVTQYbzlhcW9LNxBix5saDReqbuoAReAHC/Svk1ynwHcAScAoQC6NtlNv3QLtN3/U0m2lw0+S2+3CJNmWSiZoLygyYn11BhH2A2rmQArdhIUT+eWwCH1JnvbLisax/r+glAiQ0d4ARgGZszgBQAX6wurJ9qG4AQ8BwwnvZaSwlEv1izld+tqyb7uwWUqYsFlqxVBOis/R3rAgD9eQuPMJL7nlLTpEW1qR6ZvpsHzVV/8CKz79fGzLGPXyOXWJzX9sHeaTdthhwAaMdCoFcy/rxAFtp2PhP3pe9o06gy/wM6Il/axv/0LzJESxqtafoB8JqNMVqs3ZYtyBDXIYBbp5MWYkx0nYwMsNxgbKAdy//cD5CSutDnxKwA8EaOjB8+rZURx6128OLNOfWj39AaZszYa0+nrud8DlYWS6R2XUWoWJCettPe7Adndscbhnpy+YbQ1SgIczmZU0TRVgXSlmJ4tq9abc4odEVdAOxQPgzXSVPci5MklHub2STJIllgSMncrzZaieJeJE0dq4qsiATMWiumBRBvmbpR3QVNTdUR2Xotuf+/ovgwx7F20cTyvJq87FzeOOQrNsVhhfcOx8O+YmyCP5OvtA0iLTj3Dcq4VLpPmfsz/i2xhAzoX2vBdBK4eIr6UYWm6oZboUgWHpVqUKpHaav+ZM8V8efXvyr58b2/lxtsTVqXcpzfTeIC6DB+IC8sydseN5acaAg60vczTnFWnQm8wjdVJ9175ubN+bvWH2tuzP3TxPU7Iz87/uI+rzoXZ8krh9qB0dvr0RLAdvu+a8hlULs+FgDWOsUaBalFfyJjEusaa7qNH8R3EHPmKDI+Y/CYeBIC3ekXxg7PhZLG8V4RDdvmH3bi6UzWkM+nARlMyKLCqwdZVpDtROpnigtv/EQ2OjVZVWStRibfarJUSrPtIrqwOKrq+5EOaUF7Vt26YoX+uxDaz/Z5t/iT/rKybX9faqCL0LDPujn1OX3Acx6rKyzCWJdxZ0esiwux9+S5AelM+gtlCAqeC9RrrzK/Y2nRtrJzZMVSPeqOXWgJiDTgHZeciiBgzVxI+s37zq1HAxEPg1quflI/fGdnTNdaqb/toene339ituewCIuSFBK2jDej4eON3OdetXH8bTIPK+q6190+PH7nP0rNQdcRdwZFEBRjIOch76yLR/vOw/3b6zDWF9zfWWFc6BHh7uck4CTgJOAksFiDxknEScBJwEnASeASkwDkhZpsM61f0Ow8U6KiffE8WPEdyrhPAahHoxEtdzZCV5ncyHrT96Kc6b0uMBu/u2haii+bZQpYXXjU9H9rv6wRIBWwfADcol4AXYD9bLQgPKyWP5spgGVrcWGtHzjGZovPy5Q5zwbkBnykPgDwnNPeHFJvJRujYbFmK3UARLNWF92f9jlKGdTPEg2A91gD2FgPnMd3yBTANAAvCJSSvJCMmLheM7N3HjRzDxZM7eFHzcEP6XgTkIcyaT8nj5M5AAAgAElEQVTWA7STMtHy5X8AoL87X2BLx8ICueHKC1lBQKAFjezoA8Ae5IumNH17tzJEBJYVnA/oS2wKYnIgF/qHtmB1g8UApMepLCaQD+PgVOmv9CPAGGMGAIo6Ih8baHu7vkNcAVBRX+pg+7JNyNkx3hVU2t6P/lrQnF8BEF+hmufv59/91ENhX2++VzEntpXyuQ1Rzn+NZvC6SrX15PRc/epiPtgSp2a9/DTlGq1Wf7Opoef5E2mSxnLR3zuvnZndp3gV+5pxMqPvjK2HpVVOpZlvyK+5WgGGtT54X+u5xtvVOBj2JrWSXEDZ2DLcEFKAfiIjf9YSC2JbYmRJYd57Vdvvv00naYhbQFj9zJxqW1OpT617PCPSoduqiu+WvFwgJzhnKQuKMyUsutyKWSIyd6y55cZGWuw52hop/svU62uz8aani4H3oAKpH3ziDQOWrDp/A+k8l6x+X9w/3ZYDp2NBsWINRVjYdRYCmkQg7WsV1+VlIhvaawmWPbKh6BGIlye+u9w/yWOaqaRZyliQqzQtujK/EJHXElFxKG7FT2mVeDhOUyxrDirmy4Tmwglg4ooVW+MndOTWbjoiUrbPQL+Qh9MkGE2Qaj1pW7ustBYwxztlQRrw/KA/eB7jbx8Cg3WftZs59u3KrLMc55mwUqIOkI+jy5z4QR3/b8o8o35MGaKTvuOTOvAMbltpdbuQW+mm7ncngfMlAcgAlc1csda+9n2S9xb7fpq/um9ux7eun3x3PkjfLlIiiFOvXk2Cw4/O9D7xwFT5UR1DQYC5y/tnnwrddvO6qdeM9tReHWdeOiNDvq+ODfRU48BaA9Mk3s2wTUTZBNduxGXiPY05gvKGdRPLXLXWlPa5uUBeOguM8zU6XLlOAk4CTgKXtgQuhJbLpS1h13onAScBJ4E1LoEOYIu1xQkg39mQFZ2mvk2faL8DZAMSARyw6SkYLyqZDW+qibSomP5bd5ikccTktmxXgO0JE60DyGeDBECJqjmbIwA9QHCIBcBoNlpsyiAdeIZxD85nMwUoAmoJuWHjE7DZowzACupiA0az4eI62gx4DvBuAbTFhAX/A3LYoKv6eoIlhrXMsJYe1APNNcolW7/tgOeA6dRxVBlwZr/A48hEpT7T//Kdprh52rRu3Wy8UmYOfPABxYS1hAFtRYY2RgeEB79Bavw5FVrN1BVs27YNOVu/9GyqyRAE9BF1oj58AgghB0gJEn0HeUD/Ea/CbnQBkEg/0WkDRAIbZfqf/kJ+o11tou1o3kOAscHGVRDa9pRpXXtQBuOD69lwcw3ypw3WtRZFWuB7gazg4BKExKprUXe1Z9W+3nLDtuSJveP1YiGczOdDRdSOD8hiYkAAbDmMvJlmK9vckulEEmcyp9DAVQhhaZrn9NGMFe1ZACymVnIflYb0uzTJ9XublGIOMa8Ye+3g2x3ZLdRdwOVpt6MLsM5uqTxCH3RbvdiYBVZDnnudIP+VXALdA4Q5nxYTsO0+l2VChjulDkmxQFTYixYREdRjpXMWbng21hWdi2kna92OyK9PHW5unZE7rWt6/LnilImPzsZRQaA6c+c5T1gs6r/uNfa0x9BKJ3asLBg3EG3WNeCMZrxi2cj9k/HGNekn5H9Ma6y3TcdFDBsRFvILJUGL2GiInGh6mZ/o4n2Kxr0784MD8qT4kFaRo5orrDnWUmul6jyXfmfOWJd9scjPvAjLXllqzYZBEMjFXKT/095SjjWhqbWgdSrSokMEENOEec3zmucFazO0Fa7diP+ClRi/8YzgN2LD0HdYab1M+XZlntfEIMKqjOcqZDhrv7Wi2anvX1TmGfN9yhDXuKKibJ5Hf6rM2s/zn7pb61EsgC6E1Ypu6ZKTwIoSgNRjPPI84HlrSXWsWRm3/L8576fvEfH6ahETPZU4mD5YK8zKqiI5VC1s1cW8D/J+qWXLu07v76/U5/XfnNlgcsFxs7nYMOVc1nPDYMV8fVyeI032qFxI8p7F+xLv7CQCd/+DMs8b7okSCu9QzBv+t5Zye/Wduc0z/Iyt4VaUhjvBScBJwEnAScBJoCMBR1i4oeAk4CTgJOAk0JbAORAUCxIUQPFa/YOpOeQDgIEFQQjCebdcPVVNfmSjCTcWTPHyPtM8fsgUd00ZP2CzxcaJYLd82s0Q5bCZY+PGhg5QGjCVZAkGq5UGwAiAb8F9NleA1mziIAustpoFXjkP0J3fKMO6e6EufOdaACrqYN2a8J1zaZetA59WK5X7Uy/awOYP902A84At1qIDgJJNKASADUQuV1hhr8ntSk0wvsVs/pGCya0vmNl7p83E52dNPMn5L+yUS92QLZvF65G5wJfPdOqzmh/WzRWbV0gnG+/EWqXQZixW7lW2lhIQVbj1uV0ZWdFWGzsCGWJpg896rCduU0ZeVmsPX+KAVbRzdFFD6IcPdX5HFvQpm2isOJD1XmXALas5CPDF/TjX1vcEi4pF5T9n/wWE/+iX98S1Wjyn4Nm5VpIeExBRVwzugSxutOIsjD2T83OSku8FNTm7Kch1/0ycxMcUjrOoOBdEtqlKgxw//vPRr+dBckBBxli39dVZy2kZwmEp4PpsARBbTwv22PXBtgN3Su15uobiQDCXGcuXh158oC4LC8X9qOmzN+fVjs6lUWXyOUGbnfWwWPULu0iLtnsVjelIZBzr16wcQ7XES+xTVO16LvR7EjHC8gXVLws/onPLc5o8RWkOiN5LvNSbiD3vsEiKGU2NKXF+1j3Z2Y7PVW/ruRbYsaygGGtRJHIizCtsx7CsKvr0TjDdaMa9ciOXK+ajWVlhjeMea6CvUNe1bbDyNIiLtku7TkwTG5ye+DAkZMmzi/6xVpCQC4Ckn+2s36z9EBu8A4h4aj8vuI7jo8qUxRxCSxxygmuZ+zxfcQXFuclKhGenPu7DSeCCSkDWFdYtXtt6SZl3RQg962qTd71y5Kc3NVP/tbOtMFUsiqyRBv4DU325iWZu0AsCXZsVPOPdoAA8l/mYiGlKB3roR/ke85i3TpNmypS9OdOfmzUb5IxxrFmIeJPN0liZZY9mZ8xD3sFtgiDE7aZ1w8qailLJhzr1453axmxzBOAFHTnuZk4CTgJOApeGBBxhcWn0s2ulk4CTgJPAeZWAwAiA459XZkODaTkm6ZAOWEXYQNc95srfHDGlqwPtkKZkZdEwpSsBmNmwsUkDrAZsYOMG+AwxYS0UACT4n/sAktsYCjYWgdVKo51AfIDlACCAH9TpK50yAcrRygR8oiyAdjZaNl6BBbcpF8AboMRqZlImwA7loxVKMF6S1dinDJs4ZkFf3GBQDzRFKYv6W1dZ6IVjLQL4Lpf+4SMm2Hi98XsnzPD3qgU3+2bwlevN0T/fYqa+bAMlcg9AGmRHXAtP8gf8/1WBMpS/mgmwF1nwyf2oK3KDlKDPRpUBkLDAsPEr2NDSV8iLT2QMkEQfUj9AJ0gia4XBJhl5YgGzQ5m+BWSCCLHxRZAfWrN3du7DedwXOUOoWLCaDbTV6LXuhKxbpxMsKnTexZRSBQeuxYk3lwuT+5txrZm04pdGfmNnYGpDSdAby6WLfLt4k82m0NgsmVWsioONRoLsW4IrBDp4kEkTAniRK2Mc2dsgnCu6gbkQwlwufoPuTV9bLXGAHurN/3ZdsBYKbasOldMmr9YAcWHrvbUnmD3eF0wdKQaV8HB+e+PByk3WpdoBubF6QJYhz3kriwsxRriHQPSkA8a3rawg4jQYigLb2yCgCAiB8OLlZF2BuyOZHdV1TiBgXjEuFLxe/viaiZmT6dGUDAsOaJFhTQFsj1dyh3Sh2riK97Fke06yWB+FgR8Gnud7/rj+DDaarUEROYOaTS1ZZcniJ4tlhTWRi8KxZiuuYXl1mjLpJiftms0xnn2sNbwvWKsYq2xgLZ2Yt7wf/BPzVtm6qYGQ4PnE7zx3aMtZx0FZRZm6opwETlcCPIMZv7wvoTjEuv8iWd5u0vc7pU1ws0we+/uieDrwTfl4szBXjtI9j9fX3zXjlW6MCv6NYb4g62Xc2AWzfhAyH8K42TC5nrKJCvP6PQfSfrM5PWBGwroZGeoxzXTk8rilUGqthkmT2CTNur4rrBqe8ebZCxLEyeuVsX69Q5n3Lt71XqLMeki9cU16UMQL73CWdDmp7c5l1OkOB3eek4CTgJOAk0C3BBxh4caDk4CTgJOAk8A5SUBgOVr0BAEEcAZ4YLcDsM2GBqAa0uKQGX3vVtOaI2aFZ/pu+5IJIgBwNmc3KgNUYJ7Ocwmw4l+V2Wnh4gENLsgAtLwAvNnYAVhwPaSA9bttXVq1/dN3GsUnBAFgORtDgMy9yoDfr1ZGC5M6Uw7WDtzfuoKhbtyb39H+h+hgUwbZAKFCmZAiACTW6sMCLhaIBEAHJAOEJ9AhoAouLSibMgDzqaMNng0BEZiwp2r8y3Km9tSQ8ULPbHjzkIlnZszc/cgSYAeZW9IGOXD8Z9QXvy3SgjqfU9JGWR5SMktSIG8sRZC/tXChnoB4HLOkDgQOxAJklQ3OjdwgU+gv2sqGl7pjfcL4QHbUF3/m1s0XG2DaA6j1KWXkvlcZ8oo+tM5/6HfGgwWp6CcS13W/3ySrYT3UKXtNfnzvbTvTP/rMo4ztqdBPFd566lDgN5+KvOawXA0drSWVOO+lmzOFF64kRQG2eXmVKCa+bybjOIsUroLYFePKyI45a0k6G/NjLWtPdruA4ntRWvEyNMlqCkRelisb4atZoh8CWSsUjjay+lCYxZtKYUPERfIskxaMU9adXt+kNw/nDv39fXMvPhh6Lc0TjznH76xRoUgLwKGFflirMVXW0ASx6ypjYlKCe0xA3HatBcPC40RQaE33vF6B9IdEUhyoN+JIREXBBIpdwTMoy57WyvK4rApY55kTuEG6aKwruvqpTdjL/VNJwSp6c7mgNVjuZd6XpmarVySJf10U+g2tDWWRGJfLXdRh/X+4VMjVZZUld1oZ5FCyEmmxhIXDCWuKnl2WnKBqyNlad/G/PZe+sN/p1+UI+rW8Xq2hKeKq8mxJQAA/71e8G6K80dBadKXnGykVBPoevC4Ic9tlLbFeJMJrZTBRbITlv/GiCX/alPr2JBseGU+jV+V7/St8+X0MgkjLlaaM55X1P5aUJt+r6eEH85ocetC30tDMBEPylzpr8grgU5BBr56RIijkDk+ERX120vhRy8SNmpH/yI7VRVsXBxerKJfw7ktdeefFZRvvabxzsDbikg1LqSfaa2fXc+rZkq+7r5OAk4CTgJPAxSEBR1hcHP3oWuEk4CTgJPCsSKBDVuA72m6+ABms1QTaWQDbDxm/tN30Pq9oeq7bb3qvBwwhGDMa3ZAcbNoAtNn48Gn950IcsN/iE4Cf8yxobrXnrak67beWDvy2EFhX3wE1AMQJ/kx9IDBe0bkfhAgguA2wDOAOoA5otVcZUsDGvwA4hFShnvZ86scGjk2adUdEPazWKtponEs9qRObP8gNwHrqhSysSwDuRdnz7jH84JhZ97qmaY2PmMoj28zMXXWTNg6Y6mPUgTZSH+5JRjYc+z71yV+sBmmhsuhL6ghBYuODcC/6AxlRd/yRIyvO+YHOb/gbZ2NLGyGGiA8CKIu7MCxcyJALWEvwnXMhK5AN/YFlxV5liJKXKyNPxgq/2QDuyMm67bJjgPpYwog6tcfDxU5WqI3t9MOvvToRaWHCqGe6mD51TJj9o7K9yZe8sV05M93nZ63GTKvXz+LhycFwf189G2olWb6Z9xuhOIu5NPXSpilWkyyi30nIkO/WysLeai1+Mt8YB6nIilTa8721ejPOspzXbCXBWK0VT/u58u6aGdnf8I6NFk3tmkazsimX1UVatNv3LBIXgLAQtM8PvHjdk7Vrj2/JPz1b9Ct1uYZizDOuWRssqbkW5b/m6gS5ICCd9YD+ZRwfE0lhCelDxKyQBcVmBaSPZElwED9oOlTMknRAX2VdYA4IA7SENesgwPyS7TyTWC5rRVAdCxRLSkMQQ6CPVKrNF8hFzGShEOm55m0XiXGVFtKGWL+WXGqtF2EhZDRL9ITbkJMpRjNOKps2lHlunxTz5UzaepoxTrqJCEdKnImA3bnPugQ6JAVzjnc83qGukmHElWHem9Lna7T+3OwHWV9YjLaZ1BdpYDaGUbFXce9NI06/f6zVk4uTnKl70Vs8kRSypjBhLi+iIafpiBco/dXC1X710fc2iaFlTcSHF+WLeiEralHL6wW0Ynq9hqkFRS2Oed2H6YxhhU7W91ajYRqVybbVBYRGx+LijTrFxgLjJnuVeQfFVRvrB++1vB+y1p7TWvCsd5SrgJOAk4CTgJPAmpGAIyzWTFe4ijgJOAk4CTwnJYC7I4ADtOjZqADesxGDYACIf1pkRcOMvLNpBl652eSHAX4AqzmHTQ4a99ZHNecDYAMwseEByKZsgGv+5zw2emQAehLHrSsmC2BYF0bswbgHWl/vVuaZh4UDJAJWEgCyAIHWxRTl2HsR4Jm2PNYpHxdM/Eb9AEapN+0FqMdygI0a97MauJawAOi3vs8toYIlAtpqBIumHMzrKZtNIBYZ1I9yuPbLCkZeNblNZbPtJ4bNkY/2mKx1xNR2Iz/qZ0kSrqUP/laZPiFw4mok+gIyhjYAntIH1mqE9mNBQbsgp2gT8qYuNvg2/9u4H/QZBAftps22v/id+0BKkNHcg7SyAdLpFxtDxL63WNKIOnAufW7dAFk5X3KAFqTFg3f8R1kXmAn552810nK15B+vT7aG1xe9iVwr3hRW0uzwevPAhnxQ7TsaXfZonJjxelo+Nhjt8xIT5qXp70deNVIwldZ4PNra17xpRe3p1RhoZ1mGta4IWnGaazZjaaj6Jbn22SiiYriZ1HNpkgatRrJFk73Uk/lDJT9UgHFzeKyVlfsCczydrc/1lwtJJ77Fshr0IjTOsoqnvIxxC+gDsXdtbzBz1S19/zx4vDXylEgk1ipLxjFHIE5dOjMJsAZYl0N8LwuU6xGWJ8sb1o22K7SyL+JCqxFuoyrC7A7qc4/+PyjrAQiLiggJS+Kd2d3X/tmW2O8RwNkvTe5Q1ibbm3F6XVptyeuTX1PG3C7S8VTxtyGVrxMLPCSioi9Lsm9GUbB/Zq7ROAPXUGtfKq6GTgJnIQEREktdZS1/Wct53+RBwjtgTuvQtXprfGOY864v9nuba3qr8RR+YsOOTPEn0rg6FZSqY/our3VRGOZq/pDJZD/JC1ZY1JTVJwSF78+HGxMx0b6/1jgUNfjNPh8X6jXlDehlqqiXZllWdPQ7uC4qsTTKHWSaKIpNST/LTZSIkGatIldRbf0Pgnm34/20b2bMq5T3KLNG8k7OOx0V4N2Z90UXfeksxpC7xEnAScBJwEngRAk4wsKNCCcBJwEnASeBs5KANPkxE0drHvc+uFTCWgLQGk2rQVO6JjH9t37NlC67zgy98agJh3jmsJHB0oHExg1iAxIA4I5dEeA/5ABWBADWAHXWYgGAnu9Wi57NmHUHRXn2PPs7xwCz2Ry293jKbBhJ1Je6AMbbQNmAUpyHtijlfkgZKwEIDSwEIAKsNQV1tXE1uAfXUSbHLYlgCQzrU98SKciHcnClhGY1crDtvULf2fwBDFG35ytPmfz2VJvF3Wb4u0ZN1Pc1c/QvnmeqT9Ee6gzIipYbJMF3KT+kvpmWxupX9f2sU8ctVNvXf+c+tJH+sjKkfZArkBLImLgWDytjYQEhRBtwD0V7OIfrCHIOOAsZRVn8T39zDPlwDaQIm2DIImTHtciCc6kPG2H6iPpYooIN+sXorkVNPL2kPp93mxZ/IEj8cjjjjzaONbdMFdLZqbIfDAr2GM+HY2HZO2R6vPHZojdT7Y32mzm/Pyh4szuHwgOaa1lW9Ka/kPcrmac4tXmvmhb8mfx7P3cCKWQJxRMIocUuX1Qfm9qAjX4/XwQS4yCnquPeR2590h4ZV+Sn5xpRISc4NTRDSSsZ7CuEjdCkwUSSjEwmwZQA2HpYSx+4ruwf1vnVgoJ/qBzm74UcR9xrvv4a99Kp7c379fx0PLQOqxcde6Dzm3V950CgZabDMtYPjDkbj8W6D6oJc5O7rYx1+Khwvd3yjMKzi6Q1OTui/w9rtFqXdReztjBzUzErfMUX97SWe2VZUEwqyM2IwMsceKfYipL+9sEESlaBfpuV/NJI/ubki6ZfxyrFQtSoKGxOR9ant2C5s5wELn4JsLbzDss7oX3f5Rjve6NB5P9CSU/mwc2Z4k0Ex+UNaijKp7V8bxY3qsWBuOGZabloMjJ28gslkRglTVY9CjQB+cSCQpZP7U+RE6xzbVxHVhKzXhAuy7A3VR3ZXyyWPu9QvuKotVRBz8/nfcXvkRVHZJJYj8W2GkjbTahNKNuwbvKOR8YC403Kn1TGepZ3wRnFrjhfz/2Lf/S4FjoJOAk4CTgJnODj2YnDScBJwEnAScBJ4LQkIDDy3+hE3CrtVIakYINCTIimCQceNcXLdpn8pprpuzGUG6iDCrQ9pI0Q4BxxHGzcAkA4MhsrQGs2W2yAOIfEcTTpAfdt8FzKsEC9dU8EEAUYbq0a2CChkW8tENgwAqyjvc/9RpUJwg3hYt0xAbYDjnOOJRpequ9oOd+ibOM1YLlwszJglo0/wUbRbuSoG/e2brFsWdynHQxR2QK+tO8tyjZ2gwUvrXsbzpuPERFEW0w0csyktf0iLS43Re0V9/zqQVPbw0YRywe0tIGIIVXok+9VH20QSMzm8VwSdaA9EArUBRmRAfuQpbVmgKQgERiV32gvGbIC4mFv5zjkD3KDcLCB1el7rCroe+TD+OA3ZEp/oFnOcRsE2hIVFly2dehU4eL86CIAbAOt9iSygfyx46sQpLNROXs8q/lBtZr03yVQcV9gGrfks4n+2XTg8Z7w2GzezFWLvqwP0jAQ/FFpZTnTFxzbWPImBwv+bNU3yXXigCDQIOSsxiREEmMCkhESaSGpfonG2wLYD4GhY9St7aNC3/nNEmAQGGecFls5dAXhFpjq5RvNuG+u1pIVkumr1lvDsrLIy2tNodFMSq3MH5iOjT/X1GdUqIhtnGkFcbrB91rriuF+FRAp5gUxLS4kYYFskCNzpK4+iL45+629Bxo7dwoqYp7xG2Qk6yDzyREWZzxq2muUJTpZQ/i+YIWHWnFnbbHuorAgQ+5td2gE8D7zWz6nrlCIba9GVlDfkXwU5pMgXS//9kOtlugJk0WSUI4YH+IvNELDiiyYhsNQXvI9E8sD2/0Kvh0rpgUus+YuAXk9pzrXVfbCSYDA0rKy6H4u8x6DJUJD86ulpYb3VKx9Xy0vTaZvJGc2XpGYvo2tTAYNgyIHgp7BWm+jWje5YqzAMmGbI6hOKeJ9PTFpvWoK5YG2JYV8H4pMUIwKa1/cFbdLMSt4Zp8yyR5j8e/WPZye2OIt/Eghr5pertTbJkRiuYfqCsY9f63noSiAm1WeUewDUEYivsUXlP9YmfdP3pVdchJwEnAScBJwEjgrCTgLi7MSm7vIScBJwEng0pWAgMfXq/WQFda0nS0TIHnZ9Dy/bta96mrTe11i8lfMmvLVg1LOPKCQsRAGgEAAq2ymdnU+OQbAfbsywLV1sQQ4bl02dbs9srssjlkgClCcZIFrACk2hoCs1NHGveCaUWXqC1wKEM45HIc0AHTnk+Noh3Ee/+9VZiPGfQCvqD/AF89QMsSIBWK5xlpsAO5ClthEPSypghyQGaA/hABAJG6eaD/WB9yH9rARhIR4zISlrca7YsbUd+814bpBs/XfD5m977/OtMaoA5YJyJjyuJbN4yvUV00Bw2ftHqpjZUHdaB/m/9QbEgGLCu4JQcExNq3Ige/WBQsWEcgf0PseZUghZE090RyHbOkmq6gz7bfkECQM/5MsmGi19RZIClwfXIKJRiNLO3b5ZBxZgqAZeo36Bv/R5Fi6q3GodV0lNM1G6NU37W58y8HIzOIKZ6wvOLJrfbhn58HW9d+opQPJhnDPK2VdURYuecT3khFvnn9grDMmca3GXIUgo5/5DvFEoj/mNN7oLxt0k4uZD9TJzlfmDnWPda4l7toF/P/svQeQZdd533lufLHz9OTQGGCISIKIBAiBBEVKWpKSKNGyaEmWaDlsWWW7ZJfWLrvWa2+5vGtV7bpk12qDvbYsqyxpJZUly7uikk1apGhRJEGAyESahAmY6en84k37/71+3/Ch0QMMBt3AAHMvcOa9vu/ec8/5Trrn///ClRAY9mxpdxeKW1Hp9rO9nW4yXol8F4f+XFsERs2FRaQYpFk/qceFV9kjjVQNtGjBRYKEvCMrhX96LMkWpT+eEp9bJMigb71FxAWyQJYDmQResnKg8uLUUjpzpJU1GU9G5DF2IDXK4xISeJ04EsSzGPTRYf9krDBXMqfTR+nHg1gmSqwJAz/s1wD4Tp0Vm8IVIvaWQ/0j06rd+ntG7qEqIi36Uq6uJ2mWKOBHX3iqPOu7qgIDH06ytK9oFhXNv/3A91cVrpf5Grm+2wmecgyWEthUAkOygnmFdyPWvH0C9W+QcdJesQx3eUV+t8aRTuducnfuZufkhDEmbkTuhXEe5lng6pO4g3KtlZddq9d2O6tajaN4zS2fI0D2ukemgeXTukXpqMXDepmK4jHNYtOv5iMuv9EwtIgbY4liZHhp0gtkreEncg2VdJg+1w2ZCdSteQBrjlBEDFawvKvawXsdFhctyeQPmFNLS4vLl395ZSmBUgKlBEoJfFsCJWFR9oZSAqUESgmUErhsCQhkvFcX/wUlQGfAifUYDdUDR93OH7jbzX6m6TrPKXbvEd+FU99w0S5M39nMAN5DUgDms7Fh1wNIRAL4BOQE2AbsJi4C2vZsxkwbljwA9QC1AfYBlCAAWMdwzQToRD4AMKaJDBhlVgp8EmcBMIU8yYvrAcfRXjZz/WP6zq4MUBbrCp7L5pPncMWgkfIAACAASURBVB7iAjIDc3gAGogRI0709RUbSMoJ2MvBJtbKQrk5qAPnycMsR3guZTKAl/sB0G5XetgFFUVMvLni4mlFS1wJ3dh7PbfwBbN+eGZ4HfXChRWEyB612QWBwV8dPvPNfFAOC1BO3QGfaTdkx/N4LnI1bXBzp0X5iF3BeeoHEEsb004QH3zS7ubyyXbFo5YT/M5RuhdYlzEgN7I0oowxYMQdchqcj7xuMRMcg7DofKPzg8v7o8dOCJustvIZNxacn5clRWMyOH39THjizqwIehWvtRp6/dh3Ke05ANGVGIe0vRFQjCOIPAvITl+gTSkPCRLLLDLMCsrKPKff6O+QX5YnfcgbscAYNPTlEBgEysbKIlX8CoE4CkVQ9BTHogjD6FCjFjJH7UxTZFH0Kr6g2DTdWZXpSN8Px2eDIl/se72VbjAxng7qu1STC3+5h3JyD9WHuHgLAnHTn2nLO5T2BV7WO1J/cuZUf662lo3l/byayNKCsjEmbA4ZyKc83pgERD4UIi1s/jewjzXMrOwGjtqVBte828kK5EFdJZMeFhSylPBiL1jLFNU3zRX5RaF6ha3W5RYmlsK1XEYJvpSzfDmhkW64l+VZ0UkLdyiMvEWRG6crUXBKVkoLBPMe5v3GGuhddvUwqPlorQaWZqRSPu+yxlZ1hgG1eU/knfEhpYHVqcbNTsWEuD+IKu8TMaETa8d9Pzu077aem9rfdmlPbHqjcI3prqwYwn5U8xK5hFr1vGzl1JO1Vn2qc2Bqf1extwu3eEbGg4VMK2R7odFpVmKQFH+kB6FUcJ0+3zdU4lhnFq7w0HBv6XXz64VLxxXW6nqvGtc8r9ZItT5CVlzMGoWRolifQ0Ve6jvr+fuVsJSmTF9R6ks+uUiLt9J68QprXt5WSqCUQCmBUgJXkwRKwuJqao2yLKUESgmUEriKJSBAETDyp5Qwc7fg0y+62vVzbub77nDj9yaud2LMxQqs3bx5STErAMwBpNG65jugm1kOsJkyF0OAl4Df1ysBcAL0s7k3Y3cDZbmHZ5MHxIdpcgI0QWSQH9eySYIIAQhkZzVqoWHBwAFLuR9i5AtKgLBsMCEnsIrg/oeUjFRgE3ZYyUgMrAPmhr9TdtMkJ0+zJKEOlJMyAerybNPs1ddBXdhQ8jvlYU22T0gL8gWsBCgG5AWQvk3pmIigM27207vd+N173bN/c8Yt/KfHdB4Z80y0sckHgoDN80+p7U4IAAZIfsPH0MqC+yx2BGW2mB0A1QCpJ4cZIx+zREEj3AKsW3vRF5CtxfXAmoV2RS62mX2F5r3OD2R0rVhSbOL6CdEa8MAn/QTCgH4KUUH/QGa0P7JnLJhrrTWREskfrPwMMvbPJjeldX8pVpDtFQXVTu+u/8bjTf9CRzEtZmK/dSFw6Xlhk4ANFjuGsQPZyDgwYo3xShviOofxY+Qf/YB2pQy4/rJ4LowJG5uQlbgEo7yME/oz+XEt19FHyTuTHEataTYlMIaBsgm4XbS7/URBkqv44k/T4qYkLw710rwukEiuboK1OAyqIjbG23mR9Quv4Ut3vN/L51ZdcCBrRpmMKwIBtxfkBmdZhMVbCawwl9J2twnxEWmRdmp+S+PCWxGNsyApMC8xfyBDi8Ogr+XxRiUwBIohLuhv9Fv69SioN2j3awVQHoLqmssLcRN+KAdQcozvKhpPk9IK70oy8lzjCSEt9L+81uRFZRDbwsmgKffkQUpXh/60yI6DCmT/rO5jLjLi5402z7vi+qFMrU8F9WqEy61ivCkeWEe1Ernf/uqJtFGLiwtLLHsu/8yDh9/K+eZdIee3qxKXCKxN2/I+x/vWzUqfUJs/IcuEB/X5iUjxJ8JKTcGr5eqpGhzaodm+0gzk6TOV66e815jKvbHZNCzyRNYMRSgOoFobT2fqU+nq2nnXCitF2JhO0yAqjq7Ox3uTXrQjz9yCxuE5kQSy3lC8MqwcLI5XUYhLLHDzpvcAEpxCcVx/s4bMvY7sjMw9GYThShA2esFkLi4yKPywffvy2Xol7UWut7aCZYgmAP3HDFHkMiDJyd8UcnjM7SrT9wwIlfW1/RVuJN+uNiyfW0qglEApgVIC7xwJlITFO6etypKWEiglUErg7ZbAf6MCAEgD8gBU7nDTH/Vd87ZpN/WdywoCXXFTH1lRdEABHQ2AanP/BBjHBh6wcnTdAQAFsMaywkBswFYL3gnwgfY+JAL3m7sO8uXgHMAo5AGg53uVAPm5BwKB7/Y8Ps0SgvKbOx0AXwBaNlOAtKY9bgAhACzAPwQCRABkCJYEXG+ECYAuxALlBbSlfKZNaQCzab9TNgMzzGUO165bqnzbqoRzlJ8yK0DsID801sgfec1rH/qY65+fcQd+uqnA5re7l/7lo8NycK0RRcgFGdN2v6h0RcfQ/YA85hTmUoX2pcwWjwTZmKYy9UM+PBdZW4BsQGrqZFYw3GtuWEyW1s4XLSkAe66o0O+wm14jRgX1R7bIG6sBczNGH6a/Insjhkye9NmL7ln++933APijTZ235fpJadA/f2/l73Tvrv/6wwfjR/ybq4RAGfRprF/ow/R1+pGNQ8YQ44F8ASUgq2hfDrPEMMCS8QKAY/2evOi79HnqQZ+G0GJskydEFuf4nb6DVY7FLmF8XRLokAsoXz70K+o4Vbm0mYjjvBEFvvxleN1IDEYYhB2AFXXeqliJUEjrWL+bVOLIC6dCydX3vnvJ809Unf9NsR1/InyRMvM8k+WwitvyQX+HfCJIvUKsFo/7Lj87n+xSLFX/ubwIIAKNQEV+Nj62pTDXSqZGXFwr9X2deoon8zsym4jVu4RReuIdvLbIMo172VbII41c2GucF1VZVQibFFXhewLhFbPG9xNfdk1yGLVXa8MB3cP7QQ/3W9cK6TMq2yFZMYjfpFgfMkhxseRUV2wcXzIMRepEftVlcmHHmtiJ4yDr9/NcBEZycM/ka843G+P3lH33rZfAJmSFKW+wFvMOeJfSAb2z/JgfxnI62Fh3naTA1bKyEDlRF1ERutrkvFs9P1MEYas1sbu9XB3LJmQfKCvBb9eJ8Ne18TyJKu4FERZpddmT66Usa0wvnb9w3F9oLTV4D+V9WeuV9ymNU9xyrucAMZEXspzKFxUwm3VW5lGRxnSAm6bXOwa6IX6Q3axoNrMa02ebM3mm4d6uNpPfr09EH7pwsjIZhDOuu7o8iG3BDYUMGDc5Ip39e7qA+B3/QfJjbJgC0sXLif1RHqUESgmUEiglUEpgMwmUhEXZL0oJlBIoJVBK4HUlIDD1p3XRh5UAIddjFOz+TMvt+rFJ7WMiFzQTN3HfTm2a/thV5/bKdRHkBHELcJ1kfvW5DwAUMBCyAvAaEI5NFqAcoKtZVvAcwHHO2yaH+wETjYgwKwkAP4uFgRUE9wGCAgqYyxWAWABWDgNODSy0Z5mGONdYzA2ex8aQ+wEPzc2UabdzHtAYUJX7ra7mdsrM8qkDm1rbkg403pVMs5I62e+Un3wghUaJAfLn4LoPazu75MbvO+f6JxfVBnOucyJ3F34PGWFtgTUMMoAsYiN7q9pwQqD1Px/mcUUfIzEtuN9cP41awFBuQGy07/nkNwuObfXl/EYSohhxY3BFZXuX3DRqvWIkG5+A+Ywp+jwgP7IHrKDvM6aQN+Qdn2at8iqiZ8QNzKgm+SCQ8wbChDbCxdgxJfoR5TKXZvRl+iV9n++0K2MD7VL+pmwWaJO253c+yYc4NZAajDlIQfoq5AgECGOLfCA0cL1GXlxHvU4S1JsyQLzo8+KhfuOhrSw/+1W5c6rKXU0kUgItVZXDG1cg7t2ymhiTimgvSdKxOAgaYah+KQRFnrj7q2k+drKdexXfyR1Wojv9dEJK0cPnb7fmM23E/EK99wg5PtMMVmr3jH9x5ivL3/nCYrrD5ixkC5F0TZB3o+1bft92CcjrU66Y9EEXewkB6zIF8FoyrRAX4SkCvTzLCQDV+EGXGsf1TNUKWyG3UEURJYl87ysHWVnEupcxbi4Zt73gV9MDRsiKKAx8zWlFXIminZIjYzcLI7/j0ry52k4asva64BVpS6B0r1YNV2uViHl97cz51ewTd+4rY4BcTQ176bKMrtVYBX9I6Ue05nxonaBQ9KS4IisExaUehlfzgoqw+0nXb0UrWRpfqE0m1eZMm5gVqS7paJVlfmcMcXQ0AOfVf35NoSJuqE3kUW3ZnWsvhQdqE735XrvyPXIhxXvBDhETjF3u1+D0WU/EQfqNLOmfF1NxRMG59c7gvW4g7sF9hMcI8q6vmUC6Ip0wzsL6hEJiufzlxoz/iGiTuNJY+cDi6XDqwvHqICC3DLRc0e84P1JdUQ4YuIwaHFhk3agcf94PI4iNz6lMK2U8i3dGBy9LWUqglEApgatBAiVhcTW0QlmGUgKlBEoJXMUSEFD4MRWPwM8A6ADzJ9zspw65XT960FWlOJ1eWHDBzLiLJhNX2deTFhdgpmnRo1lt7p8MsB4N1gsID9nAhp2NGprZuEDhO7+ZBrdtDgFD+G6JQMCQB+ZeypzrAjRyLxYG/Gaa3CM6bK9wOUM5AQetjOQDoGpECoGmKSPWHAakcg1urNAGJz6Hub2hvqMWHUZWDPxXD5OV3/42rW4+LaCxubOCoLD87Hr+brqg2nfV63PXO7voZn/4Ztd58QnXftZkBnBtQbxpu/vVlk8K8B2o0l/pMSQteIZp1ZOVWZTw3SxZDFw11btRd2AXH3+tuHqyCr+GyyfkZC6VTNvWAroDiNCHAfshBCAvzBqBtgDwZuxY279m826m/bwhZgRtR14kxgGEhrWjgfmU1cgoroOkMDdu3EJ7W5wTyEv6tREqEIKMHSycOIeVE3lxPWMAt1EcnGNcQXDyPAJ7IwPisgz6n4DTUBrf1U438wSgCiv04nYvnZI2+LRc3MT9LG0IQ6k1GtGK/OxX5dxCOqFBMt9Jo37m4n5QzC4UxZ1hxzsae/npIJAPrTRrCXUkjkW2zcG3kTN1JLj2zYJ99p/uH3r06ysP7jzVm/sh/X1GJAYyQUYWx2UomvKjlMCbk8AwrgdkcSLLiaU8z3uVOFwWSDquWBZ1Ba4QtYcbKMX79ZnXsXfTH/IfpWtjfc2SxBtXHIu2vldkFsR6yVr5rrUEEjGxmdDt/cTTBFSVDKcF/E4LrJ0VnrtHzE4u4rStuWVXluR7gjg8nhZFu9dO2q1OcmJmyi3IUiyX+6j+r33pxf575nYw75Tk5Jvr3tt5N+3N+ynrM+vVJ5TuU3rQl6M0H0Zc0erzLBZpURtYWgQC80UcFGk/8PqdvFmfJH6FlqckWvNcf0XzfEvzPdazrOukmh+6XXFYfL++z8sCozu5tzXXWh5Lls6MH/KDAtdTw8Pr5WlvRS6oIlEWXY3SgVtO/bkfBkIHayXnTIHmVbIZXOYVK34gM6BK+kWN4EYYpzMzBxZ79clO0Fqs18VPXqfLHpk+2D2y84be2vGvRxPzJ4LxzooMOjImCIWuU5g1rC6o/8WjKKZEaf6cF0SZiJzf0vnLek/ZzgYs8y4lUEqglEApgXeGBErC4p3RTmUpSwmUEigl8LZIQODgrXowroieUMJi4XY3dsfNbvKBvuuexnA8djUZNRRpV+TFN/U7Wt/HhoVF+xuCg00doKMB2fhsB0A3sM7IBm7DWgGNRHY75vrJrCf43SwXeA6uY9j4QCTwNy6huA+QHvAUYgSw/4+UHlACIN0IAtjGE0CYslrMCc5zvwUzntN3CABkwEaVZwO68mzqyfUANViUGLALiM86a+SEvl4sv/kJ5je+DwK9KgE6891cR1n8De61fM3SgnNNqdKtuMkHJSO1BRYvR/8h2unmSxgiBgKJtoG8uVttekZg75PcfKXHkGSwjfVrZiPQht/NguJKH/luvY82pY9YmtN3+hhtxrh5nxJ93PomwD0EmcVtgUygHeib2w1o29ixcWwB5Ufbhj5vfXrUxZm5P6Oe5jYN6wnGtrmPIvA04xBChrHH94E7CyWshOjTjAdcny2pHwfHVv9DerbyvZmA0tVK7PflQqmRymuGbCkylaKtO/saTfWQ8MFZUfPjAOi1nfazQiBiI3TFVEXBt6tBEdXD4ubcc51GrIgXvo81A3PKlgMr/+ybPzgqL2TFPMdzTqj8N7ezxoFO3lhVEPQJgVhcS1mwTKFflEcpgS2VAMHFCbwtoo9187iGzrNh4I2J/Eu8wlMfHCyaicYYxIXcQyk6t+dJ+1sgqcu70h6PCnm3l0/9psbbmGYjxuhlaXNvaUXe/sw8uaSrR4rpobRX8nvPwGJF1o1SWp8MvHBRMmxospqUC7umFkTF3MmOCeRdUMwdyNaoWgnnZybrK8urXe8tIEvffom9w0qA66JhcG3AfywbeT/GApD3y8/KusHFdenuDFxBaQmSTzDIizCupiLVtY6JdlCHaC/VfFlHiGh3i7JgyEQSxHE9mY/rfd4lWctZ93if5T2WsXROKwHPvLFS7+1pzrQOiOVwSU8rmBYtjceKgnrPEOF73W2nLKFkaai/Gb6s059X2tQdlO6gVI9WGr1KpZ60lN/LUa3/ZKXRv1UuocaiOInCarJb1h5Rbbx3bPeRldvkIEqWH1lcaXrz6R/Gt8e1hq/YFq7X6rgs7a+/8KpyA+uL4aF5Y2fukj8fRfUvP/Dxv3Hmy7/7v5WWRO+w/l8Wt5RAKYFSAm+HBErC4u2QevnMUgKlBEoJvHMkAIgIcAqodr0LJ1bdxAdnXe09Cq69S96tp2X7PiZgcAJgH2ARoBGgErDx2HCz9FF9ArYBypkLG9P0sgB95lbINDPJBzCT33k2503b2uJUYF3BwUbuXiW0yPB7z/PZpFEmC+ZLHUY1xO35oxpnaLAbiUJeJHNrxCegKQAxRAWbSrOKYOMF6Gr++g2cHbWosOds1DzlvMV+4Dt5sTZTR+ptBI19Ul+rB8AQ4C/Ab8s17qm46gGVsX/eHf2fIFSoMzIE7IasAQhGNrTpmyIsKMTlHtdKDIrXk8cmlhWMF9oQtw4QVBB5fLd2h5zgO30O90y0KX2MvmZBremjg7GzwULi9Yrzhn/fJP/N3CVd0oWS6m/uwQbg/LAvQvDR3yEhrlMyMg5yDauDF5Xo34w55GV9mnlh14GXf/pcpfL7Ugs9Es1XPh7LQ0Y7zYpet5/5AgClDK6Uo/YpKwXP9QQiBakYjbTXr9XyIMTnhTzxt1cVmLvws+oFF/R35e6cVMdbcotjgZnfsKwu8wbGMe3JnMjckw4tKsZUbFnMeMxhELs75aPnsRnBT5/c4fk//4GJ7XZTdZnFLy97F0lAXtSKNZEWXQ2aJc0m5xWCATdrfQGsgVZFOar3Zb4kJNSTg5qi6IvWawOH4kRN0bin8sI7qj9Zt67F/unJtRPkRF1ETlPExbhCfczVqnFb4SuitW5/Urh1VTRqvZ/ks7JLqcYVwukUqeJYrIrI6Cytdb3xeuWl8UblRZFGHcW5WBNp0S8tLa6eUTYkK1BqYR0i7tDHlbAG/F4sGXB7JHLCRVVZVMgd1AC0z/OV9RhgnsWeGsR76Lej+uKpyUNpLzzamGq/rL4zEcTpOa1KrG2sPfYeq3XLX8mSIOi14jP9drxX3/tFNiAjBu6jZL2wpuf09XxZ9ni8NwxODxPvGLwfjyq6DAwvBmSFV6zp85j+bIswqUzuXlmKasmznZWqL0uLqgiMsNeqyHIiOSWShZgs++Jaelrr6Xxzpjh83T39z/da2dzJb9ZvWHlZvq3S0CUdOZBKc5EXsjIZWJpcdBH1Ycnkz+jefy1ZtkrXUFdP3y5LUkqglEApgatVAiVhcbW2TFmuUgKlBEoJvM0SEMCIiTtaXjcpoW1cc5MfUgjJmxSec5e8qlQnXP/sGRfNLLmwDkjB5gnAHTD1XykBtH6H0vcoAcoBzPO7WRyYxvaoBQLfbcM16gYJaZjLJcgMNM8A4SEOAHW/qIRbGUgMgE/KAhj6lNL3Dc9ttK4wCRuZYBpfbOwou8Va4DuWH5Sf2BCmFc8nfwMskoftysw9Er+bCyo7Z8TD6HkrBxtU6oj8IHwgXIjJYa6UqLP5tLcym3uqpoviFedJzLv/4kF37jf7rvU0pATtZ/E7yBOZhbStAOiv2IPLz7dMAtbX6bOA8PQfQGlcPH1dif5M38AFEO0N2ACRQTJ3SRQWIuodBQyOEB70R1w7UQfqC5BDXRnDRmZwHqICoMVcQkHqoAUOmMN4PBxki83Z3u+14+jcQSl/z85nH64nvZlpRbvti7SQjL2OfPAvyAl/JD/xYZIkkVf000D2FXIPlaJFviYV8U5R1LO02C1fOPt2JS6aENak/DeSi9vRSYyEYb46R6BjBd32l9KZOYUIOCal1nmVQt5jnNxxuNqdY14qEPPiPFaCmdvRJNdunhoPbQWGXlWfez7Ls6r+hrgrosjP5By/JXczMBQzAtqFlsolFK7ZRJbrur6G0ZL6qMXP8Yjp8G4MvK06vaqDUNdON/WmJ2pRFARhEHrNvsf7h8Bnz5+QjHaJwEBxQJG4vVhK8XWRFF4UhLd50jwXOXE2jnzkN67vIle9U3IPxXzPeM/Lcf72j8khWcG7J+9QrNcQFXcqqUPIykE8XhBFMuBLB5YVkBU6WlnSe1a/+fpf7p481rDBAWmRdEO3dGaif+6FHf9yYs/KnxMREcl6IpW7p0REwhMiEmSV4/Xby7VDy2fHdq/NN1MRHXFroV7rril+hDoSh/Jv8vxv542FhWuLvOA9w949LebU4DJ5ZxIJkTqRJRdkXVFUx3pnpnH/NNG5W8+75+yzs+ejatprTLfnQj9b66xVZ8T316b2LOe695DKVxU/M7XzhqwnwuTk9MF0/vjDlft6rZpbW4idAoOLrLgY58rKWVEMi1vzXvYBncBNJMoX5VFKoJRAKYFSAqUELimBkrAoO0cpgVICpQRKCbxKAgIT2ej8kBJgKpus9cDUe//Ke1x1T9P1F1eFD4oqmOm4YKA4Zu6SvqHvmLMT6wGw8X8c3r+RnDArgVFLB9tQjbpLMtDQLDBGY0NYMGDuA+wnLzTUjRgB/PyuYdnMf6/VdZS8MHDSSATuI29z04P2M8+ASDGgmEqbNYYF2rag2abZxrOsLhvrz4aS+6xePJs6YAXBd7PugLwgX8rP8wFrIVRG8zP3V+OKerjm4v0Nd8u/vcE99gOrrnfaLEy4Bv/I1AMZ/ZDa+JsCkXlmeWyhBF4jRgVtxriCdIJUw6UElkcWgJ5+BjjPWMKygH7MbwBdfLeA5pflimsLq7RdWZlFFGQoB26PkJERFIw1i5NiskNu9F/i3CCPI0G+Ij9Q3xqX9URNFhVZEd07Xw13H13rhIe78qudCDQRoDq+1u430zTJAy+r1aIk9yOXtNJIlhjOV8ThjkwsVuTWRiqkBWOfMWhE4XbVnzpZzBy5bvNucHnQnQgWGzW/u1shBPZUhfnQR2RhMTlX8377jrHB/ENfGBCfAjPTbY6xsV11L/O9uiRAf5I1RXFW46FaKPiLFsW63NgIZ89ngsKT9Y/XzJK0OiA0dI0smXTOncUyQ3+fVmc+qfuZu2xtv7pquI2lmRir+hIUbEVD8SsmFT9Hmump1+kXhyQfzVNFtZcUmt/zRNew5jYl8IlQ2u29LBds7VpRFJ6pxEGln3hj1YpsXeTmZzj/meLENtagzNokIGJiM2HQp2kPiAopwHgfl6XB/WIKRCwMXDI5L4xlVVGTS6ixAXmhY02kxWm5h2rqV71/YTXncNFpSieD58i90r5TT+2+8cLJqaNxLZncd+uZJ6JqclQWDrNhlD0cN/qdM8/s+klZV+xsL9XHFANDfUsLQ3bpYabi6L3PMwUY3hfN5aixGomekYucCJo71roiLSan9y/t1rndxF5hFZ4+sPTe7mrlkNxXNeUOarLbrkBu8D56ThYfzcDPBi5Rg8BVssLJMqTwx3Yk1cm9yfVTHfXheuReeqISyM2hKM98ncBRBHLFxvkrYmt4F/03kvV/RE6ytCjdQ5VDsJRAKYFSAqUENpVASViUHaOUQCmBUgKlBDaTwKd1kkDSAPMAifvdnv92n9w/SWOw4rnmLZkrMuki7w0VSfC/6Hd2T/jbx5UL339HyQJnj4L2o9YURlaMWh2YOyXKNKoRZsG2rawAv5xjA0V8DZ5llhDkgfsmwE5zH2XPMgJk427PCADc7rDRAzwG5IesASQksWbyTDOtRwse+VjwYTa0o66bLlUX6vAK8/xhpSgvWuaAmICykERYWfAdzT600dDI31gXyrpePj9UebK2qx9puJv/78A9+kmuNZdT1OeloWwAwmnjXx4+u/zYHgmYNQ59BOAJKxf6FG2C1RF9BsAekB4XE3wHFKHfAnBgUUC/NuudS1kJbU/ptzHXocXFRcukEaKHvkz9kQX9FXlBUACQIDPIO1xKcY0IjLwT5UvZmHsmydKxKa9IJ8b9HQvnwpvil3sTjSSJp30XhJ1BwOAsVCBTX6DiSuaHtWSACXqDAPLSV+2uJOnKny56i7uqYkGEyOj8lsv7b95OzFHnFMuCcT6n50PCyM1O4KV5I19OZ1XfKGkq7oYAzYWKr3nI8+Lraq7ayly1EQz6wihxkYu48Eot7G3srO/+rI18X87z4jmBlm1B5mvS+F+SbnhT1kd7My+7RRcpgkWxImJCa1+hdbKY1zWDeDo6Z5rcAzd170brikt1g50zDa/dQSnexXI5t1dzh6/g22u4p8tlzNWsxVhz9To96aj7ritSKJAcBQTL0iwpVgUIj3d7/Yl+GitmyECOhCg4lqZ5XSYZjO+kHN9v2yBkDWd95jPRXIxdw/24f5Lrp8gPFGBb8Sr4NYwqslyonPGDqKbVZkWWFhZ3iYWGtWvgwmnD0RQB8Oc6y9XnlYrV+QbX3C0rixsV26Lq+flJjceg34liXTctq4rNsmIg+gAAIABJREFU8hhmKcKw0HvGOtnFO6O5KYUo4RisZ+qoqaLO8D57TFYdp5rT7VD57u2syA6xksjxU3ZwbMfauK5rzh+fXpXbKrkt81d6a/HXFPC7O75r9ZZqmO/S79giBkHk3l+fLFp7b8n68v50steS3VDiZlbO+XsWTsXaKhDPYqjHow99xXr7uNJXlc4M3UOVpMXb1sXLB5cSKCVQSuDqlUBJWFy9bVOWrJRAKYFSAm+LBAQcsskiiCAuhdCEep+rzXlu5/fv1c4sd8GYIglqPxRMrYiswLc+rpggKH5X6RNK36uEuTwbPLNauLhZ0peNFhSDPdTIeTYu3Gf32m+Wh+ULaAeYyQbOgl9zj13PcwA1AYDt3GiZRq07OI8mO6A+WqJowQHqs+GDXCAPKw8AMudsM2gWD6a9NlqXjS6gNquLkSjIDFk+rISbKQNuWashgog9QUBy83Fsazjlogzk01ebCHttnHRj7zvgdnxy3s3/jgU55j5IJcBeLGAeUFv/hoDjLQ8srLyvuWODZYURc2ZNQR9lrABaAB6YxQy/8xsgn8VCof/h2ox+Bhg4cP203TEq3u4G21C/YihPxi+kDWQd/Ra5QhJCWCKvmkgIYlNnijlf8YJ4rOKt7pOnfX/SrxXteO6gVzRqhV/NZFOhGLfJajXKO5q/Wr2krRgWoZdq6PQyL1z2gl1FEHjP94PZx7vBqXs0WrYZJBSK40M2Lrqi8rS8x9znkplOp3fQOxBkPeFiZ0RWnJwJ3crZzL9elZ5JU0+KtT5gMnMN4z4UmMk84QjSa31ls7ZUXd7uJi6ff5VKAHJBbo3MUlFBtItFgeoNxVSZUjxo1o1MIKM0xjXS5EZNiCdzE4TiGQ1IuYMajE/WLCzGrjngMVaUchxkKSgFuvWV6fH61Gq711LsCjGkfscPpOVR+H614slkJZvSZDSmW6qSbSKR7klkkrG8lqw264ncwnmQP4mgY6G+hQJ5j75CXaUd6N1dLN6zdrEWi4S4W+3zMWJUVJoTetWKFI6kN3AFBR4fxHEShPGYHwRNnWBMmBXwukvV9fc0yISNx4JcRGFVeY8IhPuZ16UONKnR9rHh9cpv4IrqdQ6ZMSiynC7i/cLir1kHsvcLyrJPRg+F3FD5IkECxaYQ0aCX+sLbhcspiBERJImIirpiZiT6Xe8jhSf3Vd+twNzdsdm10+vxvAfvo3xRz1blasVykLqnFMPii60LXqs2mfzj4mSxJycwOFMHlw5uE9Gx/i6KAgfv3J5Ii9LS4vWat/y9lEApgVIC16AESsLiGmz0ssqlBEoJlBJ4HQn8U/2OJj/xE9iQzLsdP3DABY2+NmGhaz97xo3f9y3t1vgdAJGNFtYGn1LCKgMQbhS8t8eNEhDmNolPW4tGLS5GA1FvJD7Ibx2cXycXiNNgQYixSrC8AVrYENnf5irKSATOW0wNygYwekwJZO+0EpYN5raJZ1r5+J3vRohQdzaJgMtsbE3TlDICRBuhYfdvlIPVB8IELXJIi1FXUIC2tyqxyRv4/x+WEXDIXF2RJ+VY3yAHkdTadqZu+jsDERaUgbpxLfKi3agD32nrv0EBymNLJUCb0xcYD3wSg4L+Z0Azrr8sfgNth2UPAAefAArm4mxLC/VOymyEwLBxOgBCRWTQlxmXjG9A0jHFpYiifMGPktPzLj64VPNW9+ZRrz5ZaS5Xeu6sF2a1rkKSpmkaBMlCrZ1M1Wp+dF4KsWlXnjG6uddZ8cJn5sLiyUf6Xvjrp7PqPeMyytjeg3rJb32QuCze4eW1qSCrVQ4Gy408aPt9fzyQivYhmV2Ed9aCyk1VvyWbj0ezwK0o4DH9C6KCOYE+ZcGOjfzctpJXf5Np6hWHWavZ/DZopo0XdT/NVFweV6sENpAWFYHlfYGQWDixzkBQsL7QrlWXy22agu4KWD+l5SbR57nhdfTDa+6o1yJXjaNYcT/qK2v9ZqeX3NBPsqbiVDSTPI073aIpq4tYRGNfOh+yUi2SJFd84iQJZb1SCyK/XfXypsxXTslD3Uo7Tcf6/ayOpUuvnxZyObXt4/qaa7RNKryJOyjWZubY25XOy9XTZ8Nq/aHa+MwguLYnf0hRte7SnjyjRpVMr12JLC/WY7B5A8s51hDWeeZoFBawooS42DgZ0r7EsIKUMHek4xptvIfzvsd7+OUcvOsxVs2t4cDV2/D5WErzbv68yJEk6cY7REqsTexafUGun3hHuU+kS5PYGq3Fuourycl+N6rqmpmsHzwgskbWJMW8F+TPx3X13vV3cNZg6kadltRfT8vgpKg0i+7cPel+WVo8mffdqVNPh3dnySuWBORK/A/iqP280h8qfVHyZz1/FeEpl1GXU/fymlICpQRKCZQSeBdKoCQs3oWNWlaplEApgVICVyoBgYGHdC8ABZucR5XuclNS8hq7c0YazAsuXam5cGpe5AWbsceHmwvA788ONzB36XOjayTbbBuwZXEbjKywDZUB+RvXptGdDvcC1AkoGYDuoGe3KbHhsoCfgMFs2DCJ5zuf5MFmzlxLGYmBqHguYDH5zSlBPFAGiy3Ad8rORorfAP4pA5s0vlNfQFQ2oXzyPIs58Fp14dlWDtPIx5KDzSmxQ6gb9UTbHhdXbDaNoKBelM9kRptZOSnbtBwpv+Rmvm/STf32Cbf4RYKPf1iJTTOgElYctyi1aHOBw8cpTHlsiQRoE9oK66SblegfJAAD+gZWFoAKnKPdcP2ENZMFob7myYrXagX1VcZMon7LWORY9YtuJfOieiN7diJLm71V/z2n1rJKR3YTS1U8PWU7jiSpV0v6+VizWGpMBe12WGsstMRf5K7y/NNub7CUVE6dKdzZ57vezm7h9v61ZwrG2MC6ZasPuYPy0uWbA796/oznZ3uUPuTnzanQzU5FyV7FMI13Nv083OFnsexC9o3JnYxfhLvkB1/+8aUaWykUQjxo+b4CIa/P1cxtoxZjW11kt4GosPmKPkxfp8+aCz9ALPq3afhuiwy3vIJlhkiAPkS7sR6KiKBfFVg0QaTX8dSvC2ZFUOzV92X9rvWuoA+y7gGsDizCriV3UAitUYudL/9OnW6y0uvnFzC40NiUVyhBuLmryX9mnaAUuUgKWVusykS1m6RZrDFcyOOT3D4Frl6VZr4f1OLYnxLZMaHre7KySKLQp026uIUats8remppObV1A3cUGB8G2YYYZm49IgLiZ0RKfLg6NiXPm9EgEatCYZMUvLr6dT+MrxcpJeujdbdPGhtmTWtWkkd1Gita5kPeHWlXxhmxrHjfQ5HkmNJNSrxLonzDtWbl+3oVZf5lzeK9nXznlMwNKM/lHO8jWEH7ioXhzh+d2bN6vnmTLCmCid0rsrQInNxCOREUsiDpnequVQ4kHem+FINyLARJcLQ23n0kCDPqyPsy8z7vurzXcG4CdZlKo/hUXCtWssQ7fvv3J1/rtrxfOPdC8FP6HeWijcdfH5aZeYR3J9sfvF59y99LCZQSKCVQSuAakEBJWFwDjVxWsZRAKYFSAm9AAj+iawHCcVvTGsREqB7c7QrZvTtv0tUOaydznZQAA1wKsUEBrALMYIO1mdbYaPwK05wyd0/8NhrngWIaObHx08gOc3/EJg5An82dBeYFPAOMZ6NnVhkG4hnAxqbINMNYA9ngAdCgPUr5Bk7th3UyV0nkb+QAdUYD3jaTRqDwO9phRkDwyWZuNNi3/Tbq48HKRd0hKig/G1yTEZp9aOWxKUSLFUKJg83iwJR++AwLCE6Z2WSvyW3/jKvOJW73n9/plr9yk8v7XI/GP/mTD20M0ESb/+ww3/LjyiVgMU74BJDAhRHkxIFhe0KqIXPGCaAu/RcN5qeV6H8W0P3KS3AN3bnBAqNb/KfV3urYx5Z7/fhM6k9FnbRRr/it2ShcWeoGzcW1fiBQpbtjqrI8M+u+MRXkfn3ZTQfn8tsrq+n4yYV8/NyxLGqu5HLRUrj3fGO1wCqG8bEthxe2/SKLpzwvOeBndZlU7D/rOnN74v5Of2dRVLr93viOsGgrAnJL0cQXKp2kvpq42+UP3xOIuRYGAf2L+D3maoSx391mANPmK+Y1+jnzPy5MIFbpy8xXlOPY8JMYPDYvlsTFtvSkrct0xMqCtmK94GCuYm6aURwG1iHGhCyDLhJ6rKGAoUaeXVMuoYgfg5A6vbQr908r0jA/U69EJwvPa62uFruLQM6iNMjl2slPEoWw8Pw0kjsoCA7Fs0g6iaLphLKvqgQLcpmTiKjoNKqVvpT3cwHgVbEeyP+atFzZup59RTnZuyZz3D1KH8aqIlRgbREU8v1lvro0JILoJuflK3Gz95UwLj4st0ozaW9gWNuVxQLzH33EYligWMMciTtIyAoO3gl4N2A+RxmINre4VbxrXs5BeVF4QVGCuZnn8I5BQXg/pA4X3z0Vs8L1WzIx7IVyCpUnCvqd6fu4XFINntVerqHEgrUv762/KxdQVREVqdxFkS/zP3Vi7HNAakJaQIiggCHPha4XxMWxiV2F/8Bne+3f+6e1fygzxt+8RFSo79I9n1fi3ZQ8mXsuKiph+VJaWQwlXX6UEiglUErgGpNASVhcYw1eVreUQCmBUgKXkoA0ltHiB1Q1kmHOVRS7YsfHd7p4V9f5UU0Klk9oc2bWBACxHGxU2LCYRpmB7Ww4TGPKwCpz9cR9ZnnBNWxULA7DqEUF4MfoWmUm7oC89yqx8eN+QDuzMhi1WqBs5rqJZ7DxZzPIs0yDmsB/pilMcF/M8s1KxKwzrC7kYWQFG0rKxmbTtOPN9RJl4l6rl8Uo2Mx/8SipYy4IuI+NMuXl2bQLf7P5pa4cbEIHIOXwOfyNDCBVqGOuNkvd2AfOusmP7HULvw+oCCmCu6k5JWubXbS9AGAsAMrjMiWwIWaFuYCCvKM96Re0Gy6ecC1GP2aTz0YcF2ps+vnE9djAMujdHqPiMsV6xZetW178FnLO5I+/d+cte3uyQ+ik3edWZR32XMXvNvy4tX/CP3W4nhy7xc8SjdvpZ07kH3yuna8ceDk/sLeV+8saqLQJVlvjsiq4IFdGo/PRFZdv440yWGsUaf2WvDsbSSl3yWWRgpx2ZyI9bU9eVIuKzClc0ff93IvzYtZPpdMexavSzF5ba7un0sxdqMRBqmRuOZhbE2JZbFPsDSNH6dv0abSCIW+ZdwCqIGiZX+jPzEOcg2z9slJPsmQuuySY/WZdRm3iqgqRG8FibvoGa8N2telrdY5h+SiPuUvk8ovWhm+2/lvVMf9x/Yj7++3nkBPtRXmxluFgrTGQ0hQBaE8j2Qduyd7N1hUaW5cScxFhThG7OPD8hVa3fzTJRO543jkFIc7k3qkigif2nK+g2q7Zy3IZYXiKyS2YWwM5yYOwm2a79Gci4uOpiWalLx3+rowyVtVbWN+3a0xvVbd5V+UjgJx+zjstgP0Dasc/B8EkZgkXUIWCaY8qncjSwmvKI9Tz47PtBdwsVer96aWz4wRtaOoftaPreX5xTiTBtxTPYUWfzNkQFqMH7212DjIad1D2jn0p+Rqwb/HceMdgzuU9ERIRAmM0/tor8pHlRCGC4nNKKLDwXkgwbK7nQBmI+f2Cyv6luJbcsu/WM2en98vzk1/wDsq7rNWDTw7KD9HxLaX3q94HNGPUFJB75paPJl967svhP28v+j+t+ByDmB/D45g+55T+VyXeUX9FCfdYRti8oszlH6UESgmUEiglcG1JoCQsrq32LmtbSqCUQCmB15LAg/qRjQdasoNAm27PT+yU+6fc5d1EO4xTrv5eQAuAKDNrB5gywJ7Nkm3kANxHgRkDjHi+kRDmQoRzFufBACbbzpCH+cs1rU82Y4D3bNYoJxtL86NrcQLMhRMgGs/mHsgE/uZZuEMCYGFDhmYb4BtueUAk0KxGy82IAe7lMHdQRlQMAMJh3gb+Q1LwO88xYgTLCMq7TiJ8G0QbZnuRuLF4F5xn82qbQpMJ5d5olWLug0wbEMsLysR5gMSjrn5T3e358WURFsgbMJFyWMKP8DeVaPuSsLAWeWOfRjIhb5Jp5dMvORgjJPqRWVKYRvI1pY38xsR65VcPQdP+575xKptfmu3IB3yUe2vNifD84kz2mMJArPbCYuW6ird44o7gj77lB9P1b+aH49Q1DXAHAALEAUDZDu3mwPnJPimsT7isXtUM9eGhF7k8CpNq0c9DKbNO+1GgYL3yx6Hguy7Pplptr9IP/ZYretV6PT44E9bCovDbAjbRpGU+ZH4290xXLkDduYEAoI+zZ8BtCVZazJkAVubSBKIOEsMCyCNHADeuYT5CjpQNtyjmyutNle81bra5kEuY55jbOZAPsumobgM3LdtFXFwizgfzOGvlnBLWKGbBx1qX6B7mf9KmlijbTWjo+TaPRSIt+o0iC27M1vq3pqvJdJGsjBUpa+OoAgJtS3mpB3V4V5MVr9HfBnWXBQUxP1bGm9Ww3e2vRrmry31bX0G2FaDY7ZNlhbhIYFpPXv51KHC5gloUrhJlCnC+KnsKnXSRCIyGxvOivi+2Ov2lOKoN5Du05HgVebrNFlXbNUav2nyHZAVzHcD/X1K6Xa66XFwfE1nREDnhm7Xvt+ugANR54feCKCsO3HD+5dpEJ++uVs+cemr3WpH5z8jdUq020T2xdqFxdvGliYbcLh0RcZGLuGDe5j2PhMIQcyZzKO28/g6+/n0zvAZLBt7duM5cTXEt76VYatBvPjosJMo5jFUjI35Z33mfJPD1Q0p/osQ76sCdlawp1vRW+pg6aU9OExca063KoTteOrnz+vmmrDGYw3in5V2SPLAcwXqDw97zmWtRsmFduCDx9W74YBrvOJSfe+FPwz849URwb3fNm1Tgbw5bOz6g78jjt5VQCuI9aluUBYZlLT9KCZQSKCVQSuAdIIGSsHgHNFJZxFICpQRKCWy3BKQtLsDM3a1kcR46rnqgJrB7RrsXAWT9JcWxOC/vtGyMBpsaHYA+ZtIOWWGxH9gwGQFhAIe5KmKTY2vPK7TUhnkaoG9VHiU6ANTZBJlVAxssi9sAqGgBaLmXfCjPF5S+R8nAYs5BuKDBxubNtMQAkueG+UFWcJ2Z5fMMAGfICAOf2bSZxjwgNfWyAN5o1fN8NomWB9ebTCifWV6YpiqbYJMLdeFa+9tICp4xGreCfMwVFeC4bWwB5Sgr5TnigvjrbvL+51yoS9M12ob6Acia/2Hyv1t94Hlpqf8RmZbHZUuAdqOtaDM22wC1kGDmd5q+AFhLWx5TMkCydI9z2SK+8gs/cee+gcXFr33pxWxmcrp/0+q/70xkT8tUofOtoFi5Iyj6h7+7OP7B1P+uerX4QY3tJkAJmqZoigLmoCmKxcVWH9K+zqSpmkzlXu+6NBnbG3neBQGYJ7ou2ZNlUUVgTr2bFgpdIedPciUTKVCHFHwFZhaHYgX4lasYgrLWBHylvl+cFcgJ0Uo/ZGy/qWOTeBVmVYFV25wS8z7nAK5sXmOONcsy5MjcxHGHEvM2c+DvKWHFZpYFb6qcm9zM8yFtAdHMzR/zInM9ZWDtok8QF4ixuR1k1MZiMefyfOZdNLaZmwHlkB/lRE7HlMx91qDPbrVgXiu/IVlBm0FG8Xmy5QXXfTMcf+b5oPGSyAvviMiLDyXwUxcJdmSXihx8S8v6VsrlDTxrsEYTw6BWjUQguuMiIa4TtC0I2ylSjj+mcxWZVFyohH611S0GcV6kqO9V5RzKFd6CAm6fqMTxalyP2qHvtWPZajTrscVQKGX8Bhpjiy5l3mBOixSfYj6s1HZE1Zq8oeYiLUQ9yaUSidEQVROCVLu5u05ON6dbe2GjxnetHmnOtL7RWa49OrFn+aEgzD+gubrdXam+9OLXDp1fnW/c2lurTufZRf5jbjgHMKeau0/6lRGuG6vFnMK7BWQHsSF456BfMUhNWYb3bn5nruP90QiLH9P3f6N0UHWpa/24Q/XqhpX0JHFpFFz7QmO6/fU89U9P71+c2HPTubG41q/oWt4zIVVYI3nfMcuMX9V3YmNQGdYGLBS5juu59mtxtWjuuC47UJso2jMH8i88+8fhx5dO+1U9z/YT1I814meU/h+l/6CEHMp3JSRTHqUESgmUErhGJVASFtdow5fVLiVQSqCUwAYJfFp/s+HB/y3AyZxr3KToropdEU6vuXAycsEkawabCzZEEBeA/Wzq2AgBwrBJMmsANthGVgAcEaCbTRVgLhswcw1FnuYSaeO95jLKSAy0ezE353lmjYBWL88xiwojQeweiBg0tcx1BZssNm+AR48psakCMCI/LCwAYQC2AJ7JE2LB3E7xHVCQ8gNocg+fAITUn+9stNiwsVEjoelmboIGmpjDfAEiOKzuo9YmtIMRJKZhRr1M887kwv2UgedwP3khV+rDRg9ZUdY9Lj50yo3dc9otfgHZUR6u575jSoBoxCShD5SExbBh3sCH9TlkSrvRZhb0nbaiz1j/KzUG34Bgt+rSzzx4eAAotv74DkXnfvm8X7Sv81zCfOI3vF5r1jt3JvZku1DkO+RHDbAFchTgKBCY6221Jn6RjMu/SF8eYGTs4ScKWeEFedqIirAmXiJmEMdyMaNxXLh2ojgWCsAb5UW9100yVwlwFTPZT/OmgvgeHx9zy7U4LILAYy4YzMFoY2+hWyjmI+Z7NGD5NNd9zP+QA6wXHIBnzJEEfQWk+tRwLLBesK4wNvhkPkZbf6tdfjDWGIu4UaFtmY+Z03keFnUQJ3aOsoypbSFPulvdvkN52Afyot7foYT8qDcayRDGHGaRZ8GtkQ3y22r5bCjW+p9DsoI1D1eIKC3wSZs1MufdveKFjymlZ/zK178YzZyXuyizkHlLQfRNrFZo641a6JQJub1qnt1mCxWeN5CH4stE+bq1xAueV/EUQDvNI7+a5kWoMZxr7FbiKJ8RieGi2E+1agc6sdrrp7S53LyF55NMgbtzn/5xca3fwvG8aT8oTzo3tK7gHYq2ZO4YvG+KbDqSp33pfviu2uy5+mTHtRbrLkt915hqu+pY78TY7FpXBMXdIpT3i8pgzZ/U3/fr91M6J8UfdyPRLsKZ1p2H7jjp5o/NrJ19dmfUXZXvv8IzRRTeh3lHhlhgzXot8pl3DN7dzBWfvVPyzsec/A2lOSXekbEWYc6jToxv6nhEFiHnVR9f1h8v7pi78A2RKfUgzipTe5dT9dSZIE6fHNvRmhCZwbyAAg5r4q1KvEPyLg3BwLzPOsC7M2Xhd87jtpX+y7PO6Nv7ZWkx1pzJV2evdxfievGvv/Ir8X1Jz7tLv48eH9cfEEW4aoVYLo9SAqUESgmUEriGJVASFtdw45dVLyVQSqCUABKQZj1ADhs0wBQ2TmwyGq7xPt+FdblSrk4rhsV5qZZZjARzB2IbJD4BD4ykIFs2L5wDAMf9xZzS7yrhgggAjE2MATKmYmaaVEZ0GBEBQGJuPgB1uB9N3YeGzxl1RWVuo9hcGXDPRu1rSoAwEBhsqtA6A+yAsCB/NoacM6sLgH0AOerE7yQ2YBAZkAFooZp1h7mOsiDggBcAYcQoYLNI/QxYwbIDrbTROgJU8DfatgZQWOwNk82oJYYuG1w3ehhpxDnTMgako/yLarub3O6feEqEBRrS5pqKZ2Clwidtv0hfkJXFIxvyLv+8tAQMGDOLCsgt+gV9DPc3kHWcS9djLJTH2ymBevcR5hzGeiy2gH7/cOoFrbngqPep+D8u/mLy44+3srHbRVowHnC5YSTqlradFwmTziORFam0dztjrmjnRduPep3KbOLXQmlnZ3J431FwCz8X0imt7I4Ue5vtflrtp5lCW7iJRG6ihIrKjYj31aJRuEYtLqSwzdg3wO2KyryJKyhAfuZ85imAqGeUmMfNYgGZ8hsAmgFMgGJGYjMPMQaYN22us7n1ispIH7qEFQjAGc/DFztzG+0IiTw6XyIf6mPuv5iTt4wc2ER+yIH6MkdD5gAoAvhBilFeDv7GfQtEOvL990oAgdtKCkDGDeVkbr74m3akHx1Two89hA/ymeO83EXRhubO6mI7bDMhMBTTxXaknPRLAFv6JGWkXMzDrMOs9YzzLdXOfg33S7hs4h0BoFVu3QKRkLmIRT8Za1QqaZ4vpGnxvEgJ8ZBuUvGau7KqWK3HYep8LxtrxieSXq5A3fmCxnBb0Y27IjQou7nbuuJxYoIrPy9LAvR73ufoW39W6e/zd1FkLqr7bmx2RYSFDGLkoW9sdtUl3cjtuenl1bGZ1mMC/Z8VMXH/8ClmFRHJKuF7dY73YEiEhv7eOT671uutVU4rsPVeBbEu+u3YYjrw/vnQsN9CLvDuyjmbJzZWgnHLfDHqTpQ6MC5IowdzEGPiKaUDKmtjcs/Kr8pd1djYjrWdE7tXb5ZFRRDVkikRGciA99dzuo6xxnzJO+9Xhp/0SxLvN2a5wXoJoUFZKY9ZlkIgQ3bzTrSkFSodm83P9lteUhlzmVSiNhIWlJmxzHsqc9ErAnBvqFP5ZymBUgKlBEoJvMslUBIW7/IGLqtXSqCUQCmBy5DA9w83IWy4Bz6+lc7IuiJ24eyEC6c6zm9CSgDuA76wmTELCQPeeQzfzYUTG41jw00HmzdMxtFc5jDwyDTT7W+LV0E5LH+u5zvrlWkQ8/0jSgb8Wz7mdooyWoBXfkNj1XwCU3ZIBMAAtF7JC1CIzRxgx8DNxbDcRpgAiHCezSFywEKDe4ywGVZrAJygycZGj80imy42cR9TYrMKgAYwZTIyEgISBpDF/h61qiBv+9vIDDTwANs4T7k5zP2KXW8EEvfMDcq0689U3dM/iVUJFiAAPObvnmuRORtS+sK2EBabAHnmSmZgHbLNWs5DMW3LB32DtqDfAFgZ+IlMqVsJNm2L2K8s074XKhCq2585vxBZcXAxbO6QrUM24849fnvlT0+38rHjj6/dvUfXfFDExSPNYHnVqm9OAAAgAElEQVRVKA/AzFYekfMKxuxpL+i0FJb3ZdEP4ikUvtWLUk8+OZI8z6JIEbez/movy0I/9GpiKOTivqjKj3pLjvCJ/FqVZcWsLC2mBIqeiv3AXOOZFvybLTNzA/MiZTU3efhaB9Djb+aiLykxx65r0q7PrawVzGnM+eTBesD8CfjEvIv2L/PkFQHym2jb82yAMubah4b5QlpTHg7KD4iN1i6gHWsAZWfOXlB+WFm8aVdaw2fZxzrxv06eEBcKazsIFMgc1h3IANZayonbMfNlD+iHDJGZuRrckPWW/Uk5WJMsHgVzFeVgzYZ0R8OcctDeuEdj7YBYh2yhbFtKCFitLhEDxN4DuIwy0rfQ/Gb9RJkAxQjKzdpIW7Lmsv6aG74tE9pmGYnMyEVaIL+WSAc9O2h5Xp406vE+Bak4m2vC6VWyHXHFn/HyPO7LV5Q8bZ0QGJ4pBMJKEHrHxEGKsPDFVXgd/QNYPVhbSuuKbW260cyZq5i7HlT6W/QzKOCo0h9YUswcXFYooYnO0qnp2uS+pbza7K/KukJuvPqHZYXAeGfsMreMHljQvS9L/H8nt1CHRVh8px/mkwpevZrnfqKbpuaPT7m0/wpIhnczxhj9mH7woUtIgPHH2LR34EsJ6ph+4P2OuZf4FE+oHC9MH1h8ava6CwfkCqoul1a36Hwq65Dj+rSxBpnA+OIZjC3eD3lvY75iLmfesHdJxh3zA2sl4xMZskYw71I53o2Yo2th5I7UJosvzV6X9dcuhMf1hsS7/OjxN/QHff/3lf5Yaavn5kvJqTxfSqCUQCmBUgJXmQRKwuIqa5CyOKUESgmUEngrJSCNetOmxF3Tw8PNxoSr7D/hdvzA97pkXhqA1dOKZ4G2Exq1gFej7p4orpEL5vLI3FmgbfsFJTTEfkXpv1MCPLDrR7VeR/McJQLIk7XKyAhzi0Q5Rn+jfAYQUyby4BqezW8AV5AIprVlpuoG7FEmAA+u4TubRJ5lJAHn+M4mik0Z5TEXWJSd38jLfE7zO2DJQ8Nysqljw2iWE6MbTO5lkzxqdWF5jlpYGPANyEb5OMiPg+tGLVQ4Z/7aOb/DBWM8gzZBnmxAIS/QfqO9yI/N6Qn6hKwBAKO26zAtXjavyImNbH+o7XsR3H+LNHa3oo7I13zhb9ZeW/EM1/vLF7OxPvmKfCv/akse847P5J998wc3qwN9vvLPNf/82aUv1oMin+35UWUpaNza8Sq5SIuXbs6fPv5MtH9Pxe98KC3C5OX+fo3v4vjN9Udn73/4L7vJ8MLq37z9tzbVxOeZ+u2yZKdraT+N4aJZFOGTRR7eKBcyh5MibyhQbyHfeyt57Lp5Wlwvv/Y1WVl0O0na9SL5UY/kpEOMRZblHQX5jQWEjiswL/7xT1UqwaaucC6rUMOLNiEVmT8hKMxyw0AntHqZE/kkMV8AKjEHUj9IXQA3XM0xp0JWmGspiFvmHOZkc6H2Roq58VrKRp6QAlh+MCdCujK/UQZIASwbsGBgrPIb1k+Ai/SLQSwk1f2YPi9aDthD3sg8tInVB8AddQX0A1wHzERbmWdTTp4HccIngCDzCGsxMsPyA8COdYk6bCnxOZxvWSOoP2Ajz4dEoe0oM2UBmKRfPaCEljRlZY2jvSnflpdLeW486E/0HdaLycDLCHB8o4DVB2SccCb00pWsCOb0dzf0k+cDlxUiHd8nkPgWnTsq0pHAxICoWyq/TcrJKZubBwoTIh++JTdz8xqfkR95USX3Bprj/cIbl++3iuynTrV7RbvdS1w1DhdrUdiSLzhzrdOHBLnEc8rTWyyBoTsoxinjkzaYUbu52njhdsyt6yJUat5ifWpxTW69ulN7xTFVk6JS7/tRVZYzUcb7E/Mfcx59FSKQQzSzt0P98UeTXjgh0iLzw2xVjsOkFOQ8zehzY7OtyvLZsYp+4Z2SAwKY+eG7hnldqrb0N8auKa5c6ro5fhCpslpp9n61Pt59oTbZiWbnLiQKEL6oesp9WcEcjVUEFhjEb6L8h5UY4xC9kIKsBzyT5/E777XXKTGPUGfKzBrB/IAMjYzlXuYS5r+6cjgmuT5y5IH0wLkXgv+hteD90iYF542HPQnzTUlYXKply/OlBEoJlBJ4l0ugJCze5Q1cVq+UQCmBUgKvI4GH9DsbLTbGbDbYePTdxD2HXXJ6xY3fX3W1w4ApbFTYzHGYZrxp8ZslAp9moQCIxfWA9IAzgDAAX6apa+uPxXAA/OIw6wMDfu3TNnK2MTOCYLQ85naJPNk8sdFip2mgDM8kf3NhxSeAGZtMtMWoI2W1AK0AHEaKmPUH9yAn20CZVQTlIH/KgLYY5YPgAWwCtDJzfJ7F/XafgTHcz7nRWBb8huzNfYrJF401ymiy2iizUWCGPCgXz3zQfbR41P1n7/P6jnYq5SN/5MOB3OgLDyl9bnhuuz6QH+W2fjBKXr0VwNKbrpdIndHDynzFZR8hJMgXeRhIbEQWfZnz9DGeY+DwgEzT/WYZxN9cQ9ua9UcuQiPTNaNydjp3xeW9UgFuoj1t9eVzdDzZ34NHvR5wvAlRYTJkzDJeALPXPt98f/NQ8vLEYjB2ZGe6dA6rhTW/dsPqWPjZXfmpB0/0Dr+v7rce9l32XDev3SZA9Pm6v4Yrtaf1DNx0IPdcBMWVyo72nFT8iloedGf7WWNJYNFqP8izJK8E8h8jS4pEoSqCjjS1C09WFmHq9/Isn1dA36me55qtbtKpxv6CjCxStWhVGtnAYs1ON1nWNVvlCsfmZMAzrCEA8uhXzOucY47HaoD5CJnYfGldA+AKwoDfmGcBtgCsAK4gXQHK6Z+XbQ1yib5DXgBsHADqNucxxxm4jkwgLVh/IGtZl5j/mG8B/KgX5QVQfgVIzDNfr+9ZhTd8MrchK9Yh1iPkxTMA3wHwIAaOKzE3Q4JjfcFagQUGsp8blvW/6hPAcKtJZOoMSAmRffPw+QCMBLvFuoJ2MVdWfEJm/OGw3NTJAMutIJ2U3avcfA3O6TA5HvRdfrNCtUxNhsutXl7t1fz29FQ0/+SFZOfOlXTyu+Vm6WO55z8TeskRERU71BHOV7wufTVzv7m0qnbcVgJgaGVBmW3e9cLA5/nVPC+k/KEXkpQiFCuhLKZikZDVOGr1EoW5CIO2yAp7HynJCmv9t+6TeZkxQbw1jiYziWItuJlDCjQiR30Te/KkPtn1xna2Tuin8TDOdslSoab5m3FD2/HuRwMD+rdkNXG+s1wdUz7NpBvu1LWBYkYU1WauUOt5a+f189XJvcve8stjinRyoFg914xxNzUcW4zNS7mCMqkwr21mpQZBxxx38ZDRnlNMjXxq3/IHZd3R0XP7np/3tMT4Kh/PofzMpT+khHUc78LMl5C7X1TCsuo7NMsfFM8iwyDv0X43+v24lvxFnZfVXx6L+OC5zLnIkLUB91l/KMLm65LRe1R/5j/qNRutB+Geu+9Heie/8C+qL8sCadeGtxHKYtZoo1Upv5cSKCVQSqCUwDUkgZKwuIYau6xqKYFSAqUENpHAJ3UOIARrAGJZBG7qO55zM5+Yc827Ki5oArgDppi7JMAeAxXZmI1aHnANwD9gjPmg5fovK2FdAcixHlPh2/EaDEA1iwIjPwa7eiV+HyUvOG9ajGbRwUaLclAPQFojXjhHfmiBAQZRNtY9ysE1oyQJgBzlImAgIBP3mRUFmyz+5h5AHDan5jpDXy8G/bZysokEjOMaNnmAUGziIAZs3TUQmvvtPsrHdXza7wZQmxzIk3JQZzak5qbFZEJ+HKNtxDMNmNvrbv2ltnvyJ9BuZjMIaAYYy+8AanzSJ7absLByGoFkQNKW+ZK3B7zDPo1soM3oL/RFQAP6EP3QXE7Q9gDF9OWB33QlwJK54Xn6IH0e4IQ8U5EVjANzPUb+6Zf+9r35377lf0kfnUA5fdDnBmD8ZjK7QtD2csQ/WmfTcGfeMPd0VwIy2tiHqMCKCNmgrbp7KWgudPzK9W2/8uDRGKx2/RAI48Ikcb28JjTlzF2NYHVv4fybrq89/d36mbkBsuJ/V2KsnRN5MdAufyPExdC6AqB3TnlPim1Y6Xp5WyDrc2vp1ESUB7vR3m2ECu/qe11VfDAXyfdTT9YUE/rNxWEYJakcnxeeXM4UbRUmyuQmaq3dd2EY9EVYvMpK4HIaYZNr6CP0MywDGJcWFwAN4qel6X769uZXFn54578ysoL+wzFor6FcegL8mWsoExr6tAfrBOS1uRRCq/eyyJ/lz01eXAv+yZG/637pwE9UTlf37pcW+wNx0V+M8/5yUGTPrYZj3ymZTqpN9ythUfHl3b2zzy9GU0d6fmVOfwOG0Q4fUWIuhcxgrqaOZi11hWIb3GZWH1hKAPTTB/90WGfm2K9GXnK06rcXV7MJ5nPGOKAgMqLvMk5Zk7jvE0oXJEfW1U1dzL3RsTm0rmCtYb3jGcwNPNcsGJEz7ci8Qz+AeJpTgvTDvSPtuK4t/W1y40rGqW7/9rGxHionz75elhJ3iDickrwm60Fr38741NMv9/d9q+a3PiUC484DlRdn0jiaJi5NWkQflIVURYSFL+LxhVsbD9/yTPt2ZPzUoS/+H6sPTPxh/42M2VcU8DL+MKsIuYeizyPHgXJDXhQChz0NUb8dBoOQBWP6e1mu3jqFC3wRFlxPwgXUm5blZRS1vOSVEoCsgJgj/Rg/4Q6qovhAYzsKxa4ozlTH8gUB7Xpvym7QjLX+/ugNxiSkFO9SAP+MiT/Ic2956cw4eX0y6USHvSCv9FsVt3q+2d79nnN5EOXjcg01Xmn0CwW27oq88DvLNcXFuAjN8H72egf9y95jR699BVkhosDFtX6vNq7QKFF2oL1ULeQOqibSpJomoYiFYo8ImXMiFroDt1BewRz4FciYoTzMJepBrTv9LA3G1i40qse/sX927y1nn602+reoLklUTZ5QYg49J6LmeK9duf7cizvGLpyYuunAe08f3HXk3H4RHOYuUM90t++8Pr9lck/+s4sv+T+3YRFgXsbqi7HLO3c5Jl6vN5S/lxIoJVBK4F0ogZKweBc2almlUgKlBEoJvJYE5PInlHZ4qk8DRnD3APh2ylX3r7q9f+2wi6YD133pGde4CaAKYIf1wgiCUQKBR/G3uUKC+GCDTiwHNt8AMYA2FvsC4AOwCsCDw0Cu0e+2bzHLASMvjBwhX9u8UG42hQZQGmExSnYYWQEIZMQGmyqAM0Az6oi/a+oJeMN5QDjTcDe3S6NAoFlJWPlHNewBW6k3G1k2XXwnTw7KDYBHmQwU4tOAKMpCOU37mM0vYCnXkAf5ARiykeTZfHIP95uLqtH2ob5WF/K6y+3+cfkwrky6Jz4DMUL9AfRoD4gp8nuOvqE+kllfGZZ9Kz8ol72DIB+zzLks4HIrC/JG8rqEhjdZGKFksr9IGG2MzbGJJYXdY6QYGohof8uluQegCOB5RjqNbNohArGCQX5fUkKj/EeUAGDpAx9V4tn/rxJAM/3ta0NZ095HBdieV77tzAuidlCf3NU7e253b1e0FE6udIMq43NAXKjcWwHcXhTva1hWAMoDfjJnAF7jyof+D+hCnSFkzut+A8Yv5vnKLz/JnyZD8mOMUX+suzjPc74/EwrV9l7tQUOgqKv7q04xK3RT4N5Tf2KPAnDv6RZVxcUdTDdo4jP2rlNCTpB6CyIhXqdcryglY3hKoOpaJ6+nT63dda7ht3Z4WVWq397psIjOTXr+hcDzdguEP6iIra0gCqcVeHtZJIVi9qaag7zED3wRE+GCTiz0elllLeh5+n05CANpavueAnBvJDAvIbNLnuZ+5rE5JeZF5p1jcsFzVFrs798Rv3zszuaXFx6a+h3GrlnNWVwL2iyVXAYuov7uCxeJ6t/T38wzzDlYWdDHIcn5e1HjYqNl2OjawNxmwByN5/+lE7/gXdc+Fv3bA5+dfqFxePzW1adaUd7f81Jt/y3NdK0fFQlk3Us7e+f/9AOLf3r2rx77v6aO1udO/6Mb/8HaH85+18c1DvJEfll0TYyVjQgOWDv6PETBK6w+rsDKgrnNiEbG3Rn1L/qfDGSKc7HfO/Hp2V9cfl/zq2Enb/SPdd6z+jsXPvOrraz5eL+oQpAtycKnl8k9WFH45wXEA/Ix1iEWXtXfrqB8trYynyBXrDgoH+1zAvnShkqMR85D5rBGUhfWvk8pIS9cDP4C7acyXDJWxBslVJQfwbzpgzURY3P6fEhkxQ6RFWMan1Enqx+aic4xBu+U1UWz4ndnm/5Kpu9RO2vsxqWb7isawVp9b+XE5Fo2/s3TvUP/OfL6R2WZcVJ9c/FS7t149hYd9K2Bayg+RVQgU63lg8lEnt1y2pH3l0Rkhb1bDcaAyI5XFeE1An5vUXGv3WyG7qDMkscsbF2hluqueW7pjO/23JhFYVwwpzFesJrgXZf24p2Re3ivwzKJ+UnO/bzpIMy+Q4G19517YUclU4yKqNZ33ZVavT7ZyRQToyPyINV1TkG3wyzRTB+n0ixQdKLLewsyK0vWytc8REY4uX6qeEERi7RQ4OtijwJsf92Li7HFUxOFAoCvTe5ZXlh4aep4nnnzMwcX61nqH1d8jpMiVMSrFShKfESExrKsRs50Vqpzp57Yc+fSmYkH5cbqN2cOLXRVh1pUSQ7PHFw6KwOMpaNfPzR77ujMZxWf5UbVZ/XFrx76RX0+vOfGl6fkQot5hbmnCKJi4vC96bOPnI2/kCUDAtkO3kW/R4l5/JeVWFfKo5RAKYFSAqUErjEJlITFNdbgZXVLCZQSuLYlIADaNLIAFz6tBLAHoHmL0orb8X0fdEU/ceF47GrXAUwA7LMx4noARNtKWcwJEyh/sxFns2YuIgCiAPfYzBkgzWaPjQgH3y0/ymUubwxM2QgCGwhnLqnIwywhLPjrQ8P8ydtiYVAewDTKwLoHaAgAY2bzAB8DFXMdgDPmlsnqxD1oz0FYmJ9eysp58qTOVjY+yYPNFSAbzzHCxaxHjKyg7lZXs6ggPzRp0SwD0GNTTB4AGxaAEW1xztM21POgEgjHAHwb5mkgOOcop7lGAXx8Tm3bcQf+1h3u5M8hFzbcmO/T3vQF+sSn1Vd+g/z1OSBTNrhA0qkrPmyjDfi1vvn/ttury9uqX/Gjt+VGsxIx7XFARetrgYC3gdsbc0disSYE0BrhNCspUO9AoLW0iQUSF242C/yw1ajWwzS/P+73bwnSgWgeFrh6hxL3spk3dzIbKwZIbxZCDwnwrAqclepkeL4VNk5IC/03RFjs/5Op++79VvPGQOfbM8mFR9I0/J21sJm0gsayyv24ynzZ7nreoGStf9JfIWTuVzqsxPkvKH1IiXEKeMwn5wAu6POXssKxvoR7oO8c9inyY55jjLyKpagUyQUF4Y4kn4HrjbrfPra/cmzuRO96J7LCrWSTrp9LKzabcBPhwj0CRO8Z1hOglrEE0EsA6dd1i4N1Rb+oTAhM9S70d4Xz6a7rX+of2nuo+vxOeTIvTqSzi34xWQmk3HogyeabRVZNi2CHWroicJNIvLEAtEiuZDSWvb7nvFhAZ0NWFwuVOFiROxlxMXLw/yYOgOUhUMyY/KASc8HAX7nqPl31uvOxXOzfN/75cVlX0K9pG4gm5iuIVsjPOSXmONrp5M9e/5PHf+v8Z1ceWbv/dJLH75WsIdcYI6siZS6MpauN21afMOLYNJzNkoxryZd+Yi7syPsGkRLBXPtYeNvq4+qjxb21rD2+Ek54t6w+tfzghT+uihhYOLL23LEjreeCyWQRgOzQoc4J/2ef+nte9cZe/WtTd+9bCceTvh/v0Xi6V+OiojFR29c9tfjYF24/fyXu0kbkx5wL0XZK5dindFYA+l1qHsGTxYvS/v/qDbWnkO0nZSWQ3lh/LJ+Kzj3+H+f/vJjEJnUORGgdFrGFfJ/o5vVpxWm4Qd//P/JUerPzpK03yB15srab6zTaknFn7olo5+P0ASUjkQAwzQWdxbWy9fzNls36YEWyGZdlhfTbvUY9WBNZsdLVOOwmRXxQsWXuFSExq+9dkTu+SCA/L4JU7qFyjbNQ7qKy0Oufl3XFzjO9A58S2XGz8jqvcf3rIjiOazxCPrIGDcaMCIwt0eA2Yvb+r+XIIfuTe/z8kVWX3cGIWj+QYSYCgzWdZ46Si29adhef8ga+DNcinv2q518jsZEYr7yr/rAS880hrCvimhbi63K3/73py+O7irYfDiz16Pu8O/IO9p+VUBjgHQqFEMYm89RBgfvKo9ixcm5sPOlGThYJxJAYtPbCialAhMEOEQKpAnbnYSURCZ1rtCf97lolhsS4jINyQmS+XvyKwXMJGi53VJrqnB/FKXWdV2srklM6d+rJPcHK+eYBlfNDIk6a88enz/Valfbhe467nTecPy2qbVqWFS/I+qPSWmjM6rPXWqq9VzE5ZpZfHv9se6W2v9LoOVla7Op345d0vr12of4R5X+7CA2qUk163l849/zsbzan24cVsHzG9wveWZclj4ldR7LbqmPFN9uL3kdGyBpuZM4bvL+KVPIf/uN/tyVj9DJkW15SSqCUQCmBUgJXiQRKwuIqaYiyGKUESgmUEniLJMC2eWwIQrMZAAxnd7Tioh37XPM234WTcgU1tuKCacDr72CzocSmHnDD4h0YODEKkAGoA9JgQYGmGa6G2MCx1hxVuk+JzRWEhWn9j+7MLE8D8UcBfTYqpmFrRAbPJm9ABzY/bBTN8gFxGrjC87iH+lIXs7IABCNfABrKCWA60H4c5st1gDXkQ0Jjlk2iuW2iDgCdVjaLLcCzOD8AoYefpnFvmpSjZvxG1lAPQAzy/y9KbJ55Ps9kg2w+15GzWXsAkluZIEkAu6wcVm6dGpyj/ZCF2vnOwI0/v+pmPjnrLvwO58kbGQKiUUZkxWaYcq6KrHi1yie5XvmBzMxlxkCTf7v9i195US95J+1mGv0WUN1cptEO+IW3wOJfFpBFH2tTTwFEyJW2a6gH3+cq3ph60W7ZPo2lvv/D6oH1fjV6+ezumZm4m0zXu2pyxSnw8/wuBSpwFQVpdXl+xE/UVLaFX4ebvqJ/Id/oQ2ixt6Q5frjvxU5EhJOrnKnHx987+3zj+huXoinvl/f/aHU+3mF98UEByH9VwPRCNe9+PsqTn7/13/7Xxx7+7ActwPtWitBkB1j6A0qQFt83fMBPjTwIYBsNUsatEUFrkuErgHmBj9SBuQxACbc6DynZfHPJcgsIXRGAfDoqsnoop9xyFZXKmmJO+q/uXLFXBMaa2xmfVgTsmmsWoZrgopEVVjD/RIk58q8rPYGLqNdyNXOqNxeOBcuH9cz7a3JX3+9X6goePLacTgWtbOLEQlF7tumCtbBwjTjPpuXzXgRTKjhLk2+WdwM/WNO5cfnA78pH1Eq3l65WouBCtRq+mGXueKeX5BAbrXY/+8yDh98MsMNcAeF1r2TzlOflZ2Kvf7sA4eZc9dkxETqLNzcenRJYTP/Figc3QcgfSzrmIkgc5kaIYObUr3185tfPK2j53j9a+sRYP493S+t2v4IjP3nLytNfk+XDjpvXnj4kiwdFne3R1owhiA9Acr7bHGfz1HtFMuw9V9nZU/qU+vGaiIdDxK+tZ+2lu5YebqxE4wd3dc+mt64+eZsIkbtUD+6dV/8+r7vu+QfP/qP8Fw7+5ORCNBN9Zfq+uBXUpw92TuzR8x//q8f+xdMaK1O9v7zGnGtzrblKuySgPALsIgvmU9bBSC6LAsmqqXE1IbB9eUf0sru58ciYAHjIr48p7ReRMbUrPt340V3/5z97qnVHbT7ZfcfznVsa+LM/VH1u8YnW3dMiMG4VvnhBfQbSordxDFyyk2/4QfMQ5cNaCAICiyzGzDElxg/kE8Qg870Rg4w1CDosLFgfuP+PqJsSazx1IMaGxQBBZq+Q0xVYgMRymXWTxuJ75Jptt0gJ3h/Ov7/5lWJ35aX75/u7bpGrtqgqzF9kzoWK3xENmMpCsPCvq32rp/EanuvvrRzv3nDnhWSXzEkj3LztkfzXRBjOidg4KZkT0Jdyf0tpXuPX4k5s2sYa268p4k0syAbrr4gLxpO7rubSox2Xf3Tay/7x9V4uiwl7zltKUozEMaJ8vI8xqfEexZxMP78UIfya9X+H/8h7Ee88vAuiCLDPD1zamCrC8dncNXcUq4oBsaxejay+KkkxVhjjtC2WjhDszF2sCxngvoiHoyIsdomECBjHAPciAxyBvEUIOJ13slYIq31pK+Ti2/yc3ws9w94/X0+kr3D7tMnF5MM74bgsHiKsLMJq2hVpsRbXk65IjAkRCyunn9mVyWVTX+U6J4uPQzI1axWZ/4wsLD789H85QnyN56+7++SUSIp0bb4Rzp+YntHnYmux/jmRMj+u8/uxCumtVlw23ZpSZ/5QW+HjVf9xI14GJEThzYoU+Yzqfmxsdq3iVxPkzbxyLIzdGZHxE5cYCKwByJk+ulXuDl9PtuXvpQRKCZQSKCVwlUigJCyukoYoi1FKoJRAKYG3SAK8+ANUAI4TlJRPgKZvuXjPlEiLNbmFqmhDFrsgelDn0UxmI29m54CX5iLJAHmKzkYCkANCAyADEIsNFSAjzyQuAmsOQAkbZb4bAWJgPvkYeG8gqmkgDrQSlThv5yzWw0s6N9BmHJZ1ABAMz5GfaaCZhi5/Y75vz6Us5GllAxy13/hO3bgHoIj64QufwzaraIdbcEQjWfjdCBMry2Z1sT0acmJjxj3Img3xieFzcNVk1hz8hvwBjpAf97ApNW19y2/U4oPnGuFCljdK5e5zLl3a5eb+zrhb+ZPHXbIwp/OAjQBW+HOnb5hrqy1xDXQJtyCbanUO6301fyBf2p+2oO0B3iEocHHDmAGopc2I3wIgSHv9ygMLX37pf/6Z92du+dHI02jr1aIxt1p8b9H0vydw+Yw36T338vTMwWTRd5tBiyoAACAASURBVDPFyo5zN/z/7L0JnFxXfed77q1be3V39b5LrV22LMsL8oIXREyAAA4JEwJJIECSyWTem5nMZN7smeWTyZvwknnJvFkymXzCg+QlJISQgRBgAIPxAl4xlm3ZspZWSy31vtdedW/d9/uW+ojqtmRJHmeCcd3P53RV37r33HP+Z7vn9/svXabqeyZblhevIDTlaMy0VUvVntmVWDzjVzPVUmDmhM7lAn5/RlDJpOM3NCffpeeNSWP8aYG7yen4oPl29maS93tbf9bUnGgmHRQInblBxiI3YtL+HpDFxU/iA34x1vUff+3Xfun5Xzr5m1YD/koA28u1G2OYccR4xL3V+5XQUL3YwZjk+MdKAKPEwvm2wMGiNPcZ73Z8W/CVT2T/pssVgt9VmQeUQXeyXnk6Va/QlkflNuap4fjET8m6It3hLZtuAczT1VHTHlkxXqSmB24QAaDzmBLa2q5Az8KlSIulWk9fNYyNFoL2XgUCBpCtCLQGTHXW/I7peqQ6VQqdlURUiraOSctXiGTuriigNq6eFLrCnahV/SGFsOiRlcWcyj2hgb22UqitidBYrpareVlhlLJtiVdMVqyD2Z2qI/NMh4IXD+3PPPENWYGE0kxP70k9u6vTW6gnIkXa7j8qIe/NByQGB2AUAN5k3FR+8lDmS+/aa47kvrzwN7x61cvIjqdX/fNdX+h/59CxzO6jqaCwuLNwcqtIBeRpyVc0gX9ZiTGGq7A7iDWi+xoxR/ors+aW5cfN2cSI6ZLr9O2F8Yz6rslWl801+aOe+viQ6gJ5yBwOkN6v/x2RFuads180x9K7jVxHmflYb6Wrtji4b+1IRvmcEsGX0VhYVVmYgyFOuB8CphFjoOmT/kdA+0anWLdO4Xn79ZydAtuPiqihD98l905RuSc6fVPbw+8fiJ37GzrHdRf6Pf1K1/+bG9seURyVhBmInTUvFvebZb+3W2D8sh40m3ALg+o318vt0biCSC9cLcm7Xj7GHkTDDqVtyhc3VRnIOy0Sx4ac2ult1TX/7oYreuP88gcONuqre607KtqXNeGwEu8OKDVgoYml0YNKEKWv2NJHz2GtiolQuElkz/Uaj4P6XhuMTab7Y+du6InOjEEkymKi0RSS2aCuu7DWigiTKrsau55qEBVyJaXvCSNi0NmderZNcS0OypLtoCyU3ql6Q7zcp0R8EdqXfld5FawtrCUpSg7M/Z0iKyB81r62FE4rEdtlw0TyStxm0UBXeqwTFc3vQ7zT0BdoS6uowad1T3mlWb+mr0NzXxWwMaL4zrurCAa9HC86Ihdc07/HSaTazdlUNtymaQcinPdHruUdmXmOdwHy4H0xJyD/K3Kz1B+J+QfT2VJ0afK7Tc2SKzdRZvpYvyweyqZv+6IRcWCWzmaNXC1pSb4i64rLyZx+zHsxpEUlqEYGS7mEHECWZKXnGLluKuiZs4ovkZ472dsrMoV393aRFIxj6tFQzhGBckDWF4/KndXZSjG2UCnEHlEZM4phcZ2GHvPi+hFqngyTImB6RVw4ipexIBJjSyRWlkutuKmLqBERImLGOVxcSc6K5BiQ+6u4CJ0uESULqWy9/cA7q9NPfib2QK3sbF67/5Ue8ogS80uLsLhcy7d+b0mgJYGWBL7PJNAiLL7PGrRVnZYEWhJoSeAyEmBDAuAA0ARowTpwXnMyvScwpQlpY8VKJr3PWh7wiQk8G1sbj8EC4ABA1nrBWhmwUQKEsZYPE/pOjAxrvm6tJ7jXunay4Lp1r9QM9FtrCksgWEKAT7vZtuAWhAIacpYQsSQHn3YXaC0mKB/nsQThHuuewYqvGUzg2s8oEU+AzTz3oPXLpg4Qh40bQL+1aLAgvH2mrcPF6sLzuB4AkLIhFza9aLlCGAB2s0mjvdD4BQixhEojmKcOWxc2p7SHlUfzc3kG2pNYTQDS3G7cxKopnSgrwPo+M/OHNpgz7QQIS14/q8R5CIyvrz/rdfuxSYOWdgDwsdqof0vf36sEcEF/wD8zbYblAN/3KSDwPcVYavzR7bedG12ZrPT4SwdC1/3fKgPRe+JJ3yx2tJta1us/2rvFzwcJr90rmhdTF8XxYyPVedNfXYltK07XSqloOTNfinX4+cFIrr7X8cMA+KledkzJTSbXIm3Fh7vvSH2t5x4jbXLIikYbyu2T6a0uBHlFbbhYo4roeL+CFHt5L/3pk+kdz+4onMRCBC3qS5IWV9g56NeHkInSDyhdiqzYnB1A0p8q/byA9KfGS3tntyePMgYh95Az4DhkxXcjaV+8QKc6g/x9cgfVIauKlbIT+8bW6qyC9tT7YmHtm0fr135JGtpzOT+7W+55jrZ7yz8nn/lDxXpaICkc6UuOT+kM2to/qURMC/zjXwBsAWCvS387O1mZf8NqobND/vRX3thxX1b5Jqeqo6flwkaGMtHJyeqWWi0Sq/WXK4UBedyoh/WgWguWUomoH3WclKS+KAsLx/f9tXrdXakG9dNTfr02E0ajp8Jkqi2IlFbVod6ytPCK2mcdzIa06ZRmeyit9RkB5VhUHDiQeWzXmfLOdoG/79d5TXQNIL+ZrMA9yuZ2pD04Rh23/hCz40jy1JEfinz2zGww0pGtrCaOOtdBqqVlXXHHYqxnckdh/Id0PfP637yInBtkBa7NlqNZ80T2oFmNdhj1TSOyw8iSwsitGVZEZntx3MhdlPzZBcyp5Get6RpzMuTA1uJpczy9y6woLy+sxc8mRErV1vacyOz8O4of23HLilTjwyqEI+AkawTzJnMhGvl2PWI8BAKD1xQE3D86/Vnnkd7boqtyTVVTLHQRX2YwPjmsfpQQWTHaHz23v9NbVICgiyuxUy4B9ArB7JudySNG/SPIV9qzXdH5rM47con0g4lIIVsM2h4QqfHExPk1+WoO6g8Zxfq15Mq6SM3SIfpnRN+DpBMWDoT53pu8Qi0dwxNZ6H/sy0f9m64dqstSgDWe+j6rxJhj/LLW4C6RuRDSzh6shVdNnK2TFR2y5tmhfnZX3KnsE6DptbsrCrQ9nVX9Y+qTpt1byYnEaFsnD+37gnWBJ0O1mpF9hSyifLNS627EoIG8wHIKElKkIURGXM95q/JAOx6Lno8rMVc/pDG8+gpJC+TLfMrYoM8wP0Ee006s6RDbfEKO8CyI4Fft2BQfyeZLmew7EO8HNrYR7zy8+/E+we/WreTVxOR51cr+15iRfaeCQIRcahzEr1Dfm9p6YxC294auFw93a+Jg7FjlHQB0xgEuQHlv8gX8l7GkyM2n7/GrmszL3sryVEdFAH+yedWENFBQaqNg3KZaijWsL0RwYGnBo3mfs/NLs1h4BmW8koOMGJfUZ1bPry6fza6KJCinFDtDAbLzCvAdXzzdFVE5WTt5z2S8cg8kMdYPzPGuypacfrHvTtV9q0q1IkJlRTEtyuoxfepYJ9xosNOLBQTjNnJzZcqF2ElF9p6MpatvaO/Nm7W5TKOOXjQwrhe8IdNduE/1d3V9oLHHc0VsGMXLCJ+SJcvKCk70Nq5gzN3MO3Vijcgt1Cta365EaK1rWhJoSaAlgZYEvvck0CIsvvfapFWilgRaEmhJ4K9SAmh78sKP2xjQN4AmXFcI1tkVmo6DEeP1xExiO5sjNnI24CbANRs1NrPWYoFPACE2xMSQYIN+VAlg3QYhBGRkk8XG3YLmbJrZwJO33ZhZcB0Qnjy5xpqAWzdUzUQGJeZ3wCSuBSQGPKE+bILspqbZJRP32LIDmrJhR8sUoAVwzboosgQAdbZlpg6gTBakY5OP/N63fp+Ny8EzLEBgiQvAS+pL/lb+9jo+7XWUDZlw/4eUIEYAX9mw0R5YrFBPEGdkQl5s5LiPdrGxQqwbIs5bqxTrd5l24PyC6X//GTP/56NqdyChsvHXaF/qASAF+Egf+YrSZYM6UonX0UH7ICfGDYATWv8fXK8/4wB5sennAED/TQGnQwp0/fdOpnZUT8e3PuBGQy+sOu8OMpHBufYu42ZD80LbFnMm1mctddSxbVz6l0r2XKzHrMjFk0CDaOqaSjTYEzUd1VK7mw/LzqpZdmphzlkwscV8T/Uvuu597vHkLbf8Rd+9Bs3y5mNe7qDunflLUxUI/OU+PGFsPAQk/9iT2YOZd8x+8UERHJ+XxvoEdZZG+VWDkes5I7c3K31YCYsJO7avtPuoz4c/I//0c/O1QWcscXyrgEtkzPj8GaWLafw3550XMPs7sqjoG64troqoOCfS4ojapjNer2Y7vdzRPzWjRZEhn8wF2etW/K7Kmt+ZkyuZdy7Vqk90efP/SLEILlZWLEUgrAgs7QnwnAPwhAQQ0Ny3UOvfo0E+vOz39OOuRtYKcQHYM9L2/saR8s2jlTCxKLc3AIaVr7xvR3j3Hz7BXLGkuBR+I9J2zbQLLnblVz1S9espBeUmMEo150TbJuteW0kxSlZNrDTrxs3JRJo++Eo0UV0Bve3q3EMKbCzgyjkn64BQLoxuF+B+/Uj81EHV3RX4y5zDXN98XBGI5Cecfc5Icd/aRFvOlCJv7PdnTHdpuUEynExtv0UWDg3iYZMVy4XnqJ2MAsWbpzpuMo913mLk+om4LEb9siaCIhTREBvGuiJ3VCRGAwu2JDhz+oW+JssJoxgYZlvxlEkEJQm6q2GhUYykXbmD6i1Hki7B2UWQvEFlYU2ivljWkem/VMLtFXOzJW4if2/8Pz3x+1s+FD3bMbS/003f6nr+qsC+PX3e9DWpRP7amFM2UbfSICQuVT9bUQGCohHXzO3tX498O3enyuEa9cUxWeaMycqgXV1hRW1Su+7+33/sL9/8oatx4cN6yNq3W+0cU3hfYNKjURMeSJtgdYupVvZ61Z3tEdnxOArhIvKzWvXLE+eWc7/fG9TkasxXnwZox/yC9RjQFpIL4vHQujwgdqw7rSvqF9R7naxgHA+r/2W6vIWCxvaCiIqwHCT3iMCIyGrirAKrj8gVlIoHfbUh+wuEBefbI8tGYZJNtzdvYhWRQCIv6nqlWfOz+h404tJknUWRGz5rOVaSDGzq8itKX9YYJr/6pSymNhHY9v2FtRmQmPmA9xBkzbo9rsTkO6aEcgNEgSV5XhWLhpchK3h/sO9uLCookPDugAb+59bLxbxsrYdojtfTQZsB2gPS02aNI6Kz227xFwevCeIiK9KaMr6s7oMyB+7y6CcomTAvkNYU8+GZoObeLldPW+KZ6pisDZZksXBEVgpfrBajIomcC3mTPySFHDMpnVcg4LhMsO3LkRWWWGXsMTZZFyFXadsVWVT8ZW4+M9/el+9UsOzt5Vy8sDLTviTyACUmq/zynL7bdxfINfrNh0UuTDGkNC8lvbjvyGrkdMfA2tlEW9lRTIufEyGdwGpEVhXFVEepnB1e3aNYFQXidhSWk6aedxecuE+fS8vtVEV5LMkFFpaoyI7373jgO8e6t9Qnc3OuXGVdEIn9wvsVMdVw4faqWPy+5AmtEy0JtCTQkkBLAt+TEmgRFt+TzdIqVEsCLQm0JPDqS0BxK9g4s5nBjB1Amp0SwCOf8ya5fdBUV3ImsYPNDpsj67YJsJyNt7WssCQDILkNygt4w3nrXgmAHhKAjRAgD1sQ8rQuljZrdfM7wAsbQTby1n2Sjcdgn9mMUHA97pLQciNvNCUhLR5WAoAgj2Y/v7au1A85AGBNKEFcAMKQjyUrKDfXsOn7pBKbU8gNgAnKRzmpC3laEsSCFjq14bAupZp9ZHNtM1nDc5ElGm6UC/nwP25QCCLMeWRMeWw+VnuYvKy1CmUBDLEkA3UlH9x0sDnEfQHXRI0TlZP+Pb7xOuImtTtj1p6knW2QcMpAH2FT+TR9R3EskMfr/bAatAAcP69E/AXrtgjZNLMMtO/XpY3uC2i9Rb7nu/Q9eDG268ee695TfIP3zNBSvM19sm+PWY7AI738IYDdpOplczrWbxQo2uTdpJn3OsycNMSrspp4U/6ZeI+3GpcDnPY+f9XUe5wnHinfkfyc9+5dTzjnvfTI5/9LHpL1V0xPZV6Ochzzld63Nn5v99cE6BbMVGLQPNB999vPJUbevjf/4p6ym/iY4ls8KXCs8gpIC/o4BaBPWdJtc3nQPMZahTnjo0qQGxsONUBvOrK2S/7p+2/IPLIl7gRv1wWHlOw4vJggP6aTaFDfImLi8X3l04NbqnOFdL2Mz+0e1X08IkRKlheVxcV3lcdjqfmS8SYFbEYmK9seE9A81+tMBwJMf1kuaP6+8mluc/u8X9UX5ojfk/a7v+MLh1fPVfDL7ewXGRER4I/FwgG5mpKWeG1Vbm2WpPW9FBivLPAZ65WS3MI05jfc8PyqSAtZWEij1VTk2HzWdZyYetKsvre5xlmtJRI5+dlIzIXe7jknpiqE5RU32iHnYLjvWbJ5XUwYm89BrKheSfn3H5VW+y0qE0FW2/pi5xKyLHnnot/XI5c8CrUiasRIVf08cXpBBsLXXSnYXgCML/VMgGSRIGbAPdcWBCkzWJ0xXdUl80DHoYbLsgNrzxgFzcYy4qJZQE7QJ0+kdzbIio7aqrl9+VGjeCsNABsCAjdng5Upm8cFAlAZMl9fOHAFdcPq0w3Y+xNbPmxkFWHWRJykg6I7F++VJVJM9a26ys+S0wxS5sVfUnqT0huVAAQnlIY0LsbfPffZ3EpXJns2Mnjz6eIO/3h6tzOTGLlm2J1QMIuqUQwT47l2ybx0yzTAeAmV65E7Lsk0d8g9VLd8JZXvkpuoJVlvZAdjZ8YFrM9eiTXAugUN62mPxpAsikI5mQ+qnU6Qiof1VNb4hRudSnnIC2Xh4O7QdJBXGeqBHxRW85XpqOKlfOqh8dL77spCxLH2smZysMYAliIf+gRxMegfuFm6GnCRuXW7xtweWaEsKzD2oOLHXKNxM6z4L9FaPW4Ux6O305lXvIoaQdU3CxAFggsTKVYVmifMVGWrWar1NlxDiXyU17wIVi9aYAMTF4EkcsQSH7i24viH6/WhDsS2CDaTFhchK5AB8w/9DWILUBtZn1ICZOV9CItWC9Ay3nG7iHxYm19tssAqdwBW0yaA0ihAAJpTRp6NC0Ni8DDXsm5BYNhYLecl8fo46Ei89zCmmb8bh2JWCGx3R9Zm3dOdI0FGMS2Q6YQSaz8y4z2acaDF00BonIsmfMUZcmdEBgwpxgOxK/JypbRNLpU2kBX2GS9DUDAWruagP0EwcNh3XkhFLP8+oMR76lJuIXP/sYe396lcB9Tp10zdmdBnXeXnPRrCnEAtlJV3Tt5BGU/0E/t+2qbg3ZO73niqLGJCsWCcYn6hdFjzxKDqXZKFRb1rZIVx0C0i5KysNxQDyXSlssU6AcYV2+KobCsm9XwtdA5jmHJ5umbr6PX+Li8WHj13JPKYX3WIQ9V8YO1LfC7eh69mTrkaGbaubUmgJYGWBFoS+B6UQIuw+B5slFaRWhJoSaAlgb8iCbC5ereS3UyDCgEenicZ1p6ump63eyYoxrVbA4BgE8fmYEyJe9nAcK0F29kMs4mzFgQABmidcx1auAA9gNzWKsNuyiEIAPyt1QGbP/Kx1gV2s20JgIuRFYjIkh5WwxQtT8A0u6GxAZC51lpKWNDKWjo0giQq8Uk+lNU+F3ABrUg+uZ57rfsAXEFZ8NrKxZI1zdYdXANwQZ3Iw7rOoky2XHzybO4bW38OMmETSd7cC2GC3Dj4zWrK8r8ld/jO82g38rNa8NQP8gESBrmjgd0v+3zfuOkRE9bKpuPWLhEW1JU60Ce4l3KzcSXPJ9ef/Xr+QA70ARLgBv7bNwPXtA1AwZ8IYCwKeL1dG/OfEtA6jBTj0hU+bK53/ij7Y/7xjj63L1w0K3LNdLlD7ouMrAIaBAVkhT1kkXHh+/2ZA0YWA2o419xWOGpmksMHP+++0zxRsyEFNj7l+rVnvt1ZW06PlCbbFTtg6ODKE9J0bzfPte0TcKvQJkr2+J2xXzC3rDz2oa7qMsTg/01/uBrSYh0sZb5APviMxw/4xY771/seAAwWE+9RQqP9gnap5HnrWtDVPWxOPymN6R/W/6lLaKwzDzB2fkcJYA6w+Vu9/urZsepMLlGvCScJM2qWsVo9MS2g/+ycv8N/X7bmHC/HKvK5vaLgo6tni3vK8n///ER5V/uBzOPP3dz2cE73QVbhEmfz8RGV54y04eXGqVoUQYF7mxuG46eTUcdPVsN4TVry56phwpUFx7wsRJxT5d2T0voubCYYRFowBqsiLhi/dq5hXl0MNGiNomu/GO0qz3qxxYIT6a47jqs6MGaZRwPJnODkV6p9H1Mg4qwsV7ql2d+d9Zaul3b7FllX7AkUbFy/NdzsAALroP8DeF445DdkcveLZ79WTkQPnhvp3VWLSrVdLobEorxkn0E+I30nzLMdN5vp4nWmrzhvKnKNslLPmqVo16WtK/QLbszm4v3jT2VvmjyV2pbanT82thjtLh9avD8qgm0+W1tRpBfTJ1KKuZMDUB0NXsYqfaHZEq5BAvRV5xpEx1ysVy6llhrWHi9krjW7MicUB+P5dNovlugnTdUFGLTgIOP/Dnk4MX4s8ubFdKc5Gxsxy0Fn2Gvm5M+r3Z2pjbi9sWmTjS8aybfxzPXDWr9RRlxPIVPWSNaWQ1zTkFXilKwruk3BUUh2WQaIrAB8f3enN/8mxXFYUjyL39elgI2XO+hDHfR3WVRIksGx7aZ8IhOGB4ZMdXIwEiz1xeqxuOuOKCZKphYEEbkgI9+pUrnWJfbsxUwqPttEWjDPsdawLiFvyo/CAPWBMMfakrpcqTUWa/eQxs0euXw6q3HSIyuJMdw3VUVWiFCT/AoqX5lxa+tqLWj4n3YGoGW9nsIyRpYYNZEe2+aqg2nJDXdsuj7cRZ/WM7RIRsyOxFFZvmyweoG4eFAJ4vQvlCDyL2cpQv8A7GbS5JNJHQLgz9frj2xYd5Enygf0Hywx7DrNfHelY9XW/VKf9HMbXwkFB/JF2QFrUMBsCF7kxvsRbYi7R9qJejK/vG6O9fgVlmja4EpQGv8iLJwHq0WTj3hmTEMc8hzQnHdE5Ms7GCmmqckTEL9LwasfFFnxNpEUibkTvaPqNO8TWSHWT9Zal+tBL5V683vv5QgMOx8158L79ZiSfUf5CX1/t8oiEiHslaVDXyRSPyX3UE8oNkVC55nXec/cTK7wPsg4Zw0tiZRJybWTFF5ChZB37lM+e0Ve7Nf5flmTVPV/JOIFDKiprkRtQgTHcVlUtMv6AkWaRQX77pd7qEmVgT5I3li2aNoRy7G1fn9bT/2PS6sR3jub52qIP8ZUUm221nIL9boZoq2KtiTQkkBLAg1gonW0JNCSQEsCLQm8DiQgDfmcNOVBOAGm0ZoCIGBTUzfRzk7TeWfM+LkluQfiGjYHEBB8Ws3/sca15wF+1o9GgMr1c5ZseIFNhRKbQAByNlrWasKSBvxm/fTadchaLdASFoBv3qTZ783bPquqSh5stMgDQJRr2EgC/lBW6wrEWmvwDEtKcB2berQc2TxxPfexced6NvWAq5yjXlzPvQAU/G/JG85TbmuF0lxeAAT7f/P35rrwXJ5n5UGZKQPtw4YTUAiwAzlzWJ/sm61e+A0ZIAv7TNoIsAT/67jostYb0ouOK99IybTfIaDlvwoUbvgpB2yy7U5f6aPvrD/39fyBTAGeaBsb1JIg283WQoDxy4qHcHaXf3wxXc+PLrg9w6e9rQ1AYdYdIFqweca/IdZdPyeta9/EQl9Rb7/rFsIKOCot85qCC7cHhUq/vxLPyRXOymUsMSZiAw0NYlfYw9n6DuVLN/nuMeaezkm7cbmjvvqJ+WRfSa5wrk0ElZxc6OSl3Z79yJmPv+2Rztu2fnzLRzbc962u2+Xvf7c5WHsCwhNikFgDh0ValGRpcXF1+I09hQrSr+jL+J4i0PbmA8soEkAn/ZX+i8YnfZLrkX2D3RFIu1MkwIiUQxNoyF+CsMAvPSAmbi4APEhLdxSO+AqwzdzUJ8KjEobuatnpaVsLt81/2/3FlIJWu2+LB/VCuTb7nYKbEeie9ILOwkl5tFiq9Z1TPIc/F6gK+PJz67Kw9ZhSWYZq9dg/n6zsqEgD/og04kVU1PZIM1yWCimFSE8JxHT82erwQIMAUKSRU6U9DbJCxMRFRNI4ZQkL5gtkcUFFv+RE5AfczCiI8JpvHOuqCXKHexJYWuiz4WDjUkF9D37lq5HZ6lSvfPvfKED4GtxAZSK5PSJptuA2ZyB+1vRGZ17iyiiTL31TVhU5gfWRncfPPr7r2NnBWLW2p5yIRaaHJKvuNm++TxrtQqJy7d/1/IXlQD0TyFKgaCbCHSaXTpmBtXkFZk2YF9qvMRBnSblpUpsiY8BUtHHXFmPdU58e+rGirITy/ZW55/KRTI8IjHfNxvtWpxJD3xFZ4RcjSX+kdK6o66k/8zNzJjEDIKTpe4xVAGXWizGl9s7q8hPXrT13nQiQW/fljkROJ7cED/S8qfJk9g1ed3UhvzU441zK4gO5QlYU4wlTSCXN0e49ZiXZYTKpJSfs8b1twVGh/WOhLFccYi/Y2BXxSu3FRKnyP6qxaHs5GWtTHwMgBwxlvsfNEgTAiGT1d0Ug7WwTuI6VBWMbl1Kj8VPKq55d9bve3OXNfUtWAM/905Mfv6B5bNu6yRLArndZyXWbKKhomwlGq06kQ1ZGme5YPWiPmI56rd4v+5m6VoFU4NdlZRMuJhIxAZkKaeK6QVmBU9JJd+aLT52rvWei0Q8ZR1gUoMGPlj7AN+cgLSAOWIsa0bGbrRIo3yYrBSaqLSqbp6Da83tTTw+drWwbhqjZkjhptiYKJuOtms7ooqTd4D8smMucDDGA5SDyY+6gnSEFnlJ+gYiOa3pjM/smyrvfInlpPQuXZPG0LxkpZGarCtbuLRgIpU1zCOX5uNLfVfq65DsuK4vypjJTDuTaIFqUeE9AJpSBDm8BYNYKni4dCAAAIABJREFU3qlQAqHcXIu7Ra45rdRw4bNO6r4E1r7KYNy8X/BuAhkC8LxNCcuKdyoR6N0edmHAWoD+huyQ2QbzH83t3+8H71u849FPv8vQq1UB0Mdu8j/du71+S8MK4bsWRMwhlhBFPn1q1RlXAaRnjvUdEvC/U4GljUgLtXbjFQyjr6s9ePdmDrPWxlfrOpF7IRlYq5s1IsT2hWlPBoAiGZx0Z+mAF69NKZbGQ7Mneg/JKuIevR9crLTMpVg9zCqI9tTima6gvTcX6P6b5RoqL+JDBIZiH3n10w0Xek7jXbo/4tWHFOib/AIRGgU9O4V1ha6x79CMEeaNgu6ZKC47pyTLEX3fEPNDv6McAGHEeHlAqWVlcbU9qnV9SwItCbQk8BqVQIuweI02XKvYLQm0JNCSwCuUAITCO5QAvgEX2NznTffb202ko2KKR2vGyQIAAHqRAB7Y0HGdJTjYbLAhYmPMJ5vcifU82fSysWmYeivZuBCAGIDf5GNdJFmQ3m7u2djYzZIF2/m0RIAlC+w1lvSw4L21dKCcPAPQk40T55vztSA/mx6IAK5jg29dZHEtmoiUC7CFstu6WgsTSwgARtj4HPp6Ibgl35uJF/tMzlvNWkt2cI5ncx7AgefzyQbayoS2ooyct5YrlNHKxGqxcj2/W4AKmVsCCU22hl9uJQgaxYXNPm0Sw7ebquKvmjp1s24AkAltNab0RQr4130IPNtcBCu/l9M+bL5GuOBFN+MvqdolgCkAdzbN+ABnk23JH+6n3wOMPyRXI4s/kfuTw+8J/qxnPLZt1V11wo8P/HTtWefABVaiWM8Yaf2ansS83M6wV99YN1kATGhP/82aLJ16/LWOHn91vwrfNRBZmpuM9k6X3djNBTcB0bbhIPCltPjNV6O3m0qk23y1+JYNv/c5c23XRo460l6+/WnvhsdXg/Y/yZTyJ/uCuaKA24oA2v+meAAfkn//n5cv/w0udD625WfM1tJpM1w61+aF/q8q499QekqkxdwVuIey/REA+dBF+hKudXAh84gSIHsdEF/tMC2t/jm508Jy6wLwQuBi+fZP4C5nVIDmuuZ/c7bMcwAb+L2eUALMb4Bxff6KHUOyOnJG65JGLdI3e9r7cLlm9nXUakHvPamqX4iHAked7EwlSPc6/qnFelu0VO1256pDsyIjcPPC3EHD3XPem74zJPJDjv87owL9fzHnd/yeyIqMzreXg1Rmpjq6JJDZk2b8/tH4yUVpfk9IKItNbqAuIpYLpxqgj0iNDdrqD/74WGWdlLAu7qyFBQSZJS6ZOxpE7joo2sjUPvdEcV9GwcRvVd85KILiZsiVvalntijQs5FGesMtEdrtyDhW9U8EEbc/VSyf3H/45Hj7WnFLtFrb272w9oP6zdRdx2RyJZPOl8xaR8aMnp4zkaBuVrNp8/htYNrnA14n5Fpqa+KEma8NNNz0ZPrnzTH/pu98LnZvSe7I/vs7Zr74mAgIwKlSKZKMPdJ5u/uZofcQu+LW+VjvlnhYGVZ8lS6v7k8+137d2Wfar79vpHx2+cNnPuHLNRNzHHO2bWdkx3zXzArSH5OKZdGnWBeZdJDf/WjnraGC0yeU/6nlaNeOmfhAOFQ+N54JCtXeyvygys24b2YApzUmByuxmDnbNSjiIlI70zEcXejrMCuKkZ6USzWCPCeiRQXLzjUCtiPDncfP1YbPzg+L2Lm5c2nthdmBrk++sG/sEZ0Li6mEk2tLlvNtKUDvnXpmj4itd21LHLsR10YKzm4E6DdcHYlQIoD0j2pKw2LgvR/d8ZEXN7su2kRcRKXnLbDQxOXKpRB1Qm/A9dNyC3WNH0Zm/KDa7lRrAzlfYUrUjIqT4kejbk6q4a6ib0cjUbe3Hob5qBepRCLu0iMH3aoCcbP+QQhBAOHyiDUJKwfkzXqD7Pl9g/XApvm1YfkiMidUX1u5tf0bCq6d+6CIiR01zWWVetIfjJ/xiElBwPf1w875WKb8C6VJJeYr5hcbB4v1PaZ85oU3P66YN1OQcBqPiyIuiE0TVb/2+2Nn453ewi2brCzsc/6TvvyB0q+ItJgw5iMbYlqsx91g/ac8zE98/4oSawWgttXax4ICCwZIDd4diBMFmYCMmJcgM5CZjSVgn98gdq6QtGD95rmAu7y7AHr/TSWsizh4v6AM1m0hbQKhiyIDn5f3VXahVK/9L+vWFfQZ6m0tiRfUkj2eZop0dz3X3lffW845TyuGxX7pDiBXawXFO3HzgfsnTwGl9y6dlYtGWYwRWPt/4qAf2XfnzRmxlm1+/uZH2RcK68aTgcP7Qr/Gdi6RqTiKMZFLtJdlCxEZwl1Tsr38RQXnlgWG88eyhrhFxAtxWJoP9Vtni+Jx9BeWUrlovJbU9WEmcD6T6izFIQc1F9G/eC9iLLB3YM49Qr/Tb8xp2/TJXIHMeS9lHWU8MFaW5X5rvFJyOjVrNL8v2zIge4g/5uAWYfE/0blat7Yk0JJASwKvJQm0CIvXUmu1ytqSQEsCLQn8z0sAEJwNkHUPxDqQMG0Ho8ZfXjXdbxsykRibCQgNgARAcjYIAPeA2ICJY+u/cc6SF1yDRqw1TQf4Bihj0zWhZINPsnHiNzYc1kLBAknWMoJPNtOctxsvymIJACsFyt5MClAWnmc13tmE89zzdfyuf+sG+Ld+LfVkc2/LwLV8tyQHGy/+b34WZeNZ1AGAwBIMzajz5nPWAoOyWxKmeSNK/Tj4RP6WuLBAr9Xos/W1MSr4fzPRY+8lHxt7hE0hdUb+bHj57JYHmadMZWqP9Du7zJb/o8Oc+ffUjbpSb2sh0+wHfr2Yr/7HJQiJzQ9qJiBsn7Aybf60hJm9pqGdvv6MhryulLxYL4CVCQATWqm0xxmlPeu/f02f96XDwjd/pPDZ+j/P/9v91bbILwy0n9t+um3b1ps7vuktFeTyRr7UBQgbadUbgZCmHD2hCMp52UNUaumgvCCCYk2g4nNCPwR6hRPXlM4sdAVrewWy3S+Li4VBZymiWAvRyVjvH8v64jY5m7hDLqL2+06k0UYE58V9jwB186X8RjfQ+Gwfcc+ZvZEXM0PO9F0/7H3hDwfdmbWuNhmEbAmX0p8qlOUSKnc2Ofonw+Wp/hczu3EhcuH47OCPmPdM//dGzAEFRj6kHxgXv6X0TZEWsyItLqpHug6SM8bQuAb0RSN78wFRAejInHIBTNfXSltk5UnV65Nym/S/25sgZUSvmOcKN8sCQP7opVAvwATwkn4NefQZJQBvNK851wAaZWFGf2j42Bb8LhuHVCF0or2B1z3qRBLVugAYHYlKsRzPK9pAZzTSU63VexSyt7vNqSuggXlh5cTPLg3v+5eUlb54v9rmHlzMoP3OqUKQoZ37FavixtHE+DG57xnPBx23AdRvTT37LQXwXhiKnTna7i2flsuaq3IDQ2yLZrB3/bslOvmEmLBWUljREROEua+ga/mdsd+Yz/Q/3xW3onqDYmhsF4GSipl6mzTOe2RF0pDpYq1PhMVKwzUR5R+ZnFtVIxdkXdEzML30weyKQPhAES982XiIUIys29p4fmAy+bIJPPVHqSr3z3pmx4lz5rn9282zB3Y04jMoFkPDcoMxcbJ0jSm0x69ZjAweu2/gB9Y8UyvsW3k+J9Ki/Ct7/mVcAeF7h8pThYnUWF1ExQ4N3rLkTlsW9FmfTI4yXx377b//SxvkqX5p57DNfdNauk3Nxvu9j49+5OxjnbfuVgD2XX2V2afF+1VWotnsTGLw6wryPQtZqPph7QEgx7wKcXkokGP7+fYu8+jWg6uqx9SRzmu3yZqCuB+Nsag2VtDn2YaVyo1PHzW1pDcjQmcgVShHhyfn7kwVK/u3nJ4d3/vCmfsy+WLaqQsYDc2cW6+fO7Zn9Ng3777+v8oK4zOyfHmLwPW3yzJAn3kj8qvRzxQrxSjGw3VJr/Qm+rtA9fIlgkTTOQHPFebXPCx3UMO7w1JqLKxuVdPFM2G1P2qCvAodVz09CSsShGE1qDod0p7u9cRQSNpZNaVXrtaj9bDyYrlSE9m2paZ+BCEBMW7XRXrBofXxZ+OacO5i8wPtwNwqgNa5S5/7jxRuKl6b/k7DBZfImYrqHRfButmdFj//mBL3897BewntYhkN+6wGCN9/4j2rxXTX5wph5m792112kgWRc0XJ8pnr648PyJKj2B2dPUSfv8jx0zqH5RxtDyHSyHOdrAB8ZQ3gXYb3AZGgjVhanGfOQ/nDusminJSP9QOZMQ4BhXkHYS1h3DKvXLQQlwiqTVGYh5rfHyAoGPv3KDWT2vSB5hhLWI9AEvOediVWcjzr++lA/owJ2hNZYarXw6wSiWv0emY81RlmFWWhoJ77ef3OHENCkYN5xZLDzEWe4jXkFMOhp6Iw9nKN9GrIyZKj9n2YNiZdjqzg2Yy7bylBWLDeQSZqxlRJI/Wd0bhvCIhdKUYn+7YvFrtGl2/eesPZM8tTHXkF5r5l7mTPzcXV1Hk3VkooQnDwv4KEx5fPZhcVcDuruBXXrkx1PNm3Y+GZ7ODqhPKnL6MkRF9/RPcNSCbfkVXG/bFktU1WFox1a31N2RhTp5SwVE0l2uU9q+pgEfRVJSwxmw/ainnGFdnktNxCvRpdrJVHSwItCbQk8L0vgRZh8b3fRq0StiTQksD3iQSuUEOcLcIGjaqrBFYvJy00+dCCtCCXNslO3sSH5cdiX7vx2gom4lmNQTbnbJoAAyjTOrDQAL3Ig/+thQX3ABCyUbfgBdewgQE0REOauqH1B6jGJpHNnyUPmjfdbPxt+awsLIhP/TZbWnDOgvRsQrmHMrMJsiSIBev5zVpiACiw8eQ3ux7ajb/dJNpn8QwABf63Zvo8a0Ogz4uUm/uoryVCbH0s0WOBMwuw8GnLYq9tJnL4ziYP2TYDQJYEsUSLlafdHFIGtNi5F1AFDfSE8TKHTOb6tKmtRo2bRMYAxnajjFx4Dn3mf8WxWZPQyoY6WasUaz1jrUGQAeW1BJRtI+rCedqY77Qzv3EOYE14XCOy7wWNdTvOLmJdQTkgBLA4sq4h6O8AB/RtBbANHtpVPH78HbUvdXwg/4nh3FDig4vdHXdHvbr8WxddL1JwCmv4oPelJVxuAI0PrbzN9NWWp69Jjj/V6Sw9rrDF35pJdGVEQORiYe25bdWZUllxlpWOJcJamA3y1UWv3RmtzUUz9VJiItb/mFw+fULftyho93v128/SSLjxAeATYL6hzQJ13Td63zJvidyvDlxNDLiz/yBmqn8uSBn5/omcLk0O+vOVb6wemsx76W/o3AbCgszG09vlsudxBeTOA2BDPgDWARwyV9DHLnYgc4Az8vvFi1zwlxRbiYCaKzbugsBXyf0j5guL788t1PqrcWfgqDTyAfsaYC2H3MbIv726seM/I1c5v6lTEEoAHpAXgDYAhA0wTmSFncPSgUkk5Q5qVCRDd8kZaCuFPf2lWqTDVxDrZCJR0KdxSkGkO2ZqlWS0vVr19yhi+kwmYhbSifRs/tl/Xsjs/3cTApC/LP/6d81Wh96GNjjWCMi/JMC6Lzp9jzTCYyIDDkvGOQXYLvfHzi1tiZ8siaSirmuXAJcvIcbzpy+hbW0DIVNn5lXmUMY6mt0QzWhzM5YBShkTyFExNmr98uW/DVdQfZHpyEDirAJnSMNe3VxWLQ1tflmJNMgKEQ5FWVU0tG4TMmIQaWG8moiii/g74RzJrZ4fXnFdX4t6T4xMzk+O7xx+Uz6d7I45lUZA6aVaj/pqF9YHiZrnFR7qvzP71e4f3NpXmj8+UJmtPdx1B+XevhzthAw/qMRagmYucxXzL+OTDhFfDwZ9QX5afBqQ20Vk1gTQnqsd+IPrTsuS4zdlUzPkhkFObqeul6un2//9jn84dX/PoWf+yfFfz924+h2IH56VFIGxVI15D5/csqXr6ZF9hx7suCM+6w5tiyfziXSYM53OouoTmF3J5xRkfMn0ytPitolpkyqV2yBw2lcLJlqTE6+wAfD9Wna5QQD+thIBZ2irI7tfnHxy2/j0XCGTnP+ze+95KBtZ7JZ1z80KNt9JnBqsNkQVmSXFtGiLrP2aNKcBxx9Sulg8C+ZNV726V235Lj15y5xGTXs9iIyaykyHLH+irptWAJAFAbad8gklyJZ8wh6n7myvyfWa2N6KwFuvVPErUc9dlOM5ZF9jvErugPKs+z+gBGBOGVhjcB33oBLWZ5u1ohmPlAuwf0zg5ptERG5Z9ntCjesBCEDFUIn3RqexJNlsRQXBiUKCXa9ZD/I2+Ph3JtecYxMLTls67kzP50ybnOPcs5Qrfi6ePqwe2ROGkZgcdA3ItVzP15bePbQ79eyp6zJPPqiYMv/qEu7l/kD5v1fpAc1Li3K/Rb9i/sfXPhrlkKRolDPXWQUPxh5yoJ+yhlJ/ZMbn7UqQChDfgLusLwC9XAuBsIHcaaxJX9wwn9v1nU/GB2QweZD/R9fLoI9LHgDCvCPxPOZe/1KE88tl8hr/jXWPuYS1qbF2agzp9VcvYFGRrxFzKp4O9ybbTcpxnTPq+8/5VW9C8Rt2S90BWd+gWA1pvxYpL5/LPiOQf0SfplLglesVHxBWNHQzKcH7i+0PVoHlcg/gXY9rsyKHsdzpkTVFORoLyooxMdfRv+bIqmIpnqn4nUOrg5FYMKDrerpGV8peLOgqriZLtaqXjOmVUESMqZViJvClSiGrEZIsSMrTRwc8kRa97X35t+j/EY3fcZVySfl8AZnq/y7FxjgswqIol1M/Llm1RaL1TsWwoM+xPo8pYbWyQ0m6F45bWsv45XyoQEb13osE/cDFFSajkPBXErPncjJq/d6SQEsCLQm0JPAakECLsHgNNFKriC0JtCTw2peAwNFmzXBbIQvQWs0pzgOk2Gv539W9Vot+syAamxgBrVcjIBuIFtAKMG/ZRDtSZv5zxLEomdgIQBogJJsDNk1sDCifBed5lrUqsG6MICkw+wbQYZMOIM49bIjZqGPKTVkBNQBo2ICxKbPkTLPLJgtAAyo3g+/N7jysubgF6W397WaOe8kHoMQGyybQuLVOoN7UDWCAsm8+1vXKLlhq2LWS85YYYdMFSGbLZfPeXBfytnXi+4a2XX+wlYP9tO1tiRdLTli1vWayopnUoJzNhBf/W7cCyBy/2QCW9AHKD7h7wnjdnqnOaeMYREx8a5upnEbzzYL9Nk7JRcR0dacuQdjZNrOytfIlc+vaik9LYlnLH+pFAqhBXoBlALXcT11xHUD9qSfnuQZghjbjO/VqaPPraMjQlq+ZIFy3DkAW5MF1gEp80ses1cuzcmOT+P0THxkdjp27O9efOBC0pW5cTrXF2/1Cvae+EvSH855iLhjFLjD52nmDFYHd5kh1/4ktsYn/fnPisWM1z6FMR7RzX3khscVX2uB+BMC959AaOGI1vG+u+EDmerOrcm425yYn5CLqhEC4r5TrqXfJ1ckHjxYPGGl6r1fv/Ie0+c229FGTlheXLj8n0qJyg+AH6y4EIOA/3e09/PC9qb8sfrL2fuYBtH6p74XjE6MfMm9euN8ohoBZ9+vP+PqIUkYawIy3fDPwtS4/CoKl1qWO+/UDZAcAZyPegkBBZAzyk7qp7Ztr5ypjR5x0/ac/PfdzG/IQeCvXUHeYXakjp4djp0cEEgOMUnZk6VsAk5t+ER3p8+MDN01ddScRLZv+wkx4a1iq72gvm2y7/PTTfxLRiFtOOX5nyqkGbiqZK0ecbNKvrpaN26aHdKSGuoPfPP5fw7HOB89sTRz//85Udu52TbBN1hNq17hRHAvTGVuIy61S5dn8G2IiK2akKX5CbsCe2p44ypxB+V5trWbGCG1G3vRXgCCICcYz8mXOQ5OYA9m2QWwNeZM3Sh47lXaIYHHpl7m17nItGUnI6qIBvPfOLZubnnwx1bUkD0Hq/rIAuJRjdsgRq8UNqfB/KbEO/IBcQ033zS6X9z5/+tHDN+x8n2bOm4kdcLBhMTBi5uUiTWReRBr2d9e82NKJ9M6IEuXcpYQPftYs1hfmP9YgztNnnlTC3cgFf0HrdbxSVzrmxcwexjNgb3zNazuoOqLNu03ExQtf6vuhulLxnx7/6NI/O/7RBlD8rbv2z8929Aycbhu9brq2ZU/ZTWxzI9XBhmsyLfW4bkq6NbGiUdO2WDIDKwsmVqsZERNqFylyrxM6tpz6RJsYApADALtB0orUKOie4+/9868tFe7JPng4euuOfL39bSLGOuR2zExXRo3GvOmPTnUmIkXcKB3V2Mk1E2HrY5C+NqYEQBipCYFdNLHkgMDDbKx+JuZXdyjAdq+oKk9UVclxG4Vvlzt7cXdht1OvpyWgo0Iru9zA2Z6IJxZS8di0YlmU3nHTMHlDCAOSYtbFBMf/vAdQJ+ZjSETIjQaD1TSvMr+Mah663XHq8bSbj+5JPbNNVFdnuZ40cgXVCI5NH2w6mLdp7zcpAXxCFED+NaxrPvblo5Gnnj8nQzS5voJ1U31FOLo3RvxgNZJfezRId6mj7FQP7lRfL4gMjeZyHUuaSyZ+auC3f11y/ceXIC0gy766qOv1ybOoI2OLtqJfUhbGGP2f9xvGIX2f8lnLH2TBtYxN+i73WjdOY/pu16mXuIZarz/9j3tYE+mjjAkUM5DzZouK9Vs2fHxM/31KySoisG7mrsCl38Xyeq2fYy3gnehHGxWRZBs2WzJxYhWQS6hkPGVqge91rMxkRgW8h4pNcaitpzDguHW/nEusJTtKJreQWZs6MhCRdUGiqrgVVxuvwo2cf91skAHGWdEfxk3z0eyGzlrAvpzsWf8Yi7x3iyAIP9/Wmy/375qrqezPqnzzmqPqqc7icDRRw4LKU93p01Ev6mfb+9dWdf6s6tYpS4wpkRe35BcyUd13WHWui5zYpbL2UtdaxQskl6ckl2tETtw3uHtuSve+Rfl1yrVUIPLmra5bH1qdbYtOPjt0Oju0+nz36PLheKZ6nwgM+uAE/U/5RXRt7OyzO7Lx9IqsXAqP+JXiTWEjpNqGo9lV1gZS77XeGVvlb0mgJYGWBFoSuLgEWoRFq2e0JNCSQEsCr5IEmgDZZiKC3C3AbsFk6zeX37iWTSybUDQNAVWtJrC1KmAzYbUTLWht3+RxYdLY8VwhcUHgRevmiI1/m0lfUzHdPxQzUekTRzJo/bGR4HnkS5ksOGwtEyx6wKaa3/gfIBktQzbsaHqyGWeNARSnvpQXcoC6kSfHpZgWq01vgXsb84LrbVBtNurN2mbNRADPBbBG85EN+g8r4acZYIA8t63fS3moo90EbtZes3k2g+nW8uO8ivf5ur3cYTX+m/OyRIslZdgm27pa4sPKhjI3y8nms/kcZdhMePA/fce2G+AE+VsQHzKp20RSkpVYr+63RU35ZMnMnKYNAf+4l75Cn/kvl6nnlf68ufyWDLMgEAAl3+n79Cn+t7ELAIfQsuZ/iDTkB2gDQETdqBftA+AHiAPphq9wDtoLMBdQEkDNkm3kYX0iN8ZU03iy8iR/6wqKvsgYBSSlbFuT9fKjH1j75OrWztP3BkPunQow3HGiczi5piDZij0ht09Rt8fMh32xaWdcrqDsIT/+uYRbvn85mn7xL6o//Pz+5KPku4GcFPh44fr/R0X7D4fP/8t3Po/HG2AhY3VmorTz1JLfc0pa/GaitOslhMXd2S+Zk8k+kxBZsd+MyxfQBkwMwAtZJf5d4l+PPxncHH2hvhdNxg2EhVzyGAUjNrvzx2xgZIrxISU0VdHof1bEBaRFM9LAGAGgs/7cL9RJX55Qog/wLOI51NfJCtqH9uuX26D5jsjyO14o3tAtX/NGGtjN9xuRMyeItyCXLk+knAJgDW5xLkYG2DlWiuRezXc61Eb7F+edQ/GSH0sUIz1Z+faPlau+QBx3RfBRtFbzBzrr5aWKp4jEruBn1+Qrvlt41E9Eql409djaPVufLbwhKjLomLTBvR3Jo6MArecUb4BDrmbeKSuGTw/HJ54aip9+qjs6V425FcbWpVz3bKjbK/jHWrowPzLPInMbhJj/IdkWZUExp763dK13uFNWDtuq9dhAR3IxC0CcU2yEejRM9EWn5LapYkYnZ83e58+YDrl/kssiMegbQCTGDyQFcykyJ4AvAC1tDnkEaMv/nxLJMa3YF7VaNCILhUZA5LfJUuAfEUQamWGZImuVWyTHw0kF5D5V3rVTYDyyoh+QH+3HGGYOoV6AwQ+vP3PNguGvQGYQG1ioULGaQEPmPwYqaw1zZMNq5aO7/mkl+/YXQ/W/iGJTRJ5cuismS4qSG/fDQj21RZY0kl22YUG1RfE5GIeKp/Gc3MRNjpybc9rXCne49VCyCiFZL6aGbdcUPlmjfkKJMfX/ylHL2ge/9tm5k2+89oEHUj+wpS85dZuAdlMJE/Ld5Dc+k6bAZPE7ShPrbWFFgbxYDyENqdvXpSt9wHPMmBxXTfn1MKjVTTXqqBkUDl3Nm1AA4bDuymdaKMC2Lu5FN8jsJhmJRGJexM3Ho15bNBppyxUrzFnBerwZLB4gqXgWWuvMmZbAZ85Fjs1WWPRHCBRfrpiCpJt/TmOkpz2yMoTLMIgxrFOwSmsiEH5d12PVxtqA5jjg/ypkhawq3MmZ1djSSikhoqItIpIxIgYmqIf1Sk2RV9yw9IbyYm7ec0snnMTJqnH7ZB/0gp4zWqnH4+qDBZEW46lU/s/UhliNbT6YI+8WKfnMjuQLK3JjZt+RGHP0UcaWJcXtex1rUbObMvoYbcq8x5ihHzB3WqKCeZ01f6a5P2tOtdaGvNvwLCw77lqv/936xPrjcsfp9eeyTrJeIr/V16FlhcGlkOqOTHmXaMT70IlMLKngCZrFamVnslp0niquxqKl1eyNQeDsl5unhNwhJeU2aaWwnIrl5jK1dHcRq4KIAPhQcR1ktSky0gnP6ZP3lEsdtDF9JyFrAxNL1RSQuhaZMGxCAAAgAElEQVSRK6mFet2pKn7Ey7XjZXEb5dkr8uRalWNU5ehIdZR/NN1V6JFlxaSeE4+nq/MiCxacSDisa3j3oR8wn7ZpoPXKCuJwuqtYGPTmphTfIhzYPXdcRIWn+2dFUCwde3jHOdV9WHnfGfpuPbeoKBaL4Y0r0+3v0Bj7reF90xPKd5/k2ZFIV/bJIiWZ7ixWpo/2b1mba4uMP771tIJxO/vf9sJpnZ+WXKsvPryjvbicGq4UkvsSbW420db1zOrMhCxaytc1MUCsI4z3S+0bLtf/W7+3JNCSQEsCLQm8BiVw2YXvNVinVpFbEmhJoCWBvy4JbCYq2AzYjSsAnAVrAUDZuJMAJwBRAWQ4z+aWDRQbcoAgUMVmgN+6KGr4UdbB5qehlbz+/XJ151lWM/C8JmRyn9xXyyVQvRo3bsSSDjwTAIrNNeWk/Gy+AR4pIxttEpt1rgMIAUBCswuwBY1tNsUQIDyH9cYSN5Z0aSYZrGsHCxKft/44DwAAflBH8gMUYLPXDHxbiwjqbsF/5ANpwnWAy4ANlJWyoO1pY2pwnSUyuLa5bJY8sHla8IX68kz+t+W2JIQlPZoJCvKxRIf95Fyz1Yh1YUQdmi05+N8eVjbNcrO/NZ/ju+1Ttoy0FeAhViVsUK1MpV3nnjTlU31svE1E3o3Oty/yQf70FfJ6NY6Gtut6RowNK0++A6pakgQgx/YVygIAxtgA1AasGWsqG/0BYIxynlLiGYCM9F+i/NJ3OU/+jCv8OvNJfsiT/mXdZtEegDkNTe1/+3zJ+T+PVhifb1T6gBIgJv0bgIl0RIDk07cWHwvuNX+x6+z23myhPdF+IjXszccYvsZ8J73TTdarcgEVkd+o+bDHXSgv6anFMKVAMdG5w5Wb9zw7f8N38Mf/Rwt/awNZwf1XGGy1/q77f7/0Ymn/jDTmZ+XT/o8F9P5woZ5JAwbjOmZb8kURGFExiv3GFygz5s+YTrmsRw25CQz8BT3yF7qdxU/95+Q/+Ny9xc88o3IyjjccBREx69YVzedxcfL2dZkeE8C22ASE0c52LticHW3FvDKu1Ewy0EaAcnsF+B+SRus7cbeEa5jNhIWA246jhQPPyV3O1L70U9XfuOW3LmW50CB56q5sJZz+ZNl0OwvRexQ2pD/jGs19Jt6dTsalXG5iETeSdiNOJR+6daG1PUJyF5brTk2dLP1CLbp/vIJrHeZod4+AdvUXp7Tsd0+fKu8eHYlPNEBrAlYTrFr++AdU9jDjrSnrOn2NOfaqYldsFtrF/m/qK7joYcwC7CLfbWovNL6n5cprprc6X4q4wdae1FR2n/fU4FBwtjxlRtrrAs/ictMUqMy4a6LvDE4v1jqXcl66UCrKXVLaaXhR23AwfnBlxDpBp/+6kp17mPMBmSiDZcfCOx56Nv/MDTuxyMtKHsfU/3YXJCtkBjgtN1TXCmZ+s0DsO/X7N0RqML4pP/ME8zikFHMYY5s5gWe/GvIkP2QGeEd/ZC5hnqReT0nzvib3ZDWRZpnjpX3bVK639ntnf179b3ihNlBOKz51MlJoxJDR/8jysKxvjhU7o586sXv4yLZTU9ZKiznld5WwELncQb3vVTrVUci9+DNP/eHU8zddv7jidc9GvSpkXiN2CsG9FZQ6JguPX5A8J0T6nbUWB7qXeY05lPlrqyr1TCysz8TCoDtSr+V9EyRTYVjzg3BRNEGX1B/UyG5Z+RQ1L2U8+cgCh5VLqLhgyyURALVKxVcWRqSF60IU3DjaztzFusxai9UWRASsHXMpifm2pH5prWAsUP8GPWdABFpH1K11iDTYfaayQ3E5JsyYYvxgFdY0PwHyf1GJOR+lCKwFeUcKZOkRmVvMx32/3iFmosuv+1kRLF1iW6QhL0ambsK4goW3uyZ5KFytZ0P/8GGTPlgy7h2KFAxp8YAsJ2793PwH2s62j33sHV1/+qJk+S82NQ597y+UfkNy/4LmmyMa+1a2rKvUjbKNrcuBec2+pzVnhawoN5r09GP6Ln2c/saYscoYjXs0lzJ/0neQIb/zDsPaRuJ9DIWClzuY9+hvlAWZQUzzPlV7PZIV64Ky70uP6P9/1jinMwrmYqLqmcmO8JFEW8SZPtqdKSx3tivuQ0oqHSOK16CVWmF0IvURxWOoltfi+hPNyXXSks5BPAS1sndG4aebCQvmv0FIOBEJcrkW0r6hLBP0uk2sjCBUEOwVuWuakPslr7QmC71K86vhJZsWghCFgkkl3ovaMbYWCRBkegqRWKK2uDrXllI5MwqondezyrGUIuLEa/tVV/oRVsf0LfopfZI5elXlHBaZ0ZbOFnMiJZhbu+QmqqjyxuRCKjuwa+5oaSWpikd8/a7o4uYu1Swu4mHb1NH+sV7FxIinK4OuV9/B80TChNmhtcjo9VPmzOHh3bVy4t3VulN//NM3flbymlPg7l7lzfyksuC+KpTBV1kuqpzrUMJqUgSz74XEr3iJ6cVlxkDr55YEWhJoSaAlgdeoBFqExWu04VrFbkmgJYHvLQmsu3yyYDVzq3VLBPBriQw26YAVAC/sSNiAYs3ARpdzAOc2ODSbGhKbWM4DtgMIcB/gH98twAlohGI4aNJLQM9NlhfWJZP1c67t/pJnIu2BPH0DUAPWsIlpbF7Wy2stLXgOoA7PZoPB86iTdfFEWSkbmxzyZ4PB5po6WVKhmWiwm45msN9qjPMM7rfuRSyho1MNeVorAfs/n/ZAngAnyO2nlQCsrRYjYBp5IkdkastggXRLCthPm6clGni21c6/WF243pqqWxDHAnj8Zp9jXR/ZvtFs9s/9lizhHr5bcN/+ZvOx5eM87WB3usjfloNr6IdsogHu/7MS7cz/AB7jJrG9YgpHFIN4h60b8icP68bLPueSnxdx+WTra8vPuKCe1J1+YckFZMtvlMcGs+R/Nvr8RtsBgCFHxhXXWUIFtwfIgvrwG32UcvMcLGzGlL6tRD+lP3GdrSNgEWUAFLSus+i/lMEZTLhO2nNiBT8EjKK8AH48tyFngcALdxa+eeoDzh+l+zpnbpqPZ7adS/aklqOZDWhDul6WT4TF08eK5ePb3ZPVfNi2tRCk9ytQ8w5VbodaCeDBAq/NbabTlz6aY23ct3ze7ZiAv/Hx8t4PyxOKil4ri6RI4HaHWARoKwOg47bm8+23mXtXHzXDNbmqCTdoMAMQvu9G9+naB6OffOxj1Q9/wzfeoeZSfLH/HZM/ce5PRgm+7enepuOX9R2QEudLnybgcfw9WYJEW3dE51mcjQdgC9ZP0x/d8ZG6OW9RYue8N+k7oNw7CIYL6fIWff7e1D/akIPgmd4jhZvrUbdS+fryvRIpccC/e6wH2ibPWN1NJ8tOX3/F6W5fcm/MLVR6+uqOv02oUZcbiZalkB2TO6iS7weZVCLmu34oH1xhOuG5kZVakM37TrziuF1SN/dioZl0A9Om2CDPyP3WUcXSeO/zhRtXFKT6rcgY8Hq7yqyg2zsExO8U+E47M+fga/+K2/llO8Elfly3GLAWR9OjpbPdt6w8tvrGpUdK59JDg/NtXYM93vRtvaXZ3ni0dGelc96tKkA2oJriWciyomq6l1fNtvGpaM+8XIgtraWJudB00G6fVmJsM06ZbxmHAMmsIxeYDYGiLyET/sPfbZDbgKf/Tv30E1gkFIK2RmwSET3R+erAbo2PsspzSj2bcQcgx7hk7DOOAV0fXH+WXWtfiag2dBX9w5rLQR0gKwCVJyFvqmHitlOl3W5X29x116efONgZnf8xgdZqXzkT85YSgbwPQbhwCHg/mau3/5Hn+scrkdhzU8M951aymZqCbVuLvLfpMlwMvU/pPZcpOMTGLs03b921cuLRvfPHHps13cn2oZn+iixTpitbzJnKdvqZyrH4PskMAmlGpEWgWAusL4w76kXbtGu0R6viH/JOJL2m6MIJN5iWKUWiUq15sjCShUnoyUKhHtTrRd0ceJ4br/uhApmE6k+O4P+6WyjV2oNAdjjyIqM8rfUnbY4GNO3DusGc2tAkV2rEGFGyBD/vPcwVKZFTblT9TSTZoIi9QcV3Ecm6hsWUlSf5soZ/eT0P3EHxnGWNoxqEyemplWTUi3SKsBBJEWxTuUcVa6O/WK5mZBS05EUEvDpOwjHB4oDjF34gkp8s1NyT405iayl0t1cd91GBrmsieq8V+Rk/lP3i51WGH9EzWHcuHFh9rPnZQ5OV7TMa8z2aK7M6Z99F6P+sDd9Zl7VVJLlY8/IbxCXWEbxL0b+t1VByT/7FM4+ft6rgGFOiL0IE0RdYwyGSreWhzX/zOwvnWeP+SOlPlWgXCLnC69QFVHM7MC6Q90ZLJ0kw0103HYOyggrjK8XVTCq/nJKzJvGBUXVD/S6QfgSiIdNVjBVXEz0iK5xkW7mowNIPJqKVxrvlJtdQp3W9AHxFTspUkl408BX3ol2ulRoxM4KqrP0qkVkvHiyV87Froyl5Y/MjsvSwzf+S7mMtgq17TMYR70aHRZoMtffnUl0jKxN61hlZNBwTedDZ3pv3vEQtJxdP/erCkGqMTx5AP2QM8521aZsS783zum5ecwnnurT+rqn+DSufkf1TqdJa4nfPHZGIAoc5DKuqiK5dlHXINSIfrCVjSmTFWhi4Gd0bSWVLjgiPbslpQLFAOiXLQVmssCai1HR+vxEaMS1J5opluYNSsPOwuY//mc7zbtGwkGkF3X5Jv2idaEmgJYGWBL4vJdAiLL4vm7VVqZYEWhL4a5KABaGtdQIbSDYVgDrWtRIbWvyKs5G37hEATNmEcI55Ga0pNj5WMxWQBs1u63YADVM09AAhrGY+9zdcjShZ4uJiYrCbWq45f29Uiq7aIhk3TTkABngOGwXKzOYDEJh82bzwPxsk7uU7mwvqwcYHUBcf1mxCkAWbHzaElA0QtxmEp2xWXracbCIt0EVZ+M69nAc0tqAVGmHkS54W6LfkAUAYAAnPBnxGJgQy5Vmcp6wQKvZ/wALq0tiMrRekmbTgFP9by5ZmS4lmYPpidbGABQCD3X1yP8+xz2u4IVmvCzKmDwCKn1EaaypPs1UH19E+zSQKZWxe08nfkleWSEOmWJeQL0DchBIACBY2SRPkBUp5tLndyNr7rghctcSYiAsrCytjS1QgLzsO6Lu0IcAg9eUZlM+SCGj/4TqFPsWGFhkCUtGelnwhP8YXhAR9ErSbcYEmLkATZAxgJ3JAnjyPvoDc6E+MM/ov/Ym+QpkswVjd1ebWU4osW/AbwJK19qEPjQs8nL2mdvSbP+H/cWb34PPX5lLxm1dEVCxGO6K+E3EgAaJC+SpuNEzXSuM7lqZ/dzXSmXvWvf6mlaATi43mg7FOXdHqfjmQa9NtG/6lrVLS1+yQhnQjOquCStcEkkchKQ5kHosAuqKxbI/Pd9xmDpROmhtK46atXmxYW9gj5lQ/8BPRTy1+2f/B8kQd0X73eKrjpraHuu/60g/OffWH2uReapO/9w/qStoMQPvJ9/+XTxQ/e16mtMXGjM5ryn9eiTZv1pikLvRP2uqQfbKAbaOA1ebNnV8w9y+/c0OZFDOgV441AGKsSyQbZJtxyxzRoXjBcpERDCvsuVcxHV2hE09mvNzwmuno92JZNxOPBxU/TOSLlaxAWhPKT0yh5HcpYnoiiEXF20Ty5XKYifp+2OF6JuP6T5bq0cnV0GkTaVKRpvsLfhjLLPl95xS8950DsbN9KWndC+yhXD+nRN9Eo/d/iXbo6vkgveHJ9I6llWg2PVw6N6C4pv4TYweWhhem2jvmlt+31pZxH7r7gASUN1Gp0UdlWSHrC5Ms4QpqzijmhOmZXzGxagOIf0AJ0Jhxwxz6NSXalvFDG3LuAmn+ctrbApqrAtTpIw33P8RjwAIIYooYIOrHNQHCgHD0A8aEBa1pT+Zw5Agw3CDrN3SGV/4P+VAXHK9BlJH3fQLUZ+Uaa1QxSt6ajBS3yRKgb1fquTcSmPyUXLwt1noNlg4EvyaehCwwnteYe2QoduYLynBKAeEZdNWhcwvkb+PmUAfmIMD3P1divfolJYD8Sx7xoHrb3xr/3dteWNuTn2jryc13ij4RaTKn2DhYJXQ0pql6Q5nh2fxB5l/mNMBu3iGYP0VImJzcIVWrIh68ejDvmlpH4Lgxoacxzd2iaR0Rn6EnMLVXU4K0qE0ZD/tYWOheR+EvyrK5CKt+3Q3LfvQLD/BqcuFgLaNOgOM8kz7PvMvY5zwHbcg4nRTBs/Wa1OHj7d7ygMiXa3pjM4r1M9EgKyRrO7fYdxBrjcVcfiEGzKoizFSqfqpUqfWKROkR2TiitEXMSltYF+DpiHeOuAMiLtq9iDcnZ1dTKSes3+CVZnKBd3xR3KNcQ40qXSPyYZssLZz7l9/1R+/o/tR/VH+EHcX6oeGiij6qz4NbEie/JXKtUAmTmfPhyRqyBQCnjflOn325cc5vjBks/uhr1KdN83U1FlT7RAgPFQXxxurVhEhhLGxYD1l7fnBdhhf7YP1gnrXHhL4A8v4PJWSPxWm5RVY0xGPfXTeS6Gq9uq8YNApNUc5Fvu1GEzcqxkMGgiEo6nVDc5UsF4zcKtU6h1ei7QNuWm6PiD9BHIi64jjk5sd7HhcZcb2ctLKmY1WRTLSXVjyvnhVpkE61ldcU0LoaS3mxSj5WUkDr5XI+cUptPam4El3RpD9dK0ZXRFhcqq3tex7vw/Zgsn9O/vqOqyxbREzUFEi70taXe0TEyr50d2FMxIqCh4fMRdxPH+V+S2hyjvXWugNlbuY9kz7XS9302VBUkjun1PaDZ+5fmuz8hmJXJNX/v67zuMN6plKMZWZO9Ja33XTmmO7p0rVZGVg4kocjCwzFBgknVY7tIjashRDKCswVlEvmK44sPMxK4NfyMnVMb5rY2TfdqcTc/1dipdgkz9bXlgRaEmhJoCWB7xEJtAiL75GGaBWjJYGWBF67Eli3rgAcsFrwgKuAZIDnvOSzeWVDwYaWDQAv6xbwse6feGEHCGLTwHeAGoBMXs45ADLY4HKe72woRpRsQFXyJTW7h7oYkAOgYAmV864Haiuhqcxoe/F2yg+gMqbEdxKAA8ADZUKrlXqRhyUoAHXY5LChsQAJm2ZkYIH/ZksE+5068XvzNVZDE4CD/Kgfz7MWKNzLJgr0DDCLNQzgnk/yof6ApWzcKSMapeRFnW5WamiLrZeTvKzmL/Uk32YN0GbZ2e/2+ciPvJCfddd1sboAflE+wClrKaKvF8gLmy91RM6ACpQJ+QHk4keb9gUwQTZW9uRhrRLIo5kIor9RD85vJkloJ/qdJY+QFWVU3d01k9wzZARer/9uNWep38XcWnDdS46msUAZuJf6n48y/d2ApHyn39CPaWM29siIZ/Id0guAiz7OwTXUl7EBsEN+jCUO8ni3EuML8gE5sxmnr0JGQXYgHza4jEf73sPzf0iJzTYEGwd9AwBjIe+HM1+f8zsEcg3L1/st/nktb/pXm8C8eLpeKN9cebKn15vZsZJI9Nejjhsv1vLpaCkoR2OpjF/yU5XKQiGeWKq77tzkQM9iopJ7qpBD4df58fXn2Q/GEuWhbFdEWDRbV+geO/cAQKB52+hrsrKQUwv/lIC1qVSksCti/L5NwWvN4eQOqTkuK6JDYNJh+QL5AAmx3Z34xXd5Xzz9n6t/e0Nxq24s+wcjHzxxx+I3xzNBfjsBhDcdtAft8xu3LT/61c8O/gjtMrH5Iv2P5QztDOJJ/+dABswdjNdDm++RGx4A4tPr9zX//LP6BwB9QbKZLLU3wHrGC2lA5M028Wi7RVYM+KFQm0iHgkvHx1wv2larOJ3CNfOezC/yxWqPhBlvy8RX5PdeOL1U/h23Q1YUq4pEHIt7vumuVOZkpzIrdzK5iGvSilIsbzpOhywsphUguHpN6uk2xYX4CBrvgPE6mL/ov2hI00b0xVcLZL8gA1m0cDBHMZ/RJxh/e3cUTjJ+DigBXN9177GZLb5icpwe6zdPv3F7wxXT5uPNX/t2g6RI50ufjNYC2gRwHbcyjD/yYWzSZjyP+ZU5on6VLmZ4sBae8B+ISPstETxyo1Q2q4rFqjgGtz+48vb/NlsdeWy6OjopMug2XcvcxVw4oYR1BuP5giXHSypxlSfW4zAw/si3Ae4rvUn9Zo+IiC6Vsb5U6409nbvtjSt+V4NkmapulUVIW8MNFPE+FN/g7M7kC19R8PKH9fu8ZItsCP4e/u3z7WPbnU/GPK6xmHQZB4DXuB1inmbu+tDmKuCKbbg0Zcar2zPFxU5TaGtT+5XMqsqjgO5G/Y6A3r+ktvuHiutCPRhL1IP5lXWcc7t8x90vMP9zfUF5RUzENUFEdETopKTR3K6eU9Uc5Ym4UGFlHqb+LfdoVTmw6ZSLpVAmSBJ6XfFdAuJZOIO9be6v/uET9V89XzfmWupMnU6t18VaXDAOWHsYnF3K/TbldIvi7uyQ7HolrxEIM8iKdrl/E3hvqw8hDUkBYcGa3ohZYX9cK1RUCpMulvyeIKyP1vz6oAZkrwaAG/EiAkHD7qjnVkVmpMqVIBkEQdSTR/4dkerquUh1Wu5pDso53l3qyLKmkrc+42x9MnfnrXtTzyzuSD2PyzIC0sutX5IYK0YElJGrr3e/ULhB7yAhYxmCy1qVMi54N3jJ+N7s3k/zFO1yQm2qmC6OL49Cic7achoXaV/veXP2pyf/oBKvV6gvayhA7cuSWfqd94bfUeI9krwhKiAYreJGeJXj04r4+/WTccaaf+GoyhFaQW9c4qP7e7bVR+pBQTEY6gOyijBr8xlZFLimc2SllsoWo7JakJe8MCmCoCKLCFcg/E4RFklZE9wiSwcNr0gj/IKuOZDuKE96yZoH29U2kFuUFYKvOBCDsjTwTejHoqnqiL4XkrHyUr2miaYeYQ292mO/yJXnRL89KVdMy/FUNdxx68RWPb9TREFWn7xbNYhCJeYD1kbmdhs7xz6PgccY5RPLT+ZYSzIyhjPRZG1v77bFcbl4mpKVBetL471Kddh6+qmRes+Wpc/LLdVJ1feNQc3rliVFFldz3VuXQpEXx2XstEXzDWWw+xz77C4tmitePBF6sbjyq0qGF4Y61rS0GWPufwnpf7UN0Lq+JYGWBFoSaEng1ZdAi7B49WXayrElgZYEXp8S4IUekJZ5FdCTzQBgTgPkVAKsAoRAK5SXfl7Wuc5q/1uQnw2UtaBgg4EGvLW6YFPMvWga8WlBKZ5l3eDYeAPcczGgmesoK3lRLtesfNszXW/xTFDiejYqgAoA3+QLODyx/h2AEZ/kXMcmh+db8JtPC5Lb3+ymwlou6JJLWllwL2AYdQY0sppvnGfHQjnYOAGSUXY0UnkmpIHVBKNcfAeo435kD3hCfiSu5xrKY8kJ6mkBPn6zLjuagSVrrWDLj4x5hr2W8xzWsoB7KSvgJPnTps2kh7Ua4R7KRZlpT4Ad6mYJGYB0+gxy5Drag2upM2W2Vi58t6SFtTixVi0WwORZyIL+1iwL+knW+GuysFF16jnKSVnID0DNkg7c/7LHumWF7fOWtKM8to9QbvoXMqGe9BNkxKaY592yXl/OUX4AKtrJurey/9MXaIOx9TzIlzoBbAHWsAnmmbQHdbDaqYCQgPnkR8I9BmWhHOddEqz3u5VaGPyPGX+71JHfoILdrvOQjPaIj1YnpzqdhVGnrTq0Gk/1eZEg2mlytV0zZxfzPSkzFeuO5OKuFzP+dCkSezDu1b42ntszV6knKCfAerMbmLfqf4gTgARk/0rAbOoFSQBhcQGEEWhSX/F7pmaqw8+Mxk9h/bAZnDBfb7uhelf+2erOylQGyxCAQqDKtER8j3f/1v9S/QVwFgtaIIOiAm8X7u9586+8d+rTf1PXA7LaA/IBcudWafPf8I7ZL5390+Efn/5Ox40NDeVNB32PPlmROyhLOAKq0oa4mrAHVkEZlak/6tQeURwLQFcA3uaDMdBwlfEv4h/lQbQvlg30k62690OqlfqJ0+ab1IlyvdPJm+7hfD2VKNUEk1erQ9IcD32Bmgq47UQLUvAX8hu6biSQP49oPUgNGH9WHrvzS14wWw5q448FqZFi3VH8C4HbjlmSBv7xA5lHfQHvB0RWfEdkxY3r1ieW/H2byvJvlDpkXbBytW6h1gmJzTK0/1Nn5Emfp+6MCebIe5ToG3+HC4NIxOQzCTM91G2O7d1i5NH8JfltnZgJsisFo7gV31LggkckBuRtLSn43uwa0BK1RmDoyx7NAeTXL6RPMQ88JDk9Igug23Ff1hXOCxxOmDuzX/kRBS9/8r6lH62IIHhuvU4QkZAVjJUrIvdevlQbf10nLeiTzBWQJDuxkJC7MU2OYUmWE0s1xanFskKkilwXrTbcF3lOVcCyc0ZWFYXO6MLzMaf8XLGeyf2TG//4cmQvMuB5kNXMR1iH0V7Me3y/S2lMiXkUwC6a9gsmpbjtE5VdZmGqyyx1dMjV25q0/2ONeBauG/y4rGJ++8WMIk44wR6do98BdjM+IBHkzcz8/+y9B5xkWX3fe0Pl6urcPT0zPXlnc2KXZQkL7AoQAiwZkLASSAJbz5bTsyzLFrZsWVjv6Tm8JxsHOWFZAoGQLYQRIMIiNrMLm3d2Zif3hJ6Zns5dXfkG/77V9e+trumZ6Vl40u6q7mfOdNWte88953/CPef3+4eBRTfRsxx5RzR+T7p4dHHlMi2Od0eNOFJsilCBtRf1vSrfUAuKUp8ScujLcqGhjnZelhdy1+Ik6o3Qm54vdc5XdCrWKLyDAdwBGHkf0B95vkZYmJLTm0IhsdgrOY7IJdjwjswRtyFCgJg7HcQq7sYeUmLtZFY8qw2n4BsqkpsJomhIbqBGcLPjud6wLClGRFTIBExmbopiIWLGE2mxSUBpWgG58xrvQpar+5Zq7lm5hdq15PhPVly/oMq8Vv1v/IHFH3jBdxvPjKVP30IQ5aaCkaQAACAASURBVHlZ0FRkQbOkoPRyDZaRtYViqPu8i7Dmg3iiHVEwQM6XncPpa3t/97mFfFg6PJXetEdk7A3ZsOI2vGTjRHbHlj8efdczml+3iNCAWL8cWYE8UG7BTRtrBsaGWT2x1oSs6B4vSoBxx7uB9z+EDjG8VgJu6wxTfmGk4pYXGs/L4iGdztUSiXTQ1ztaDBR3Qd4Do0Aul0KRFMfDwJueO61ljVxFKa7DqJKMA+JljZnmulQWGdOZvkpVsSNO6ZrpOPC1pop7FftiXu+Niu7P+4F/Y6OS3LQ8mz8tS4TXiAR5KW0loyl3q8gS1ujzIijyIi9Q/mBtxZ6C9wLrC/oocwn9gj7LOKXPsL5ifKLEwjnWUfxlLmRdznzINd/Uu21UwbjnJvePTckShD3Kyho0dkYUf2Pw2a9ed+SOH376eVlT9PnJYDydc7aJpOktTvdkROqc0nhizcec0G4R1FJ6cjNSJFiUa6iDXrJyjcwe22XBfbTXZcfXSxFg956uBLoS6EqgK4GXnwS6hMXLr026JepKoCuBV6YETMvZXDOx+Gaxb9r7bCIA4gB+2CSweYcA4Hczy2YzDtjIdxbyaC6xqOd6QCJADDauAOXkz4aI84BTLOC5jvvZiJm243oaqIAogMJck3CkZOjgBaIxpQ2MYom+GNSazRx5G8nBZoX6oaVlFiH62ATJeLaRJgbcUw+zvOA6js6dWDsxgGx4JtqZyArgg2Q7Fj6j6ctGik0X8jOgztyGIBtAdspqwDQgLZsu8ichc+RCOfm7Yo6+8hwS562cZhFidSF/5E4Z0d4nLzvaN1G8X/nNrD/a8+G8XUt9TROWdgOMu0cJoAqQbqcSMmwnhCBtIDfMgqL9uUZsWL9qJ42s7yEXAD+TX8XJXtXvLD0mrzn93If8kAN1Rc4bPYxAW7HcWemvlJ/PBgIC8ND3KBebYMA52oAAy4yJE0qAP2hSo1VK/wbMAxRn880mGxCM9jVXUffps/U9yswGmnwYc1yDfGkzygJxCIBGPRkrjDPICMAeyiHQzMnO1uPt5TAe0mdIADbzlAO57xyKZifeHX/pya19x/r9vsaOhUy/fKrFjnzUB25PPLCrfi4aipdOnU/3T1T99BOR635yJtE3+a0zNGlT7g8oASQjL9qE59Oe1OGlHvRx5gvquHqIJNgji4T/ef/8e77wo5v+0x/LrdIXOh9Ql0uUbxRekyp76UdurE68kSDhAO3C75skw5g75ZyNx9r7eW450fPaf3nV3/uT90x96WO9wRJgOG5LOCAr7PjlciKXvWlpX12EBWRJ5/G/dOKUtKuDqfrW5KbUJGOQ9qH/MP7toI0Yb7+tjv6khk5R5btFZaO+tDGy44j63cX6uxNfoQ9AaOBSY0rXvVd/P2AGXarXYMoPn01ExbIsJwoiKLyU69fFUGS8yE1Ks9ytNYJ8b0+61Ot6YbkR1f1Q7nDiKCXyIlFJpPvmneQtarjnRwRiFyNnSb66n5Z7qDOKZdCQJn5DMSx+Vc8EPGTcGolIGenX9MeKAPw1pg0iMNYR0SVP2RxF27S/axgntAPzJGAnY0DBxl2nnEs71WzaKfbmi5PjI/S9Cw6RGg/tv2HnV2547thS71IZcAgSincTcwHzFYnjuwWNjKRGRvjYfwP9jjgQuC/LeaVNm1Jn3nlTz3dOPrZ498F6nGbMIzPmjssRAVcqy9XrBSSH0n6nrg9ovIxJ43+rtP9zCqQtrX1ZIvnFWGC1i6u10dSZZiD4apR5oRrlH9Bn5CULi+oZpTVI2yUA4ybBLUKK+cesIZgbPqPEXEj/Zgw0CTARgc5sUorIyl3ay045UsBtlQGrDwLSQ/r4Ded9uw6fvS81ULum4uboB7wXzFryAT2wLCuL03rIuSaUH8TlhO/L31Ez0HZaQee3avTL3YtTkIM/VySGK+OKms4VU8nEZDbrnS1XnWnupR/88gfvIFaNyZA2otw8F/CT+R7SmDo9qES/6xHJ0ieSorYrc7Ahki+L3YacxzTzaHMzx1zP/M/8zFhvWqvYgz774LGE4laIU3OrCq5d14d00k/01oKGp/JGVREsIkZkARP3KW54KG99cmcV1QTsBlEY7sjKN/91rjs5FSdziunBOGkpTLh9J6u7Gw8tvvPYlvSJJZFSW+X2TXJeIIYFljQ9b+7/ivfw4jvOFYO+bZIZY5A1xgUuyjotK9TOjFtkkZ5/6C1D+wvXbf7H1/6zvrnUUP7t018/nwmrd/UGxTfIek1tvSHg+neVF4A044jn4/rJLDttLWgi6/59UQJ0WOZm3u9Na4iGLCwijatEOp7vHQkKyczSIVkNaM3iDsgNVJwfqKRlsVNU0OmiyIBsFLqHTz239ZgCbe/p21Q8U5rP7pQ1gSsSwqxKHRETcWUpWwkzfkEulDTKwuXCSCmb7qnreck+ERxZeoTuGYmW0yOKI7OofNe6qtpYq03LEVR15sTg1Yqh8diO207NiFyBTOPgnUifY41lbp9YS5MgAXjf0ldQDmD9xJhlTcFcD4nRHLOIqSWvOcWkeO1Vbzi+7+iju06o/ssag1gE36krliWf8Rfu2/vYTe88MCfy5m5NbAcrxUy8cLa3UK+kWO9AaLKX4V1vR3M9C9+ovBKu51/DlCQDlvbA26wpUXphjvlu3z9tj+5+7EqgK4GuBLoSeLlKoEtYvFxbpluurgS6EnglScA2oAbcA3YAPKDhy+KfzTZABht4NkdozrORYLEOAAvwhuYoi3AALeZmwGQW5ACmpnFvYBG7egBZ7mfTRd62QWJBbxr5pnnfvrC3HbAB9tqyDUqtOp12vBybmnbLDPIHXDPXRmjsUVaA9B9Qor62EWJDc6kNBL/xbBLPXiFLVrTaOdhsc55zbLYFTDaBNjaU1IlE/TlnsmzdukoamIYjwBabK9PApS3arSTIH9KFTSGbNAAhKxvl4npTPe5EDDhPvgCiRmK0g7lWJiMoeC5tbKSSkQz8DhjTdKWiZJYTuG5hA0mZzNWWWU8gH7PYoK7Ipj0/yo6cTMaUxcgjSAjuIS+AerOiQFZjjrzdNMkKqeVZBfTXyK7LoiYt6wpkYy6yqE/T9UfrnBEE/OU8RBx9m/EBSEQ/oky0C7+xmeUvhAbuQJA5edP2aCJzLeAMvyNHfjPXUFQBwJY8aV/kyBiiLAYIsiFHmx8ihHoCyjY14aUZuSA3UH2vG0z0nZqs3ykgg7yaZNdQMPv0m8KHl6/zXrg7k50tzqYLxUxQL5aTmXzkJ2p+FNVn/d7lRsJ/MvK9BwU4PV5zk2cFskWZz/2WuV+AtPgdpd1KWLwwH3DOxshqGwACdgJeVK7jIF+LI9MZJP2TCl78+YVg4GjWKzN+/5ES89Lf6MzkYGZb7draqWN6+G4aPCWRiwBw7kx82/l844c6L7/2ZHa790zfLU+8efbBn2/JGoJg9YDsUF6/MFo7v79FLqz9eaXNhvr8OV+a6vRb+g+Ayo8r3dbxQObQ3xQRMHp9/qkJAYWfkML3r+ickRVTSadx/Rb3TP54tOvQrf6zt0pzHOLvRtVFLGyTgpFLF3m98cKbi87WfbPhzrPFKDfQcP2cov4uCpetSFc7h9ebtO9mpD0+Vm9EQb0SyOGX25NMJ2tzDScxIzCpFHlnhN4mM55zejjlPBm47rEni3FdwKYw0YD+CsAM+ch4bj8+pi8QPIxL+txLAV1srqLd+czcD0nBuKJ/407rZ1vfm8+Wy5mmdcVSX94RUeE8ccc165IV/fPFByrZ1H3F3txXlXFRALARFUZ8vpTyNstghEyHpQX9ljH/TRMSLUUQZpKA+B8RkfXUtvSxZxSrYemL98hQ5k/niBTk/biIifvVP+++Nv/M8kx9bFPoJIK8V5xdCgeG67JomG2MOgoSfXxL+uRCJcw/oM+HFHT9vOq6nqLARkreJC9aCdljZQGYOKHE/PULyajh3Lr4jDMUzzpf336PJsTvg9xpulLCNRSuqtxafG1jIde42X+u5+nCrSUh9TKK8GZFdgA+0vcWFHx7+kknX7w6Kgm7j2vJpFv0fX9OhN6IeIiU+kyfqIxedZ2MOLxZvRqm5Y5eZYrlssZdkmXDsn6/0J/YyjuG9wpjGU1u6gFZwmfe3zkRvOeHkucHRVoMqp1zM4oFPJyYapItxKppHczzEKxYVzTJqk6rpKH+nKPxmgiDMFuu+Dm5rNK7JB7RnC1jqbjm1MO0iDq8W/VIAFW94CqaCxSGJhJR6WRFYjS2OTX3Fi9xuh55Fbl9O6xYFsz3p9X26VPVXX1y+bU0nDy/JJKidzBxXlYsCdzS9WxKnPkHI8mzny2H+f26FhKcd9NF272dqGi15Q65gBrcUzrWK9d56QOF67beOf/tnz7Yc7VzIrfDOZ8ecXaXjjk3LT1nBA6up9rnE96B2E2QmAMQHHMP7wDkbf3I5Nn9u1YCvO+ZowHpm5r+kBVyceTMnfbL1WI4K7dHN6vv3KL+nqgWMydELqSyvdWaP1yKBdLvk3ujgcHx+feJAHNlbVGArBAwr5gWtixr5jdans9WtNqMRX7gBspPpIKC4jtobMl0Kadg94G3JGqtl7dB0zXbyruhnfy/VNvR7hAP8lmlqV5uqnqGl39Klhb36fsJdR7W6livMreYNTb9g7Uk51hHoRDAugArClsfs+biPUF5GIuMZ+6hXA+KeBnYdNXMtuWZnvrZQ6N7VH/mKdZcJ4nrcv7Y8K5vfea1D++87dR3ZFlRnDoyMir53CQyhnXIW1syb5/PKUtFigGHg1qpX1FzhpV0ypbSzbUcX16qFeqlZNj9rSuBrgS6EuhK4GUqgS5h8TJtmG6xuhLoSuDlJwGBsnKvuha7bfnst8IaYAsQxyYCEA5iAlCVlTdzLkAsGyV+M9IAIBkNOQgNQCfcoXDOyAJIDvIG2EXbkIM8uQbigk0EADoLeXP1xAZmPXCJzYhZLbCrqkq7PucExYoUKykjIHETuG3lz7MAk9AIZyPM/dSP5xg4baA417aDrgasdZIk5G1aunxmY/SoEuAjZaC+gDNcYy6ckAX1Z/PEJsosFwC7zCUUzyc/wGk2ZmyeIFuoL/kADKPZZRYjXMezjCjhftPc4v723VJ7XSgDmzxrU7uO+62u7bI3LTKTk/nyNpdbRh6wSYVosToCPAKEsJG08pCHETHUDZmtR0ixuVvV8mvVi3qzUaUPcg95IeOiE9erjicxVY/RL7kX+Zplx0Y0/8kL2XNtU3tUyTT5aCM2wmx0AcysP1Mn+pBpp0KGQSDQXsgEIoKDMUGZaC+uoR823R4oIRs25ORl7tB4LmSEuaMiL8ahaQ2amyvT0Ac0hShsuhqoR3HxeCnqVRRJ4XFOTgBqSSp//JQbdc97N7nPystTY3ct59+INrjAN18xK6KR6sLyOX9AVhWp5wei4n+Vq4QjJS/b+Lnbvmia1siT8jKWXqNE21Emxhz90iw/rgSUpb8hP/oMlgSdmploafvn6tvoM4whiBL6GPV9p9LqMecX7jmZHP3G9eEJxpnAPAXwcCedt/oPOstxj3Nv8H3Na3WesTQp1yUjv3ztry3e//BbyffvKD2tZERfE2Trkfua8eppNCo7D8bPOclvXgREJKsEAKO7lf6fVn06r6ev466qnPeWk5L5XIeQNkkQP/uh1Kc/3usu7RA4+xZd26wfxIlpbFfjwslKVBiXL/qRKDl6znd6jwVhZqsaWq7vo2UhmwNyAxVVxGwobolceyRc+YMS0iS0U16yZHsyL/fk03k3OtCXip+vu86+XXnvZMl16o+8oz/6hJ4nQJ7+Bgj2D5S+0lERQJ9fUvp3SowFmwfXEdFFT9HezG20tZHk9B0+/10lwKA1R6Ag4jMjfc7x3ZudF67nVXHhkao3XhBbt29keuGJ656fOBH4fnPMbTRIr8i19ea+1QdBvD11asl9zbbemL/8oM+R5MVzGAP/Qemvc749kHvKrb3tuvzTv/3f3vTRKxkXVyLPC67FXc9ffeZ9kfrJtCwYJuQW6mSc23dXPUrNVaL8rMiJYawa1MeW5C7qyby//M2Cv/is+vHSd0FWdJaD+jI38d5iTqPPPKRn3jbYmPvHA3PzzomBceepioySNOqWvT6nINdQVcVaODE8/s7kRHDNzcVnS0O12an7h97q1d3UZgVwPqsYNICPzTgdIzI2EPFQSSb9WO6eKmoUWR+IC/FieZOKd8l1kmI/OCIyNNFFMhkJolpdBlGNRlQUoVeWy6X11hi0rc3rvAd4HusVAZpyU+MGM3f2fvOwHvAjGa+6TQHLexmjEC3EU2m1PXX/AyXievAeqK3nQg3Coliu58vlaKAnl+oTSyEe0c2kUomluBb4wm97ZVjkplLJUK6tej1ZUyXCaF7n51XIuvDQRjqKEte4lfl9TkZxOpx+LQaaFloiJo5Vop7ZoC6f+5K/RHD94cpNTjHo1YIh4Sg2kKM4F77IintPVK9ivNfoN+2N2CQp/sqqUgHjk3UNwC6T6duRjUiL53/61O+86+m+W1/fUPCEJSn0i2ASc1px9heud3aVjzuFoMj7jgSBxVw50ZIN8wtgM+865hKzQHrJxGJ7+V/Fn+lfrJE52tdJTUuL5RkvrGiK0uceWQjkPd8pi6g4JoJhrywsBvV3XoFdNiczwXVygZRaONtXrSxlckvnFc8meJGsIHPAe4H5i3KFlBDJQZDqipfIbE+mFOpePdRPhJXaclpkRfN5HLxDUebY6GF7A13vOtVi+oDy65d7qR2ZQu1+ERf0NfoHawDeu4wn+gyfedebIhLrMuZi1lXkyfqItQLX8c5nDHMNaw0+n5GbLHfHa05h2ZGaOznwlAicourXVDgRifOO0lzupufvvYb3HDWDrDQ3cZ/VZ9vvmEUu8wafxyQYOaZTpJxQIT5ejJHFnoO2uqwCzUYF172uK4GuBLoS6Erg5S+BLmHx8m+jbgm7EuhK4GUigU6ygmLpnNbT2mmsHEZY2NzKzoWEFjlWCYDyf0EJAI9r2MyjWc0GAYCVRT3XQESwyAfkBZxlYc/BYh+tbLTo2DiY6xPAKjYjLPbZWABG8Bsbjc7DtO9XgcUmLh3MhM7yU+ecnmv4nU0M5Tb3SahXm1sqCBI2DZTPANj2Z5gs+I087HmAbHw2QoC6cg2WFMiATbgB3WaqTp3YMFEOgF5kZpYIPJM8+J1kxIW5RWAThkw5jxx2KhlxxKYfwLgdAANUtjLa+fa68JnyQW4YMM91Vg+7l3LZwT3mYopzRnoA5tCuWFJQbyMPQBIBZvkO8A+xANjDJhLQnvvNxQz5sqltfwb3Nd0aKZlFBflwju/IDgAMeXA/coYce9CpntjthMtJp/hkJyho+a1W6hIfTB7InbajDyIX2qfdUobnc40B+XxmLADe27jgXvKjP7NxZrNKveh7jB/GBPIhIRvKSVsD7vE756kvY4U6s4mm/Uw7j+vxjQ7gQxkB2xmHfWerce3RuXDn+Vo8LsKiLxvX5grhYrniZTaPJ08N+PlGjyDzcjYRK8SFsGxHDq+FaIuoOJVww8/PZXrPzrq9E7KsKHWAbNQHUoRyYkFAne2gfNSt3cKp7eeLfkQmzAto3kJCdB6QRJChwS8d/a1IsSLQVKafGRlk47R538M9N9Q2B3Mf6w3Le0XSfATwcElxeI2s4BoBgsmEI4fucuEz2b/1awK0zwuYQ85Ybfyk0k4l5qK+sp9LPd3baWTQBKQ/o/Sp2wqPnLp74MsZgZe4BONe2mK9gz7Eb7MLwdCM5I62MXWgbzQP6eTvLDjFv3STv69fhhDXqozN89RhxdrDB9AbipzkGWEgS/LaMa8QFEPZpCen5Gn544/r5XqwUA8d+e1wMgnU6YOGm1BwbYUGaNRqDT/jepXxlH+k14ueTcqqIozD02OJRO3OTYkYNJlDbV4XCI886E//TekjHRV6s75/WQnwclUrewMxKqg//YOxxFjnO/2G/H5MCXda9q5YfSTWFRW5gZoe6XfOyLqiodZb79B1n18uZL8VJrzHt09MLe74Z5MX1RbvCPpOHzTy0chhZB38la1u+Je3NCOPu84KSeGKrDBSGwIjfqb469FS44hoIYJ7r4uz3iEXUeOSKe+5C8r0ElxprVv/9pN6VrNOclc2qjQvAqyp9p/3nMFeZ2GQgLpg+OpXX5ETmf8uEP65pOL1fg/JCisOAuHZ9CXeGTNeHD0ht0FnS4n8e894W78fS4+ZcJMTSau7ESebFgqLPYFTHRvduVgedCp+9oZriy/s198pER07pbX/VcVMWPjq6DurX/vRPdHXNM8qaHagINp14fmxyIlG0vWfUryHstzTKFd3liWOolxU9N+05sRzssAoKxBFvVoLLhZHhMHHXGMgfa9GoML6VGsDiZnsnuwLN56s7dkdxAmtY+IM8UCyshJpI6ru1b2McRLrmXXJqsVi1a3Vw7hcDTKJhJfNZ1PeUrnWr8ab9xPutIiVjAgXlm5VWV+kY8XckBVJoxkM2XeXFIC7LA9b8r8ThrfGpRNnnNRc4CYG9DNz6V7F/+j1Xf+cLGeOSK6jvhMMK5i5ylp2xtMTuAS76tbCo7Xp+lj146//9QvJipX3rmm1Q1Qwz71HCRdZO5XersDazvbKiWbkoFKiB384zqbalFOWpyAsLZ4vXP/Qaxaf/n1dhxyYI1kvfUPp60qsFxhr5Y0Si5ft/H8OLnjioU/Ft9/1QbOUZVzxPls9aiV36PS+7LneTc54tq9+TtYQIi2iQRkqLch6Yri6nB6W2yXIiHjxbG/i/NFh3Iw9rTgUb0Wn6UWMvZnlEVlm7ImjTFlKDAVdlynJUZniOzjJtMZpMSPXUqLg1059rA2Y79qJC9YNts5sd6W0Wm7yEDkyLrdQ5TD0ege2Lvap3LhnY15mDXW/EnMbawD2EOSP4gT9lDUTLwfeKRx85j7eKayrWDvxmfubVqva/oSyEDmpeBZ5xfTYcu7wyFnJ5WaRNle1gmqzfm23lG6+F5Ta14RrCQhF5FYMi8jVS5g3d9s7gTqz1mMdT126pFyrobp/uhLoSqArgVezBLqExau5dbt160qgK4E/TQmYNiSLbxblEAuAhQANaMax2Ee7/dNKbBDQCt+lBGjFRsFAH66zzRP5GCDN4hzrCjYtTykBuLN5ABQA+OZaA2lNYwyguyxCJYRYaQmDcwCczP8rBEHp2Yqz9ed6nL47duo7ICAAL9eY32vAfzZ1ZjlCvXg2GweOdpdHyME2VbYR4TvP5zrKafEieD5uIig3zyUhG4BmgHw2S2xSbONEfqaNZQAGZbS6sInhM+XjOuQ+0cqfOrDZYaOE7HgGQBBlMTJCH5sgMm3A7zzf6mJqc3xvB0+41+q3CsSRkY7270ZWcI78KSfAOsA8z2ITx0aRMptlCeXD4oA+wn1cY5YlVmbyarfWoZzch1zaAXH7jnwpL9fQhjwboDDjNJZyTnKE64zkMALCLBda1broH8pHG9NXAGkgmagffZTn0SaMC36nH3MeEAeCDCCS+83qCBlYXckDcoW60nbI4oQS/Y/rDHSnLc1CiELSX3ke2oQ827R9AYm5h/M8k77R1CqUVn14ZDncPFGKrlqqh6MysujNx6XojsYTZw4kr+4Zcs9Hhex02sk0Qj+MZoNkQl6Wg32x5y4u+vkDRT93vyDuRelOIofOgzYz9w2UBXcU+BuHNAJ4N9dk69z64qkOsNj6GCQc7lN+ruNm6s24Cprav9Ia12fk/ttK9Ct7dvO2qpt69x/1vv75u5efnd0UzJ/oiUs7+uQWKiP7gqo8w1jegZPYrdgW1272zm2b/tzCjPPlfur7+0q0C5rDELMjCijr9AU09cqheBfzxUQhP1CfLwYpP3lj/vFRAZWMddoOEK/zgOj9IyXAOvrmtFwEzeXccrQcFz4pwPij7Tc8G9101T3x/cNqE5mIvOitBndQElRacXYfmwt3PT/vXy3vToWoUQ9yDS/tZTPybC9v2dIyTwrkTLgJr66Q6Qm5xxfIFASZTHIpDhtBWpq2fto7v8mPTvYkvIlQZMWewcx6wAkPp28/pNRJWFDkf6j0hBLA46UOG+cG1jBnGGFMfwH87GzzNflFnteMW7EwUDg4P9ADEHsBKSTa/dNBwj8o0uKRWjq5cP0vXZysWKewRjZCPDKnMH/UfFEUX5iOj6sxzv/FkaaPf64z13+GRNVvKXw0fHLpV/eVwlOv1avqEUVpeGPHMwDHOIcFGnPHGnnjYup7QVp0uKqy9zjP/mFZNXyoWSadlWOxpostHf9BADvv5G8pMUdelOC5TBs3f75MUGQjo5dFbJVO5rb/znyy/5uHC3t/OPQSPz/mnBxKpqtNd0Vn6tubQcvPb97iXDdx1BkOzjvvO/v563NBaXgmNZJU3Jmn+oLF+/oai4EapEk4EINCpEVdMSmKGgg1WRzJCsE568VuPul7gTKO5TZK/+KykNWq57kNWViY8kGz/G2u6+T+boF2elgJVzRXSU6HZUHxvFxn3Sg3Wlc9s3znTQpMv30gOdsE/0UIiAtZFR9zPXMyIOk0BODF5FeuKsqQZF+uNc4m5c4q4XvS7I7FvRBcm5gbmm/lEkoFb65d5ByqIRzUF4mxRXUcUHs2Un5CBGjs3BSXgxNB4uCjiQFIgLuVdmt+0bwUZ2RNgbu3WZEVwzszhxyRWE1iSKTVrTm3+NqxVANgdqnl9sn6On0HpRPGnPV95kUsJ9cciuHsDDbmNVcuOvlg2ZlPDThP9t3mPN13y1NfH/n+e//2sY9/856Zb3IPZD/uQ1EgQcbIpgvcXqyDXPo8HQ5i+bFWG61e7bp+de7U2PVHvpXq08sqMbpnekDWFOlsX2VSVhFyB5XMzU32R4rJ4AXVZEUkwbRcHV2TzGluUMDssJ6QdcAqCdGjzwqI7eGqbOWIfKcqSwxZXTQtMDrIiuYVSp2WZy27tAAAIABJREFUrWssQS5eNbeAtUd0YnD/yM65cHjnLOsd1gDm3ok1CHsPI74Za2ZBwTjhXc7zITpYI5CY29l3GCHOeon1Wb+XiMoKRr4kYuQmpdHSXD49f6YvIeKioHrt1DWsyVgLIu/J1rOaLjZbeaypCuM2qJaToYx+Y1lYtB0T+vxtpS5ZcfHG7/7SlUBXAl0JvOok0CUsXnVN2q1QVwJdCfwZSMC0INnAs7gHSAKEZ0MAIMkGgPNoGrERAHwDxeMzGwG+Mx+zQWEj+qXW71QFZARgExCejTCbeTSvAFs5AEvYtJomH5pTfOeZ62n980wjFVa2T2FFfggerzvpsXknu8diCLAZBtxHCwvggE0yLmeoI2WGfOF3wGTT9jLrA/4a2MwzeB7AMhsUNu4G/vMb59g8UT82TeRrpAp/uZf8uZb7DLgxII/ncx9gNhsjyo98uIf7dyphtQIgDODFhosyGGhH/oAA1AUwje+UnXK0a5oZMGxbTqtfu4a6Abr8tesoswH/+rjqzsjAacARgHcjgyBwKA+bTLTfqJs9g2faZ5OFWfGQN21j9TLXTAYMmksA2o58uBbgmr53m5O9Ou8s75d/o6wBiuRn5My62q1c0Ha0A6sWH8IsJ3gOO09AaeszbJIhEwC42fzyDDbVlAsyD3KJzS1lQD60Bfdy8Bt500fpnyZv5EZ/4EB+yIC0U4lxRb+kDOZi5Q36jO9/+guWFicCufv5/dON0r1TjT4pD96Ejt+C17vlkczrk7KkcJ1EXM0Ksx6sLDweZPygL6r25eLqN44nx3oF9h8QWUEdFgWyNTWy1zkoB/VCJvRPQHqA7buU/lDpYhYGF8muWXfkg0sp8rCD5yNjnoV8m+XB4qMV7BmQ5neUaKtVKwWuWfJz7zyVGvlEJq7/h5qTueXO6Ds/8TfTv+n+q9rPrynDXu9I+oeSX9z2C6nfeE5gK3POogA7QMpZAX3vr3l0OTWaADg75O6EeVESzP2l/saCtECTuHzBAu1j61QQWf4XJcY2890EdfmV2z8RvvML7+1/PL5trBSvxXS+Frx9+HX+d5w3+w87Qy5DeOWQFjx/vlWNev9dI871l8KBQilMb02mUhkBJIlqParIZYyMC9xKKiE/UJ5bTPiu4gu7U6VaHEtx2026ibp+P5dMxFPppDebkVFGfyHTHJ+4OeooP+fpg5DJn1RaAbxfPJj3zG2OjdH2343gZB5jzoKoYz4A/Hyb0tUd+V30a7GQ/fixPVuG5gcL0yIvcN3VeXxWAPxndBJyqDkW28H7TjKggzBj/mFcmvVaERc8Otmn+B57064zfqIcHzlfiReH064rzfyCAOQwqEfLms0laqHVrrO8J/djC/uKv/GoXMEPyGbpjR2atZT3tUqQbGblttHqv5TrkD3zCDL+60rv7MxEECPuinjX8G5uus76XpAmGymsxpr6y77S2/7rlyae67vx2ymv+pRXCnd5cbBb0L+b80uOglg7FcVrcQYazrsPfF0hHlJ+f2NxlCQrCzcbVmizIxqvWF9VyLNFWjQJYFwr6S/uoLJqM8nclTFCZOC4jGGa7/OQey5SZn5nzUCfHZNlxSmVaVnuql6rWBCZ7ZmjdyqGhTOsuBsEsm4jK8gOmWJFwFrnomSFPbdYqtXFUExVKvXj+kvvG0n53i71FF8kRp/4OtlPhLCtSREtvCNWrD7cuJZJ+RPE56jXg7pcYDm3BkuhCAvGLWsw1mzXiKzqV3BwkRYFT+W/phz1NK1r5KqsWW71hS0DwfzY2b/fW3XmlhjXvNs56EMoHDC/864irsy6h1x1qanmm+6gDhaudZ4r3Ng4nt99SN8Xhxqz11T9DGtHrE0gQHmH8D5tX1dcLOvu+YtLgPUARBOkMWsB1iOYTTuen7wnbLjDi1N5uQ1L7k731ML+zYspBYyuJ5LBrGIyjJ3ZP1YS4ZAS4cBL6AbFdIgGxxd0b+TIHdOkXDP5oYJZKZj2AV3TJ/Ce61Zeijp0blaqRKb001lKW1PTzowl+iRrtQvIrs4bm+SHuHdZgSw8/42rD113z+Gn+8eWNiezjR9QXx3Ru/mA9JfoS9SXtRTvf5RGrE/xviUxds2ylfKwp6AMlBkCoum6U3ndKmuR6/rGin25vupMaT73UHEmr9Be/nbF5WD8Mp+SH++Wo0qMK+bWdoUaqwaEqEgfWUM1K7KqI2G/IwfWiO1r7E4RdL93JdCVQFcCXQm8iiTQJSxeRY3ZrUpXAl0J/JlLgBW2afwb+AogyMabRTpgNH/ZcLJZYOEPYC2vDE3gFRCTPNCkQjMP7U0W+oALALsGZrKRYJPBpgHAk00E15E3B0gd83unNQC/sdBn08Rz2VxLDUyuOHJX6dqVrU4rP54J4Gna+z+qz2xe2CxQfn4nL9OIJ28D1A3MZ6PFswAIDCTnnGm7s0GijIY6ch1AtFksAFJ37lp4XjtIQr6AEOQByGFa9VzHZgyXU4B8AIhmAt+eJ8/iHsuT+2hD2sYIn1W9uFZdKLdp4HI9wITtrIxgsM2YAfnIB9nyLOTOedqbMnGezZ/Jur08lo+1DTLi+UZUcF874Il82RhyDtkYQUE5LTYE9SIPgBXa56RTPpBX9IZNTm2KfGljI3IoywW7RirTcRhJZYQK/dFIM36baJWFvOlHbDyRG20EmMN3wAPuA3xH85++DeFHe9DfyIf7zd0U+VBf6kOfRPuOMUadKbf1K+ptVh7cT7kYl/xO/8CqhTFUqkVO+shyNF0JQlfRC/oG4tLEkpO+ZpMzVd+VOFp9e/CN6tbKidqCl3WK2VxlIdlzouEnpObrHgxcH/BvjgDb+rveQZuYSwSeadZEfDYNbfoGdVnNYwOBtxlPP6bUbqFAnZEvsjIrlGaZWqQF+TNeAMBoX4C15iFA4+Yns1f9m7OJof9zMeo7t2mhce5otJs5Z80hy4udd/iPV2/xn90a37tiRVb/vaZsn1lO9PzEqez4Pz+d2Xb34/23t5N6zTxG6tMjdyx/u+emLU/dpeC//7A9ZkHbQxhLyAgS5MhosLC4q37O1bPyD4e/PvDv639t5g87goGfUczda71Da8gK1ejLisv7X6pRoeep0g8ecpP9Y9XkUL+82Q9oxusTYFkRkJn2vURNuthlATAlRa2opNKJbCrhx7VGOelK9TyX8k9JU/uMXOHMJRKJUPfQHyErLmhv+oBAfyM9IUrXO2gz+iUALW1uB+OW/k67Qub8oBJzO30XwKqdrGAMcG3nen5eJMQL9VSiPDU2eHD/jbvu1ucfWacQjDtUt8nHNFc3qrFt7xJIQEDZSJQeE1MxLxdafQnn+uFE3N/nO/1Hys6cGwXy+xSPqK0LAr+XPM+rZmSyou53Nu2NN0ZSrz8z23jqZOCUJ0VabF0pxGpR3qwvWOJANjK/rTm+V1YWypT5j0JBot+txDzCQV9E4xi3WxAVn1LivX5c6buyrOisy0a/Pzz4JsZ2qRA7+/1sPVeLM6P1OFOAsFAQe0fxNJz5UcXhPRf69cWEsxj3OdcVDzhyJ/UmPw6ZX/+mEn2vR8QF9Ws4990RQT7K2sIs9Wrq82rV1bUBxWu+iy5BVmBtEWvempXlxGNy5+XcXnioojgf28/Wto3uzh68bmt6olk+WVnAX7W7giJ/yoT10dnLudjaPFKIRFi4w/25cH6pelaBtl0RiWkRLm69Hg7LisJXnArqMK0YNYMiMLICpAnCXU0nE7OMfV0rC1RvMYplghLJbOT9hLFwFlT+poVqLcreMNvYFA8kZv+HXEBd15eYv45yY2HBvOVF0Q/0LFfriSDEEoxjpxJEMZZmjF2UMS57QFoodsW959JjwQuF6/pmUkNPH87v7esJl91N1fPzb5x75LysYuh78Qpp1T2+GwnILVQkt1BYWPCeZGyvEBY6IuInBPXdQdWpKqj0gGJPzAmIP57KNBTKyCnPn+4fFSGwWdYU8pTmeCIp4t6R5fqmq6aXBN6Hcom0rKDTJcV2iCuLmSOLU73HRCJMahRtF1HB+p51z8WUGtqrxbxuykw2F1222npGmhe5XFSNHXlk1+Gxa84H/WOLBwojywQR362OW1HsDFkcrXYjysI6mrUCayHeXZSTfQLrMVtj8X5nbWzKI8zFvLuSyi/h9USKyqHwLg0/qcDiLxDPQ2XhHcPaCEWUtyjx3mB90rmubM5numE5DBqjTDlN91ov1pYxZa4hu/3/sr2ge0FXAl0JdCXw6pBAl7B4dbRjtxZdCXQl8PKQgC3AAYMBgtlc4sID0AkAgMW9AamATwAeALL4z8fROyAJ17MoZ7PAOQPj2RSwSGcDYdr11BqwDGKBTQSbDq4BBGPjAfjbCaaZpjkbJsBwyhw4peelQF6wWAlmEQHwSxkhRwDM0MqiLgbQm3UA9TRNsXYSAxnwnWdyD+XmmbbZMMLC6sFfk+F6G5J2yxC7jg0U5SZfIwAA+tgksQFFppA9kBbcgzzNdRbXmQUHIIURLDzbSCY2ViZv7kfGpt1ldSEPI246/3ZqgpkLKGRjcSnYqAFUs0kERGaDaKSFWWjwviYvswAxmfG7ubsC+Ke89CnqTrvZ860OPJ9+iOzZpO9Qqjj5GwYUeF2o1neouz2bTSrybQdTee7FDspGvyYhJ/5SHtrHLAssNgd9hnah3pSV6wB2kB9yBQCn/9FWtCsEA22HzCgXwCXn+Q6ozf03tO6hfNSB9iQvyoUVhVld8NuEEnKH5DAC5FQ1cjb3+2Eu7TlySu1uziUqzwwGUxPD3nQ2n1gqutna8ROF0ZGqk0yGCT8XeJ6e7U5IaORDmS+3kaYsWAv8JyXcAnE95SfdrUT7k89GD/oFxJ4RCo/rM9roHIxX5hGe2dkPkTMa9fQD5olVwsIefCY5+G8UXPi+x9zbH8w7pQ90FuiR8PVblelfVIJY/arSEQFpgYC+8NcO/OMj+XD5sZKfv/uJ/tvpe6vH9spJ533Tn8vetfjg2yoj4ecnewfX/N66EE1MxuB+xQd5TM7ny+9ZesxXbA36y+gN3v5b3p/4PPU+IdKCPtw8ClKgPh+POHLj5VztHiYoMqc/3oizBypRf38pGlicD16zPJjK5ZcVPbkqn1AiIOJMKrkplRK2GcUzshDAb3+PtLWFWkUNJ4rLqqP8UzhT8pN/Tn7+lxSoWJq3YdCbT1+0vQW2BgLSaesHlH5YCa389uPH9QUyg3EPcGYWaswNEAD0UzRfuXdnx732lf7ffqDVzvtksZTPfPmRN99UP7lj05sUtwLA/wLSSedoe+Zuxuhl3cusY13B+ILogKB/vTCmUcHblCnq8ZzF3oRzTkHshw8tx9cu15yxW7JhLeE6O/EtpFgMQT2QmnoUv5BMpubGE+9fErj8ZCk6/uFyNPlP4jhotxjCygR3Or+p1NmXLyKaKz7NvELZGVOQI5BDAGwczC+QFRyMT+YuEvK73Ji/4oJs5AYB67heOhA4yT/ZmptYVByN0f3lWwvFoE/WFXlHlgwSreecyo87d5171Ll67ihkhSLuNPkV+tj/pTTRqht/mU+rIi+q6Q/eYesGyAv3UuTEemVdiQHyYWeievXstxa/74CCgb9ZVglvgawgWDlgPzErkt6qAYXN1VhU/ZYSRNBlrSuwbPryk5NxPpciLsWMCAsChysmjrddXKPibDiKT+PmRUqcDisyv3Dlfcp3CR4ug6poOa3g3KIrkmrASPOArZ+aVZJ8mcumFL9kQQHVR1/X+80ekRXHZS2CtcMqySKrpdd5Ij0qufQTvUsl5iTcYGGNSp/dyMG7g7XUQwvJvvvumn0w+dDgm+4+kr9quyzRFCwkV/70+I/PnMlsLv7e3/iZi5HhG3lO95oLJWBkI+/d1cPFLMd18+oleXnrcqpL2cFmYGzmOteZkGVEUkD8qrVEsz+4cTHXX5kQeVGVy6jkyK7ZBT8VTgm0jxVTYlpuoz6zPJfLLk0VhuUiCmsb1qQbPVBssYN3PH2w02VUZ17vURnfUF7IHj3x1PgLC2O9JxVvYr53pHhtGPjnFD/jcK6v8rhiTzyaGyjjco+1IesQ8mWNiAIJcxzrKvYk9FPmYA76IWs4U/xgfTcvGaST6UZlaPv8meXZXFly6JesWN/do8T7h7mVcbbeO1/WKrET1KvnG9Xy7o6A2zyTtQptUCMGSWdlu9+7EuhKoCuBrgRenRLoEhavznbt1qorga4E/hQl0Aq8zQKazQ+LahbygK2cA+gAZGMzAOCK9hIAG9eaaxgW4QBTACZsgpruFpTY/Np3AC3mbAAuNg5sdrgOkJr8uc7IC85ZHp3gjmnZcw9g9IoFRFAUgrADiw20be9Woh6mnQ2QTJ5oCwL6AlACcrEhN211fVwFRg1kt02JESNcg0zaQXSeYdpWZrnQvilv18Jq3+QYOG5yR7ZsiCgXGr/8ZdMFwcImDAAEANSIC+pvZaFcyN4ICD4jfzaxAFftGuJWBtsw8dfOISMOiwHR+rr6x64D4KN/cFBu2t/cX9DmPNcCMFMWK49ZnnCfgZt8NmLJSA/6FX2F9qQsBlgbYcPmlw0oIAlA5ZATSgXXS0fOwoNcS6Jd6BsAcrTPJQ+NgYjo861rzbrCSDbIAvKjHcwCxVzIoHlnvpn5zfolgLWRH9Sb/mygAjKijNSPNuY66sRz6ZsGOvKZ6+gDgIzcD/EGkQPASnnMigbyKnWmEpVm6vGNUrevZsPigYKzGPb5M4d2JI5sbSS8Ui2dnnD8Sr9iJDwvDXaBw74CQzTB+iYJ1BFkez2ZUR7amud3Alps7CkPbbcRrW3aE8Cg3SIHkhMXaMwXEBY8i3ZcQzq1ylkTsGjywgUK8RBWD7SHBSzeXU9Hn842gv+8LTz9kVPR+Oq6cS4elHC9v6bAtB/ViEb+ZVk/nMsuOY3f2PN36j907o+++ObZB/rl+umvTqco5spxdfWgMz084JwsbL4lOTi3eT3rCsVUeEHyZa57UPE0SsPBoieygnENULNbxMQbb/Sf//Cc3NATaHhfdL0z7k5SHudotEudvuRsdc+c7XGX9yv/TRlv6YlasPe8SAtF2u1N+mXhgL53XCCll8skqwpFUmgEEcEo5Bgmzup0X7XaSNU8b8ZL+oeDqBlgdCnpOacrtcZ5aWovFmuN8J23bLkcgEjfpG+8KIB2ITvOT0tD++DeQ6fN9QdjgD7AXAtpwbjZufaWi367V7/8sdKc4lEcfuCeW0+c3ja6PfQ9CM31yIoJncfC6BtKyJoxdqVAEOWl30K0b0cjNus5Z/JePCTSb2E8FS/IwuLWpBPd3udF1yuowGnfVRR3BYfRbFECNdb02SNg7bTEfrzPvXk6dOr1mjP7QOyU71I8i/YiIUPG+PeUsGgF2CZP+vC7Wm3F3PLBi0gaGZv12Ea0pDfYfC/pskXpIT9zoHyrPOfHMmXytsmqIV2P0k2yDvdFy8mck2tUHII7J8W/tY035Mm4Z37/y0oQahD8k8TJaAk+ktVF/It/5bIxNtYrfGY8fXzwvSOf3BTEyffLndJbIFCIV0HcCtwqtZWFeeo/K2HxBXGCpdqG+uK7b9saPvDCdKO3J12X7URvrdZIiVislCqNYLncKIVBNC4STd7G3GllKCMgAnq5XhDGC0G5sag+e1avrsVsJllTTIz29UbTUkSyqH38Az91Ll9f2C928yjBsTsPWVf0aJz9oOasn9Xcddn3Zdv9f6LPEEdSdo8K45XJ4rcHXld+dPD1pxeS/ZtkcdFcOypg+u2f3/ze/SJQ1gwIy6ctfshL6kR/jm+ijzE/E59h5Wi6JAqdsFFVHIqAcZ5jZRMrWIw+s/ZYg51wuRpvSeRELZEMR+R6qSeVqxfVyyqKd8Faf6Z/y2Je1hiurC2WXrh/b0IxHr5B8G39ZiA+T2b9yNzP+YvhM8w3ppBwuWajHyqWi5sTWdKzMNk/qTKNzp/qZw2ciiL3UDpXX9x+6+R1yWw9k0iHVf1OGVgjMf+Z5Zyt61gLW7lYy9pegnUzv7HGOinXWLk9rz8+c+jBPQ8VpwusP5lnbA1nFiMXDiJdpLGYTqQykZ9MTgS18s6VJWXzYH5gHcna+bJE5uUE0/29K4GuBLoS6ErglSOBLmHxymmrbkm7EuhK4OUtAVbWbCYgK4wI4C/AIRsEQFMAIQAstG4BXgAF2By8WwlS4JASGk2QF2i/szllQ0MebKj4DhiL2xuAbhbxbAbYPPCZTQCLesBOA9I7wR37zgaCDccKQL0spdzqaYACwG9AZLSqyJeNi2m92/MBdpruEpQAQ9tdFLWTEfqpefAcA+Jso8JfNma2AedZZkVgZedvO6lAXvYszrcHYOU8m0nAW/JEtoDiXMPGi00ez7TnGdBoJALl4/nIlby+oES7seFs16RDblYXykM+3Ec+5rbItPrtdyMayBu5kR+faW/aHxKIfDgP6Ej7mussAAsjTNoBHCMxOMdnNnG0Pf2PPoLMqUd7P6AdKSPX0v8ARAEqcQU17ZRf2OQo3iGFbt1v5V53c9m6rv0P9xppQz/nQDa0M4l2MK1AygFxADGBPGk3+t1tSrQjZIpZniAXcwVAHcmLfEwjkOtsI/t5fYZ8wP0ARAifIQl3KkFQ0C94JuQF9/GXtFcBt3sema5FSSdMXReefvTmxgPP5RPzI/NOb/mm9GNLnmJt7gwna6ec/mrNTZwJHe8xCZfxSVtWL+EKSj+vHrQldUNW7aQTFyAPxhaajbT/6mFuoTo03Gkf6kg/Z47goN1fr8S8gBVK+xhrz7L5WWWGtIAA/edKE0p/o/0iQMVN6cnrj9Zu3id3JLOnnHFkuHp8JXiHc0v6mV/XCfrRx5W+9nD+7hNvcu7LfHLbB8d/d/wnbqu3YlnYTfcOvMN5Z/xFZ+LqYWdLujzaSVik6o3jinbtKTLu/VvKs7PXeyeQMYAI9UTrvSow9iPDilHRr4DgaQXXnhdxcSLa3gRAp+Ph6K2JBx8a8uYevMHdz3z6oNL8p+b+I7KXfEKvUm0sjQzmDwWNsEeunerSwlbMEndzOuEHldhdlpuZnFAo1084pbwisCaSTjWRTBxx3GhO2tkl3V8XyXE5ssLcb0FOoXXNnPJDHY2wyw+iO9PyO1VPJ59L1Ro363f6+y+32u6CNus4wRzyMSXahX78YDWTKj93y57Eqe2jw9L+Boyj/693YOED0cB99N8NAcStjJgTKKcR8rzTxoUvDQvtKyowSD4XxddsSxC7whtUDItspR6kz1Uag70pL0jH0dKKi3JXccu9ayT3XoFTUSqzs28kmQ+qtbnHQ3XfFcJi9fiwPhHn5TtKjPfv1UFdmIfvVMJVEvMRc/B6B+Dyfa168/7bCLH4vSrnBflgZeF8buH0+caWxjW5Zz+/LX18h9wV3SArADFvviN3TLWBganHxpcnd/lOuG0dctDA9U8oc+ZeCEH6KVrcvKvoG8yZl7W+scK1CCDyvUqE53uVXiuC4C15X68mtTl0AUdHWXgmrqCwNiJddmy1C2O5XA8HerMy5omX1Y/OVmsNTdJBulxR5F7NpamkFykmTdhoRD0pxSFKKPB2oxFP6doD6UzytEws5uuBLKo6niuyognMfvAbn08uF7Lxd+68Lpgb7H0mSPoQw6tHulYf7FtY/usEuCei9wYOiAreAyZb5s/wgaG3VP/Jtb+aEcHLeIJohEDjfciakPmPdd6fNUm2geq9Yi6hnzGO6ZRfU/p+Sg5hEYg2FWieSyTTspRI059t7WJzH2OiufYTSI9FRSyiYkDkBesv1jq8e2ivg+rzva4f3yoLjH03fv8LE1NHhv/70cd2flVEAlZkvBOYS1E0eH8rz/UEyFxuc+7lBGzuW219klEsDeZP2ba5PZne6ra+oVJJwbL7ZREysjRdqGQL1YezfdU5lZV+xzqOsrBvsTUyawpkZYftPVirkHjPfVGkQyORUpTxSuqISJGdOofsWIfZ2vJi60lCF0n0QSFs1HdGgbr5i4QFsmaNQzttVKHjcjLq/t6VQFcCXQl0JfAKkECXsHgFNFK3iF0JdCXw8pdAy8piBfxfATEAVlmgs1Bn84LWO98BEdkMsAFls4JGIwA3C360Xdm4ArbaZoh8cPOBhQAbBDav5s4HwQCoszkhTzZU3LeGpKBsbRLkOjS72SgDdq7EBKgczznVk3znWsoAYWFgNxsOkpExAKuARgAaPIv6Aph1kgs81srC+6YdhDAygnsNXLd3kt1jG5v28rcTDGyeLAgfcgGYA6BFJlZ2ytDuusmIAf5Sd9NOR/4AwFxLHsQDQE7ImnLxG4d9537KZ6C+lZF77dkGSJtcIB9w12REEW1Pe/BM2wxjmg+IyHM4z9EpV3uWyQs50L/IC435nUoA3+TZKUvkR74AdBAEbK5nnMSANqZe2gmXjYTiGtqbshoJ0SrO+n9aVhbI1LQEzQUabp3o72ZJAfnA8ykLfZd6GPDOM43cQMaAVxAC9DnqzfWQeZQTcI2yAe5ArJHH3a1rkB/ADv0czT8+Iw/zp8w5xhXXkdCin7z3XC15sliPR8VbHPD2hl5Urqa8ys17FeJgLHP2zNlU/0LRy5YUr4I6kCaUKpfzta5r2g/qTbkABQFJ7SA/5gqLY3EpAJl2JVEvQPyf6HjGTn3nOZAzjNNLHfR9ZApZ9j4lZMm8M+a5kdOfnLl12U9XKm766zq3Ruv8fzbe73wk+dvONu/0NQSf1e/XDrrzoigaW+tu8sMqIQDwmuM99c8744NH5GefZl17jE7Nx/0Ly3O9iyV32+mpobHMwlVyjPdW9cJ7lBf9AVDkbsBO3D+lNW0qvob88690LQGjzuHoKq8RJEvno9FP/4vMR8/s8E4uu29njrrDkXubJtinILtJuX8qytv4kcXl2o5sNtWjuArZUiPuP+Ol04pbUkuJsNiW9ReCOKjIQfds2fOXvGpQ1n2yC4ijwycUW3x9UE7PAAAgAElEQVRjBxV9RIn5if69RoZBMvFzyz3ZreVs+usiLP6Ffu9089T5FMhGgOR/pcR7AUuaJml59Kqti1971+v4zBwIEc68uIaEamXGu4ay0D/I70oP+h5zg83rlOM6nRzLOPHM3nQ4P5p0/OGkm62KFJILrZxeQ0m5gvKELdf8hJuRFOWSS17eXa8WZBKDIoB2Z+L0csIZnhpJ3PX8qUBNHctj1Kqnw+a88CtKP69E+TeEDF+qYi1wnTpQFwAx3Gn9U6X1LFK+rPP/Rol3hrm822gfuFL5rnt9B2Fp1wRLQf+Zdw3+/h/Lu9kOWRzdsByujIect5z2NlXS0+O9nxqdCW/LluM7ZA3A3LveYf3k+/TjbyvxjmdOYD4CXG8HK9fNoCVP5jCATkB93mfXarzOKw20jBM632eA9/9TiXm8aTF3heSZg5WFXEPVRTTOynKqLGKipDE6JKJCbesu9vdmchrOiYWFih/GUUXxK3rTSXdOPuDOybJqyRVRuVisBub6qkVUMI5o6/HBuaVirlLtGzm/0BAheGypL7+GsCj1ZIfkU8qpCdfOVmSD8SLQ2imnf60TgNiMT4vV0XQL1/fupvUEczbP5C8Eha37kCmxa7iGd9iafreBOEfrttef95OtOBbMzzYf8r4aUNBnAj87QbXixPk+BlO7dS9twTqHc7RDVW6Q5tTk0wLoG/4KYUHfIS+UDyAiWHsURGa8KZ2v3bbtpjP3ieQ4evD+vSMiElhr0eaQpJci6lhHbXSuZi3BXMY60JSOmmtVlbGaydeiwvDy3no5mVA8Di/bV2n0DJXnNvec+47vx7i9IoYMFpdWb8YlazFzewlxQr6sO81qnPxvVn2emD42tFxayLInoBxGal/KMoLfAnHWpVq5uL1RWZZ1y5rpnTEzocT+qUvYSQjdoyuBrgS6EvjzIoEuYfHnpaW79exKoCuBPw0J2EacTYe5rjDrAlusNzcuSlgyABywCAcc5F5A3YeVcDnBZgegEQ1aNlQs0smDDQMbIgAVwDsAakgRNgsACgC6BtaSZ+cGiA0EwA+bH65loyTb9/KSEzfk9FpOrj0fwJz7DDA3LTSu5X7KC3nC5vsdSgAcPJ/nGpBqG+r2jbUREJQTaw7qz8bH3AQhl/bDNvCcaycvjFgw7X028GxoABHIz2Ja8Gw2l+0H91BOAwaszayu3M/GjI0RzzFgvT0mAvkZUcFn8jNNVcpp/rjbNcmsLmhQA7Kb5jv3IQsjnCgvn5EJYKORLSbHdvmSJ8/mN8gV+gJtyuay0zrC6slf8mYjvSLHKDzjBEtFp3bGCDezNKGPcI423+hhfZ8+wqaePo3sIAeoK6ALz2WTS7+mDwPcY80CMEBb0sf5TFvwnZ0rbWrWQ2yEOUc5kTVtxLNoN9qV+xk3AJBcu0LKrbiu4Tfy5XnIGbAX4HYm4zvl3eXjmadr+f1OEAzsz+x+nesHbx12zy8969w8OeMXzvWnz6UF4nM945c2JA/THNTHDR22E+8EOxnTjGUOG0+rGXaAlfQDxst2JQjOzsPABYDtSwK7rQDR1IN2QFufOAH0ozGIgZTCDOzKHHrD6erufZ01DVVMrBu2ShlYGtzfFziJhCiHzbqntx4nL9DszziV2tbC8XS6v+jkRViYlrWsKpxrD5x0rnt+wlU069szQV1xKGrn/NEoF9c1roUByoHGW1UmA4PUmRrO1f7hE9+fuHfH0+Ea/NCZjLbslvuqrc+Ub5y83X8q/rVP3dA+FkN5c/LPTi85AjdnwlQqN9VIFBqxM1SNE9sWIz/veonkoBfVlwJ3bCbyq7nIOdtfqxd7vQjXMfWRXD7+qbddvSGw+uf+7R9Gn/vAW0/MjPQPRJ77TU1l75KLGsDI5qHP6Znhvg/UMskPNJLSim9csrl+Ubfguof5lz7N+DBrg6hFVtAnPqDEOwTt3XawzR77kD4wxiAtIdw2VJeOTsZcheCxfumRgAcVqD7O+Y67NxmcHs9o9DTcu6XTu3VrKi7Ir4qbUITlSiPyg9hPpJJ+RRODq3AC6jX+FrVFplwNj4oLOllLlfb4cfYpxUt+Tccz36TvaP4ytgHRr0gTvyMvvjIn0acA9n5YCVdc65EVyBlw7tqWzK/YCmCdZ1/xqUu4/olzz7xvRq6gfi/n1f9RTvEhOOSpD6XlO7/5jtseu/bAid+95oWTHx+eXtyhZvq7+pk58GLHT+sHrIJYxzB/nxaIj6XSguLUXCBziIpWHzILL/of+b9lnQcwFu19CFnx35UgzpAxfZqA9RfcpvwvKS8CcOsC+rqCbEdnk0lfEQNSvXL7NijLi/5aNUh7Cc8rl+pLUuGYzWWTy/XQUTyaqFpvhMEPPf9RD9dXOnjn8j5lfDAPo3Xfl67W777tiYNXFZZKvY++aa0BzvRIf2apNy+youZkanXHlWO5tuPT+vy7SqyTIIGo5xeV0GTnXU257QY+MxfT13hf8Y4j0QaUiXcm75+NAteXlFn3x6YEeH9DDNGovNObRxw2nEatLCuLipdII/41B23YVP7wE9HU0I55r39sSUvn2HAV1lisc1nD3a1ksSHIaEHExfLo7tnkiae2LZTns4q/4vI719rRbn1JXra+NEsD5vgLCtVRRtYSrI+4zhRueOUml84XFhr1RJ8CYwfVYkYhm5ykXF7d0juSP9kzvCyLw9hIWbKESERGxPD5PaU/UvopJdaHjHEmm+aEo3psUX5nT+3bUpP1CHsDrEzoy6zPeV90kpVW5OY+QNYVM/XSYkFBt1uXrtaIupjl8Et5V3WIpvu1K4GuBLoS6ErglSKBLmHxSmmpbjm7EuhK4JUigXZgmE0CmxoAaf6y2WTeNSAWEBcgFmAPMICNMuAqYMwKkbCyMeW+duCYZ5j2n13DxsQ0IPm9PbXLDrDr7yiZ1hh58yxthHRLtDzteH1s2igvoCzAGAflpqz8ZWNF/vjuB1AycLz9nWKgBNeZJhrlo5wC7ZpANUA4GuZsxpAJZI6Ba3YPz7ZzJlvqTP48b0ernICtbJqsbO2Egm1wbNPWBDVaz7Ryci9yoIyUC+sHnmOa+fw1d05GBPF8A86tnuRnJEN7XQzk4RkkCANkC/jA9RNKb1BiY0h/4TcjckwDGFmYDIy4QG7kQVkBsPlr/aOdtGi/j03vPiUAEamyKTZA/XzVmfmSuW6iTxiRhFzoMxs6WlYW1IH6AurxGdKC/OjngKvI3og1wBnqgqyQJbLhXspAOfnL5txIHcgJkz9u0siX69jQ8pdnkj/PgrQgbzbKbJgBiJAlf2lLngdQxn2VP5hsxPclrk7Pp6pbionCjXI1NCRPIrlUunzkSLznuBPVz/Y608fkjohNOOXm3vAlgL08D6AKDVvcN9lB3f62EnPBRjbljGHkhYYuMmo/GA9oWCKPy+aFhYhAQsgcng2Y/WbLjMC4/YlZZyx96kNn6tsXa1FmlQSciHY4/1/9bzu/kfn7zoA7/wahIeNy1XT/Pf79+78Wvn2mFhsPuJJbyq+5E/kdzvXunCPserW846emndc8cWjFnYq8zCd7RIVE4c+E+52fEVHxVW+H886O+mFNMaG2WJY1x4R+29n+e8NJYvHxAyeiHYtKT10vu4vW7zbe67V6mIgUUOGFOFk/2shkvIQvbX9nPCftfzrjTD0oD4Tuwa1Z/6Bc7y/lEk6xP5VYqDeC+uxCeV2gXKCujUsb+7RP4f3/4/68gl/nvv3662+eHu1fJSuszNLYdhb7epy+hZIjd1jraWjTnv9e6UtKjFMDLenHkSwrHJEV9G3Ig/cqAY6+rVNmre8QzVjLQFbQD9e4H7vIPU4HYWZzEn0WbXrxPU5GQok06cRjcruzK+2cKwVxSWy4pgV3UZN8MohdvyZGYrHUcLMpb2gw4S8LUFa08zgp4iKrOOdDnuf1JdOFUtodeTqIiq9xNUw7YlkwbzG38d7YUNk769SyBGDuACjEmo73EOAbhETngayZL3k3MJ/ZHHYxUf1Zna+nvBrjnffymvGiqA4fOHDDzm8rxsLk6+efryYbwb/TNVhU0HbMletZXVyn87iK4viMEnPoEfXxWZEWqyRtS5Zp/aVP8A6n79EHL2bJQX6MD8YQlkdmdcq8uC5bdzmyggwJwP3UqaXo7HTR2TTUs1hrBF69LgUM9U3FppjyfC/Zm0qmsgq0rSDcDd/35SYqLl5/7LP17RNf8LcsPce4ZP3Auxf5Mcczd2IRtRc71WSduBvrH8/fuMvZffSMUyiWHQXh/hldBdALwcYYpc9gtYIM+cy7nbquNzcjW95REHLkwfWMa+REfQCKLyqrixSve/oiEmhZWSBX1qS8k7FYbFrr4ROQwArEUtAc1p4D71sB+9H0wPjC1OjumWS6p0acIyM7jYzCCoF5hfUJaxnGJ33sVlllbN77pmMPP/fV6/4grPsQhJCmHPQX2tcUb9rdMPJCNSUX1r62pu2sHWOReRKygL5jlrbi7txEUPfzxemenAgLR5YeJ5dn8rHiaxTGrpnaoWqy/jXChDJTXtaW9Fn6HgQecyL9EhKBsi4q38lqMe3PTAzuUKDv82HDhyznucwvlyNXkHFZPttmglr15jZXUFYvxgQk0Uua7zuF0/3elUBXAl0JdCXwypFAl7B45bRVt6RdCXQl8MqRgIHDbMhZrEM6AI7w12ISsBlhM2BuagCG2Xzwu1k/sKkHJGEzxUaFa9hIoGlufmP5bot4nmeAWbvWXrvkyIffyJf8eRZlVD5h5NSnrnYSfYDDPJPnrGo06zNAmT0PoOsjSrZxbn9u+/M6tXupA5qCgG+8g35d6S8qGcBhWmFsmtrJHz4bOWB5co25dQJ44TsyZnNjWmV8Xm9TZxpr5MvmCxCWOtBOyAaQnQ0SbWTtZi6NDGCnnuRtmp185zPlNGsT4gOgqWpADPI3iwEIIfI0IgRZApaYNhkbRPK/lNUKzzP3TYAbgPRsFNnMrmfhQX0pG+AM5VCM23M7HLeheK0pns/vAE3IgGT5U7cNHS3Sgmt5jpETyJWDfkO78wzKxzXUl/Nsro1IY2NvhAvyAUyH5LF+gWy4l+/W1pSV/sVvtsE+rs/0YfKGCOQ32pNkfYr+5P/J+SA6shwOyZXR2wNPvlQSFTcpeFVa8Xt8L4j7UzMzgi0AjSAazeLmsmTASrXXHJSTcgFgUU6ej3Y3B+DGTiXAk0uq2reuB2DBKgttRjse04ePKk0oXYn1B88DUPsdJaysmsA6KplDyfPO1vREZkvqpPtHMz9Rqsdpc2Hm/H7jR5xrvUPO/5H6hNTsl7f1uYsf/MHkl3//j4L3/KU1tdaXN/Tdm9qeOeYMeLMN+X13GmlFh9Bxjawr6A1R3nPSucBJDqso6jnoq7pDF5IV3COyYmeuUvp/9wRHc9u9Uz95Mt5m47P5WLUVWuSQNs/+4n13BP/ybpSbm4cr1y/hD//eIUXdzkYn3BxtUHADd7csBO6UNYWsHlzHj72FVORMDzpefsSPTu/NOtNvO/tIyV9ejH/0gx+KWuTEioheJAnpa/R1azvAW8b52S2TM2+9/TsvbNt38+4ZBcNu16Z1suWac2LnWBPsHJzFIdWq1wvmIOZjSEPGt2lZ05+Z+4Lf/FtNbXTGFHPWu5QAlLYDuNkRKZ5BG0GkyMJy+6ExJSD4pbjXsHnSSAP6M67u9oSxm9mWCI/3BjXfjVK9OSeuJBxZJHnJehjEhaUo7g+8RKjwH/m076f8pFtQ/ADq0kgk1NKuggt4ztmEOz4burecbMTFz9Ticz/eEcuCfmnkqpG6q3W93AcB64w3+gqgIxYigIzXKFl/ZR60+YrsIHeYgz6rhBUb74QrGVeXK9L36nd7r0OudBJ8mxWI/VaRFieHZhefv37fBH2JOQi3YQC0lyIXKN+PK9HR/ofSP4C0mNi1OXFk71Z3ohFkGskE2un0Rwiftyt1WjZaHe1dybOxJGXualqRXqFbvXVlBmmhH0KIC/11FWumpPgWDVnz+GEUu5WFOTeXiMN6rdQoOgONGx/7Vfems/+rPxlWmAMoO/Mv6wFkAmED4Lx6YP20Y+KcAttknGdv5dIXj6N7tzqKbfG5nuXKfxw7O0u/pI8x/0A88P6CAOGdupF5nfcm1wFWQ5Dzl7Ua5WG9xhhkfXaxdd6asnW/XFYCjHn6IYQ9c0GPnCc5UUPvKLknSmV7HHflVdV+JERYyL1deNZLRPtllcDczPzPGo65kTWprX/oU/QJ2o2/NX0qDmxZSPYMlKcXpwq8d42wYH4yhaU17wmdN5enZmnDOOtcY1NGxgF9mvKsrPNW1olNy02RCxO64uaglpQFSXJcl5eSmSBdKWb25gcq50ViPKgEkUt/M60D1kyMEfof73/WbcyTzMeLyk/e/eLG8mw+K7ICRSZ7ATG3MAZ4R63VYKCkK4do7OBQaX7Kj2Rduc7xDZ3DbeWiCKaXsuZaL8/uua4EuhLoSqArgVeABLqExSugkbpF7EqgK4FXpARMC5y/LPRto85q3MBgNi5s8ln0G1DO9U23CK37jJgAiAXE5eCcbQZsw8p9lrjmYot6QC3AYbNEYLMD6NtwFh4uOsPv6ZOLIGF0vllDkA/P431BGQycY3OFex824ha3wZ5pdW0HzPnNNCn/UKA2WtxoVbGpf62SaYgjB3s32UbMgHvKbRr25MemjXLib5fNE3mYLTmbfOrIhq1dHqYZjYzN/N/AFZMlboLIn7wAp3HjxG7ViINWlqt/2stpbcA56oJbFpMLmzWTCZtbzrOBpE6AZsiX+/jMbyYHI25M9vZg6ytsINHoo/4ALdqArsYoae8XRqIgczawdScKXMUuiZzyiYZTPkg5qKfVh7Ihc/rMFR0t0oJnUycDACmnWZ9QR/qVWfiQP8/mdxsXbPLJgw0x7cymnr5q5Qd0Bey0PLm2nfCgT5g2NHkBOnIN9UO2fF4FHp9aCN26lNu5ThvvPxlITV+7GAzerZQYz09kev2FeQWxBXRCLtQreAnWFSZH6g6BgpY78WIYGyBggAz3tL6f0l/rr3Zf+1/mDtNobj9vbkc4t+HNfcs1FHMMQCIA2S8oAZI50tx2xtMTjmSRliunsuInrxIW/P6x2j90dnvHnWF3xjkU73X+oPFegNALjry/3LTWSCZqSSHUzd+HZxYfz1Rrr83EDcdXDGEvI6hdo9Zr1ytdL7OFeG7k8FTlxt7nDv1Y32d7/0Xu7/1k52X9jYXRu+YeGvmdbR9aEGlROTjy9vihsXf7n/xnH3G/PPtI/+To23fIFd6KKwsv9bOe/DOpDzTFJoi/33Od1FI57Fl0a6WRpTPVNz76815q7qgjwJaxTVu1y5cKYSVFP2M8Mp7eqkSfnRVi+rObz87Kz33KmRwfaZIidiiOhXPk6vEmYSHw1xG5IUuLEID8ASXGyEQrTwvUG0nLPW6B7zyXee4tSt8v6d2q1NeI5O1NXb0RJatzwUgm65Wdgr84LTdBXD+p7y8VdGe87VRiHNB/zUVbRYTPjNwN1dKumyiWaxKfqApfsF7cyCp+RSid5UpBxIQ0kdMaY3XX9YJKQ2MxbEylCplez4t7VPbtfty35EU95xPxwNmaM4Wbpna3dFiO/Felf6qE5cllYyuYnNsCQqN1DCDHO+AvtGRnl7WTFbjyAaSHOIIwNaWB1bbjw0YsANbc8P/PFzoUaw0sLBi7ncffC31v38N33XxQhAVzC/MxcxBjlX7Mu+pSB7L6kPrtuXIu/QkshuYHe8dS9WBXkEhco6HDe/QuJd5DF9P8Zu6lfMgVCzmIE2JWXGqeu2JptawtHNy35R/7RFhYOpaoJXr8xNxEIr9wJJ2uL0RxrRIValO8WygzfQAZUAfIWvrHBQexKbCyYHx2EhZcrFg09dnhXk+xLiZkLcY7h3m+Sa6v50qr/QGZtTMm72fWHrjh4Z0OiI5caV9keK8S6x7m6ysm7a5YoK/yG1pWFsyt9ysxb/8UVhUE325Uy04oEF1eAk0K9FXWNBo/7iHFf5iplVKHRFyczg+Wb9N5LmTNRDsxd7NugaBjTDDGjFgs+clo0/ZbTz9x8IGrDsrqYY/eQ5o6Rc+GHu8P3rH0oeY7uO0gH1vXXqxlmAuYp5njme87lVfo98dUReqqNZMrD1heff7UQG+ut1rJDZR7RFhAzrKesvU886KtW6gn+dP/yHtCZX42jtytIiwU3d5HSaf9gMTBmgoSsLM+XDfdqJS/3SgXP7hO+Bd8wX1NCZm/FIL9YjLqnu9KoCuBrgS6EngFSKBLWLwCGqlbxK4EuhJ4xUrAwCwz/zfNfANO2XyuOJt+0UWCuYthw2puE8x1AN+NCFkVSkdQ7csJy0BgwAc2UvwF+JQ350cDZ/lgyclde05YHc8x7UI2SDybjZhparFx2aGENqX53V8PHDWQHXAEcAtQdos2g+TJFh2A741KBgIDAprlicnLyBs2X3wmUW7ABbRJkSHabJxjEwWJYi532CCyKTOywGRKXpTXtB2pm5EgnEPDbZcS7UG5KacRHO2khH3Wz6vWCMiTMlJngAXqidwpB3m0v3upI/UAmDBigrw6j6bGaOtk++aTcgPKswnEBQCyg0wywMjkb/XmL5qZkDAHnKiSc8KS75SeM2LBrFja3WtR9is+Wv1S/pljs8qhTNSdMhgph6w6rUjMsoJraDeABGt7xg4ApaEH5G3jizIaqce9XGNys/utvZpjSmVsgrYqoyvCguv7pX3O868bELAurfTFkeS5c74bHFFiPEDSQYYtfJcgm/Xjb/EspXZ13X+k7wAF/7cSY7QTWDbijDGIBj9AdfuBTAFM0BjdMBDY8huPXJAhQDna581+L5kMY2XRiFPOjsyRgfnlTsVPx/m12i8p3kXdKcV550S0vR1gbpZNcnQGkgLi3UbTaoMjW699e6w0d2Bq6+CxwajYmxoKb1erjXgXZr+mgqH0+eN5R/G9o1/eMnna2TV27HDPNaVw2c+vAUoXkv3/6kDP9W+6dfGZJ57ov/2L189/q/6u0tHEmcymnp8qn+wTmZH77NYfjb7dfwcyXzGPUtEErDfLWAirX8k5tQd/7ORvLXx44r/0pspn6H/0X0hB5gj6JlqnlNi0ZBnLgKAkG+s/CdipoNrO1slp585v7XcefSM81cpB7AqOp26/2hGoPJ8vVY/3zxcfEskBqItmqYGSdYgKrlV7cRPzCWAmGq3MxfSHRC3KOgvBoMiKNH+j2caoYobI+5vjHZqs7Tg0mjwT6Rr1oyuOXWFAGGMBcQHiMx6bAJZcPr2QCBpTmZSXz6WS89V6sCyiYjGhACdy7KTqyIbClYf/MArrQdSIG2EjmU4OpTLZRkLBkhmQCiigEDLJak9q96FStN8pRz6EwYdXhbXyAVIPsuJg6/nIo+OSNV/b507eMVgEAFIz93aOH7sRq5F/qwRZQR2ZZ+1dfKln/Vn9Rr+gn0BYfkrpg+sUZERWAH2yyplXbBXeFfQt3lOQY8w5H1H6mxergPomk+YvytLgF0en5p+ZHB9+KleqvraeSgyJaGPOMXDzYll8RT/8ohLvIMZS7bsgfdc8o83iaWWt8qu9NvcxTgF4zdIR0pn3CmOYa+jLF5Cd61SAftDUgp8dXt+AZH6wsO3RN9ww+NzNe2Z+7HfvLdlY3UiHID5Jm9s1ytVuVbhT3yG1sdZCzsw5zP/MOczzFd1rChdrHneJuCcbKdafp2t4z0KgoQRB2gphEcrKIlJMBawtXF+TqOueFtHKPNCjANO9i+d6fcVteEvPUOnEzoFTuIVivcT6yaxpWaNOKLF2MGtR2i2ra71NV03vTKSD58++sIlONVKvJCeXZ3oeV957wsAf1GzfaS11JW3yOV38AaX29yLjgzmQde2cyvAXRB7nZCWiBU980k+F8oQV0c+xNoEkMwsN1gXUi3U/fY26kFhrh8qD8rPuQobsbSDcmGfZHxjRgFwvICyiILi3urwwLoZIxMYF2wjmKfLoxm25kpbvXtuVQFcCXQm8SiTQJSxeJQ3ZrUZXAl0J/NlLoMPHrRWoufoWIGqbZxb/7YCzgZEGVhuwbJrg3N5+75p8X0KtAUcnlNh0sAlg48SzKk5YUcxcKXUtPpJ2hlbV/diMcB0AJO8MQF02EHymLuY2yEDn9UgLzgEavFmJTTjAGt/RsgdkRx58J0/yYeNjbrCQD/dwDo0zNj6AdPwFQEI2AHZGqHAOosHcOOFOBSCm3WqDa8mriU+2nk8ZbaPFPfwGGIm2JRtQ6m9Auj6ukklmjcD9poHGpu20EmQFgC+fKVM74dJ0t9MqB3/XkxtlaCcejMRqv57fAVzYBLaXE/nRVu3vecpKGZAlYMeQUz2ccmqTc875PwDEQSbmioDPnJtQos+85ANri9bNocaBEUVmTdJJxHSSMrbRNfkYWG+bV85b3A4e026FYi6u7B6T2wXADuSKAB9XboZS+ihl4ejmcpR3b85/55msLw/oUbKR9qrmfswspq5IJusAUha/AyCMg7Fk5B9u0tBCpp24rp14oM3pPwAggH/tx//Sl0eVyNPcXl1ROVvPxJXJf2vlg6/7JtEwkjzrvK73PudcfbyilJW8FDLZa46BI9G6Ssmrz35L/x87Y6lJJ+2uNF06bnyr3y1NjPUvSLm+/K3UeNzvZdYNIL6m/JAVzSgi6hmYxGTkpv7GuX2D7zvzueCT2z50gWb30fzu9y0m+/amovp4ycuOFRqzzs6wNHkms3nLo/2vGzia2w1w2Tza2cfB+vzhu+Yero3Vzjo/e/hf39LXWEQjHyKHCnxMiXmHsU1brBf74AK5e1Hs9BQrzg3PHXME+DpfeB+cxtrj1PZNAJPH9fsDg3PFo0Mzi033MAKZV4iKv9Xs44xtxj3p/UrMiTtlnZAIxbedrY07c8Gok1Xw5fONzUHOW5a/juCFlBs+cqq6K3y+dBPMEx0AACAASURBVFtKhiMZ9fma+uVGXNS0i4gxyfOxdADwNkBqUiTP0cFGpVQPk+5A0l+u1YOzCoB8TO6etuolOCirETcI4qV0IlHQQxMCv5vu3EqNaCgZBku5VKIujFB1iQteVIj8cHg64eU/G8aVTsKC8gDkQfjR59ubrlOkJi8DrgF9kRvvHoie9Y4v/W/23gTIsusq0z3DHXPOyqysUVVZVZJlDZZkC9mWLMu2DDYGbBrsBkzLDwi6oaEZHk10tx9taBoc8WheBPAIXtPB5AZM22awMW1sYyxZkgfZlm1J1lSqMVXzkPOd75ne/926K3Uq62ZlpkrCqOqciJ335rnn7LP32muvffb/77W2TkKGMD4C6C++UMD6Cs97oU4jB2wsoeJ6HRbicVz61AkJJqDfvNSwl3hXAYDzfvAepQk8gRL5ymgnEmdhZMCp95Xk/RM6AudvlmfQNbWBMiGhbBy0z17PZvX6bygxvvIOEaxHpipnr3blebaggvalDoxd9GnqSqL/sMKbUGnYNUJ8vU4JMop3i54xaHpU4NMaGvbmw6jgxfHr1Jdfq3CBAL9LR+x5r2sXvdPtYv4RyXe/80cfW0/fWv5Ie49g3LGV7oDI9DveNRjvqQf1htjseHIonfcuYSRIRlz0aNHzTyE3I4kYQ9+55GXRqAlLT+RlkfP0rvBYrtRf0me/JF2vzfbvlGeY9t5JNsjDYMr1O+/66Ld5nqF79CfeTe9XggxAL9FdgP49Yztm+0a3LlTlmRArDTZrhZH5E8MfOfbE1jta1cJbeSN5nod5DnE7ZbKQmujTm/Wuc1LPTwbGa51Nw0WenCkNNjfp/Jie2dIn7/+UnT4EYWFjHX0OL2lsP/XcQj6Sx1HdZ+FvLbwpz2a8YPHQBXG1+FEeLIMKBaV69qwlxArj7nwWDup5akF2WyaBTAKZBF7CEsgIi5dw42VFzySQSeClI4FlXhA9X8uZHPHunqpVB1hdgQhZd+WTz3ZWVQFkAryxMopnAb4xCWEyNewc+q/HnGt+C3CdcANM/C0Egbl/QzKYqzpgvk280nWy2ZWRMJSVCQ55EAqJerGinIkOzzYQhQk4YDplYyLE5JuJEhN3vlNGgCYmToC7TL5YBc59TKq4xlYAT+o7YBorf8nDyA4DVGzVGPXjPiZZlBEZ4QlBmCry4jdCklgYrTSBYOB4ur4Ah/wP6AisCpHAnhKAzqzC5jfGXvLl04Do9Iw0nW9armkvCZMtdaNM5IfMLHSVeZSk7zdSAjly7HcaR29wzv4t5AFy5zxyQr7IhXyZXD+O7rjf3pnwXtKRIi/Ix3S99zS1+6Ruv1jPjP28/NbRf9TX4ryICcUL8c7Uo/7t2vr5iID6uU2l4/3ytmBVMGESCGFy0TKvUUjIGN1lQs4qcmTNJJ9+xcrG13TbEzDKPLHQGfogfRjCgtX86QPwysi751tG7qOt71cCwEGHfxiPA4XEcjYWTjvvmviT8kMLdwsM3+odbYL7XvyArNhSPKKCRR3iYyKcrw3G9V3b29OF3eHJXUUveLfHls0XOVi3GkkSiUqWmEXQLTmp/sure8f+/cHfdt4w86Dzr2/5wwty+ZMdP3bjm8/ee2MlN+AMhHXnaHm785XR1zofvOoeZzZ/YYSK33385+d2NJ5tXF95+n1D4cK2UkQ3Wzq+oW/YFQ7sTvoAKKb9lh94IuAF1tlQOydXA4GeZ/R9WEp3XlxvbcC9ce/1O5/Yd+2Ol5da7eNX7zvWuPPfPJ2IqOCwtqWvQ5KQ6BvvElmxqRn3OafbW53jrUlnLhx3pMt8/5zabXhT4fjDOve5uXDjTe24SPkBgSAt5gRmrlVXeL6F3euEulI6qgQJ0IgcdyZXKra9OKjXGu2K9g6Y83y3pu/zIiIGxHA5DYWGjxUOTP3S9+IwV22L0tDux6pQxW0FC+0wmk4ayWJfuRAVnZ3zSfxlXdwh75avgsdLDGKPsQrbhc4urwflJdHIMGqQTIwdEH29QpMgY8afP1WiD6JpvfLlun+uB/Uj7BJj2q8uKySeRLTb33Vl1pAXQGfhgQgB7BH9/b6jOyb8jWcX7vPD6Hu1YfdPzG4YcvTpaN8KpzJY1ubw1Y6XQaNcLMvromObIeME4F8gE5FU9Imv67fPjM5W5jeenc/tmDodXf/e4522Sm1Ub223/F2CcSjtnWfEP5+8D/AOYcSFLcCAsGAcB9wHfMauMg6/W+m/pQq5WuA5u/ST+gJxVZKX1N5CKzys/jsXe/4F+/ToGvoH71DH5PVTu4SxAjnYexrhdLD5jAOQpOgmfRh7zzsQ73UYUPoj4/xa+3NKFFf2V8DwW++8B9lhT9Cnd5pEWrVFgeqBMzC+pS+J47eIfJ2RAbta4PxM0Mo9qb0fnEJfe1L/o3/0J7xgeN9D79AxbCS25F3dPGknruksBBIXGCsEk68kZsQJS0PNO/uGG18c3rz41cf+/oY/CNu5H9d19IHVPJh6NSILb2wxitlDrpN9cLV/WbJQKLcDeXmM1BfKocJaLcrelkS7+NpSiPcNdIkQVbyz837LOyaEB3bGFl0cCZq5b8yfHN4ibxPenXt5UvQkK/R+13Y97xXyZCk+t65rqRof1jdsmXnS9qpfdi6TQCaBTAKZBC5jCWSExWXcuFnVMglkEnhpSWCdoZ2eT+Ww+bYalUkUE4gjSoDVTGTqTu2JqjN33wPO6N392seCSQcTLiZVgANMwJgwgd4xUbZV8pSFSQ152ETZQHcLoQEoRz5McpjsAHABqHAPKwgtVBIALtdynok59wBImOcFzyYPiAXzFAC0sBW2tskgZSXUFKQFHgKU28B8rjUPEeoFYAw4TJ4HlciPMvEcJpUA1aw6JT8DhI0wMITG0NbORrjdvACWARaoD7JKe2ikJ2+W13LAxggKnkH+RnKkn81vyM5AnTTZwfW2+pR7bJUm3z+vQMnbHK94ypn9DGAfzzKSCJ1AZhYOC3DrW/a+0CUc/ikAmGgif/Jgn1+9YSg3f7wVl9z5YLz9RPXb4psGvrp3Q+7ss44bL1xiKCiJcukA2ELfaCdWHVtIH7sAMGxSyTxd6EsAD+gqn/Sh5QegI+0JuHapMqOv4XX0ISWIml/z3cjp84Tf5hLnDSIh/naaRdgXP+7Z/P85k6V9KoznlLyG8x3VrzuDcaPfT6L+DVGlVo5bFyWjkprz5fiE801tEx3oeztpOb/QgS9S/Ia8J5wNwawz0Trj3DH7kPOlDTg2PXfU/H7nh2/9C+e7Tn/SGQwriuUBLuQ5c/mRbngqC1IlI9eedq6p7Rt95cKjHUA7H4dLIay6ORpZ0avivcgKwCnznOGepwV4nXbj5AntWVFeHOrHe2BpZboA4Emlt+ncQrNc+NLXXv1ytSXRiTp9GftG22M7AWUnld4JWREmeWcxHOmE5cKTRRujaydTbREejuZFUDSPtnYPVqPBV4mMk011/4Xuw65CpHxTpAVlNBu6WpNiCwChiWlFuW08oEWau+dOh2dahdbwYOnMQF8ROFtkn9cs9+W0h4Xj5qO43HaTpi4eD7RymABhas/2bORsHSWciuc2tUFyEIRR0/NGW65XOiFQ7SvKu1fYnh/RechkCD+IvbQXm8ibbTntmTJc8NrfL0zwO/Q7JN9hpZXICuoO44UNpI7kfXEmbTVp/dP/TnkZs7AFaa8tK8nPd+u1X4D6MQB19vb4/dT43V9tDCvuW3Xb0TP/XTukf1Mhn35VhMR4rb/ozIwNO6WGwuTgdaH15pZpL7JiaLE2e92Tz+7f8ezpL7WK+c+XG60+eRhtK7SDAREV2ChbYGAUJDpo7xXmtWmeMbwLoP+MsVxP29CmAKn/WwmSgMUFkFu8R/xHJTwQ7rmEJkC/sL+QyYDOT4hkrCusFv0Z2UIo4DnaISN18M70g93z9C107VK8LJAH7TilhBx4DrrLOwXf+TSvEsqJVxCEqoUdvYSqX5G3YsvQHd7d0M8NcSSTIjX3tYdFFAVOoTSA/M1+jMqrwhPQf+bkvokniwOtaGTL4oR27UFfLBQpdpY24p2PNkMfLMyRvVNjU7HpZ9Uj6hqNcsX+9lvltfDAwFj90MKpwePss6Tf1/seZvaZZ5M/esH40e23ST1fDKPyULOSK4QlhaHa1qoXgvJgM/ByCXrNPIHrsfU8n75pi30IsQa5c0Ijx1fCVm5E4awkLg3y5wg0FuwgT3SYPtrzUNitpvauqMXBeYsC7FqeNdnN76Vmh1eqcnY+k0AmgUwCmQTWIYH1DnzryDq7NJNAJoFMApkE/jlJQCvk57RSnskTYAyTbyZltmIWIIDJzIjTPJh3klArxXzICkAbVvAxXlioJoB9Ji4A4ICutgrLJhTpsBDLwUgAJVahAT4wETLPB7uXPAEiuI8yMdFiAsQKL37jfibuJKuDrTrjHLMe7rFQQ3h0UF4D/fm08jHZZzIFyPiAEuQEoUBYzcZ1lJFnA4QBfDDhs/qkyQXOpZOV91adhwxhCbptpG3l0Kml1XLpshkZwe/p70zc0t4dVj/qQrnShBH5GVnBeQt7RbmoM20muYQHnYP/mf+ZXJMf8ua3c+TVOdALXRlDdyjQZX64WpE+XIsGbzobbL5dQpxQeJ0p7dvwzGI4mjTi/tMD/sKlgE/LxUfbADIxsSdfwIt0iBragHX16PDvdNuIPsjKctrsvJX53bwAbgHKzsVdurSD8gHe0DcgVtgz4JOeInwV3abCxHjOrtIzzrHWLm1Uvbwo5x68uXDMGc1NS6Fip19sw1XBSSfUsk2RFM5A3HBKcXDxOFKJ8xm35PyO9rSoipMYU62fSY6KdA2d/1PZ069ZQc1xSETElj31g+X/8sx/dd533a87D4/cJm+KqlOVVwVHXRjjX289t8B1U+u0c7r43OLqtJF61cI3nEBODzm5BEBj5DpbsFzSgc39GyX6E/3oEwJ/ta10rV5sBqO5vmgxzPkwP+mdO7AXb1TCfnxKgDIAF7LiHLYIPViKbU7IEOltx3tFocycWjzgVMKRp7TZdl6hn3IiM+aDJN8UgWHeZthI7CXAG2AUhCx22bwnVqowtoYEIIX9pUyQsowTgKWV9/ddk7yvvj/YuXWkqn0ppuM4OZDP+SUJUxvKOuUgjH0nCBI/n3cb2vS11ooUxiouFPI5hQTLb5ooJHuTIDweBLHGmGFtTLul7RSmiMWOffq1HgX7bp1DAW1/GUDiWRGOBW0Qf42IqbcFceEOhcS6RV5StMUNaldIPfJLH4SXgpxDFhCIrEzuiaKtJBzOp/YhsMtMvYxMTt++RCpeasie9Mbf0hf6LXVgZb6R8ennIrMvKtV0LXYGXWD8Y9yYVZinHc1ycezsxAjjwhZ5FTwtT4myH8ejasc9B6/pxZWeL5Xrn5xyFM5sg8iK2/urzVfII+EXBfYjY1ZNQzTwLGSNXOgbjO/0AcpN3zaiAl2DCADsJYbaTiV0Dn2ln0Cu/1sl+gQHNnN5255fuJX/+4x+ghxDP3g+5eW9iOdMKQE8t/Zet7Ot8E/8f1/3HGU3cJfceYfgXojANY+dy8IGWinREfo/fYx2pQx4CiET5ICt5zu6DWlDeembXGuAseWVfV5EAl0vC/SKY4lkhrQI2g0n1v46imXYITC6x7n3L4VCmj062t+uF2o3ve2pQ/KOwFMJe2R9Ht1Ab7GdnXBoSkZAGHlBlrxzc9AvblKYqVx5qPHIwunBRT2D69d7sJiFPoV9tAUz9Hfeu9Gj+XwpmCkNtsoiLYZEXuwR2XJWoaDOKPHeATk41S03z6ceJMpMn2UcGRRhfn2rVvzy6QMb2XPjh3QO2dFveQ7Pu/BIkqOKIVWXZ0W5Pj8t83ABH8Ecg+fjrTyXhYNab9Nn12cSyCSQSeDykEBGWFwe7ZjVIpNAJoFMAmuVAKvGmOQ+psSqJ8IMAMww8WCSUXRO/1XFGX/HZmfzPSzrBRRj4mCr7w2MZwLPZMhAdVA9Jm9pQN8ma3YOEIIJGxMYJmyUhckhoBkTGyY4XMMmhUz2GKNsBSZgBCvWmGRxHWCCeQwYkE9ZDDk1bw8mgJxnNmReFQb261SnDgA1rJqmDkzwOceEjHv5DigHCICMAEKMnOB+DluZDABjMaQpJ3J+uHsuLQsjTNIeF0Za2G9psoJnpL1X+I17aQvkx0TSSAojj6yMXGP1Aci2ME8N58hv5p3KN5AjE1rqzbW0CzpBPdAR8qGdLvvjZX2P+yImrhMxIaIiFyt8USSyYkibTec1IZ/XSvW5973qf16q18JyOSJnAxcBtWkfwjxNKQEM0J6g7GxeSVgSrqVPAt7RZ9LHp/QPMdrpX5eMsnczpr7oPuWBvPo9gb0/k/faihcROa/RfhZDuQVtVK3NeKWij1Ru1/ec8+0bPq7V/sMOq/77tX/CRDLr7AxOOZvDGUdeFc5QXHcK8lyAyFh2ALyBhkK8HJT2HVLGD0uDYxEX+fiYbmh1dP6zStgEwAy8QP5GHhsTW5on37+pefruX9v7K867bvvrJbJi+UPSZAW/WaPuqR10XicPjZfVnlFDRNqDdNVFnch7eVguZE896FMQrYCHf9ItJ+fOkQKJ0671l04qEMhKe8SQL/dx/IoSNpcQSNgWgMnOId2U60lRoZ92OgLpnUo0Ehxp7n5gPhz3pL+xPC0Oqh0a8qzAYw3Qk5WxVJnnAqxhW7Cb2AlbPWvZpz/RTXRyUglbwf/c/1UldGNpL5kOaXFgf7Bjy/CivCWO9JXyse972uDVWYyceMBzE1+E1+x8K96kB25o5orthu+faTlerR57czvz3uGCE52sN4LgzKE3hQOveIh+grccYwN9IX2g7z+ldJfShxVsC9JRWZc2KBTWPQqDdaO+X4OuDedmHXlcoLtpUt3yguhARkZYmC3vJYsLzi0jKowYZ8ww2dJf6UsoFQk9QGbmhXjJtgVPiW67UD9WPzOeTnY/zUOPshNPnv0k/kAJ/USGlBO94ntDXj79SozXN8nDgr5G+DJA1xUPQkVtOTnrjM4uOuNnF5TmHW3QPSE0coJQaDp450i7ZQHm8wzzErS802XlnHlhrvRsIyv4/fmQFZA3/75bFhYa8HzefyCUaTPeB9D5mI20f+dnB5ER4yL6yO+vVaJvpJ/9S/r/S2qThsgkyr+mYwXiij2WeA62DjKFxLiNfcEGomeEh0PHKBfkBV5xgMrYi+xYuwTMsxSCnvBG6GbHYrYbVe1j4SsVpv18sS3vT9qbMfk75GnRatUKfxo0881kqHmrAH9j9eiD6QO7SdsZBrP8d67tEwn9cXksCMwvF/XsKZ2jb9o7dppjX61mae8++ri9Ixfw2lAop1klT6Np0ctHrkiLaQ0pvPOzKILxjfdj3oHRKWwV/YB3SUhk3kMUycmdrc32udp/49WFclCQHO7v7rthodmWl7EWx1FFm5k3arOnrw1bF6yv4Pks0oCwp+70x+zIJJBJIJNAJoErUAIZYXEFNnpW5UwCmQSuaAkwAQAkYPLLCiomugBjrI4FYGfyu+DMPzgiwoKJGisIv18JUKGzulCJ2QX38T+AtwHoCLbXKlI7x3XkQx5MfJiUMBliRSX5kQACKEfacwBgh5WKtioY4iINCC0nRoxAsJASBvab14Fdb54Z5E89mMj9pBIgHDKCSAEkY+LGNZSXCap5M1BfIz8sL+4FxGBCCqhAaBcmjDbRXA5KLf8/XRf7LU1eWF2QPe3DhJADmRpZwf/UnTJxDTLlPtqbT+T9u87BX3mLPpHJlBJAEqAjKzchWajvHyuxPB1A67I+APoGq7818L+qP5Icj7ad1krsAwI5bxjy5ysCek/ta9x45N65d0Slj/6Xjhye72roFVbQ0gboN7HWIYuInQ04nQYlbL+CldoBXftzJfSC/nmeXq2lvOkV2sseQl4NyQjd+T2lAyItflwr1l8xKLLixv6HtaofzCXRUuwj2ux5o0I/1Z18vq1doI+1v6/+mUKsmkBU9MurIi+PBfYlfS4I09LTIGQ+ogRQyDOxEW1pdeDmtL/BHvl9PbzU7/9MvwFSGthL35wXafGLLb+4bUN79kd+7MgHbvvjHT++LfDySejmsDsXPbQPhvPTh/97h7AYa8+myIrzREk7PdstI/2K1dh4edA+gIOAhLYPDIAXnin0JfocwJYdicLjJPX+Em31j0rYlf92kQIu9yzAfp9zHeEBIoZmA/hVBR/3GidEYBTacaGpT5E7yacl67MiNgDk0Q9AZwhhCN83dssMEIoeYk+wfcgT+2GVRxexL9gy5M7v5EedSciXtkh7aCRHTi40t4wPzERyoSgWvAXfc2Z93x+PnaQZaE+LBQF/+Vy8LZfPDVaD5PSJhjNfd91w0Y3nNztBa1QblLzvntsIWQQIi6z/ndL/o4QtY+zgwD5z4Cny63wR2TQ9G0x8XsV/uzyAciJxOhuQ71JospwbOvKUykO4dQ90DvvP2Aihgw1fF1lhGXU/6SfYXcYpxjI6B2UF8EO3Aa8ZazrEgBIkyYwAaXtmT5ZstT7cJStoJ/QPO26A6Sf0/WeUls/5AOYhQxmvsPmMGZSZT/QAPcGuvEJEBXkx/q54yJPCuenRA86IcHV5DrFHi+Nrr5YuUbHSfSuF5lpe1nOg8aUf6D+6iqwJI/UFJdqe8Y86Ek6J8Y7rICuWkNQOUfHY97HpPQdtBClJv51U6kXq41kJudbUfUffe/ADpnA9ianV2lf5cJ8t2IAkBMAGUH+TkhFVvHfwXPokfbxjF7vlvWRCrFPzy/9AN+gPeFuh85B74q41bmnvnVyhLMIin/aGI5Qjx8MiK77nyCPbnnn5Gw8ckecC4zkLYRjL0wf2Ie2iZO+O6WvwVJjUiSG/EM0K/GeMwBMYu/eCYjdBs3Dj7LHRE+WhVlLoC5pxJDbXd4dlBbBbdygxsGCzeD9E7+iz6D3eoNgL9Po1I9sW3tysFfPter42c2RDvVkpoofUlfGET8abzqF9QM6265UnqmePvyEKAhiPZSLqeH/R/xhj7H1++TXZ/5kEMglkEsgkcAVI4AUd9K4AeWVVzCSQSSCTwEtdAjbhZZIBUPF6JUA1xgMANSbBFWf2gYecOBzVzIyJCQAdoBATFSYoTDyYIAMiMCEGOFtOVBjIbuB+B/RUAtDifiMsmEwDkDAZYnLP5IbVjOTJLAZQh98Be4zQoKzmfcG5NLBvz7PypFekcc5mRkZ4UA7Lj9+oI59TSuz3wapJJv+sRjbiwVbIpp9lRAJAj4F2THy5BzmlPSTSQLR9pxzmccH9AJIWq97qYtfwv4XKAvjifz7TcrBrjfjhEzKKuu51nvjhB/VJqBBAKyamtD2/oQvIXmBfpx2Q/2W/QvO7Fr/qFZJwcLhUm/5g656plpcfOty+uqXQUGfkdeFVouHVQuVITGs7egBTHXBegCUTdPqk7anSK0NWNuL5AtDIwcSeNqP9AVG4/wLCYm0lu/hV7N0h4A1bALGALr1XQPhNfX5tqCyCQmq4MJqbKWxOjj3mtAt/po2153clxxrj4YLW/bdep9BK1wu8vNZ3YlZlAuago/SR/6HESmHTcwAe6gBZiA52Vu63P7wEXND/6B8k68foN3r6TF9UPzjRPvvoT079wU2vmv9G4R8mvnPjA+N3/YdTxc0AeD2P1859ee/tsw99uuWVPr2xfWZbLiFUVYItoi0AlO1ZEIMA4/QRAz8Ju3OvEqA/AAv9luvwBLO2oI07q7PPK8AffSxiHwGdA1QG3PrBlcq47PwSWQHxg/dA0WtNH23telwhoGang02JvAzQ2Uf0+zfDJEdZKBM2hr4PmIScucZWuE/qO+QLgD1ALp4s6b6PrLGFPJt78NToyFyJduJz6fpuaCjn5HS1NbltZEY3twW8aR+LZEFcwXQxCrXy3ttxTDHPG4G7uxZ7SRDFh08J6664bvRKJ2z927e/rGOvpXuB5MSz0Rc8id6bkocRFx1vE+Sh+o5r/4rbFB4rV1D4srzb6kjJVTgzQphtzJ+cG8ufrom0oN0gljhogymldYeBSpUFPTznqXjOngKEI0f6NiQCMsTeQgbwLAgN9BJdR8eQvXlhpLK98CvgeeogX2tHA60hlmh3dA6gEfBx+UFoJsg2xjmejX6wmppE6DnG+xUP9eeTRW1CveXEzPiN3zy0VWTFWLne7GzAzbEKWXGxrM3T6qIyWMeP9GNkzLhG3TBYgNK0De2BvvNeYl5D2Jw0YdfrUei6eV/8tb7fvfwi6eNf6tyvNKL+P1F4sgX1SfQDu2eenDyjqTGhJ0nV46FG5NpYQb9DxygH7c37G2M57WkhNJHlNB4aeg79PTsuLgEjZ5EhY5XcB7WhvMJC4QmAl0W+3B/7uQJtmT62qKe9LGjlt2gfh0/nEvcxeVk8rguwqeickXO8D5IYGyDLludDnn2yFG/U58m+kcbw4umh/WHb74whSvZubYtluB6iHJ1g7KHPGiHC+/lyT8zzCi2C4qS8Ix6ZntowomoW5G1R0z4ch7QBOOMD96KvjIXYEMYq+ss7unWi7Id0X14bd49tnJx5enpq7GvaD2PIdQvKT4b3nA2y9/7Os+Mo6KvNnb45DFqbkO2yAxv//yohoymly/79c7kAsv8zCWQSyCSQSeA5CWSERaYNmQQyCWQSuLIkwAS3pT0JWtrPAtARsIIJAau3WAUMaTDjNPZd6xz/H/c7V/0MRAUrzJhYMUFiUgSJYfs5MMFPH1xj5wzQN4CfiQ8TIPufyQ6TGcB3JodMtAF6mBzxXCaOTMQhASxf7mHsYrLHxMwmcJxPT+Bs1ZoRBTbJs/8pC4n/qRMTKib8tjLWVo6x4p0JGpMoI1EolxEC1N3y5ju/MVm0/KmP7TFh5AjXpQ+buFpe1I9nmpzI00gKAzZ4pnm3cJ+dZ4JoJEZ6Ykv9KD9t/Cnn9IdYmYlnDW0PwAbYCvDHCmPKlrAdQQAAIABJREFUi24AEJJXW7riSGcuy0N1c53W8cJMbsgb1SLwICqFU609k5VkKKjGA5HC6aCDveMwv7ASoY0eUKLd2DfmF5QMMDR9BkAhsQqY1Za3K0FYAMjRXgBwS0vHX8jidQFS9AtyEZn8stKEAGJFxtAmCiI2FUarpH0U8m6p6tQLTlgN/YP1uBAPhPVTIiwAzgCbqRuAOSvmCTmB7tmqduvbFjZuqS4C+9NHmpw7D+zTZr6uPCxqB0avnn1s+ObSk0PXbxVw+Dvyvvj1DrifxJW2V5i0zLRR90feNH3/R79t/mt7c0l4XEGUntQ19AmL6U+7YBdsZTykkRGw2Dprs+fCPZ3LvFPG5STFMqCZS7At9LdfU+K5rJheIiTOq3WPf1Sjx0+0d/zyyfb2bz/R2nFtLRrSjtblk9q3AYTrKf2OV4iFa0JWgE4PKaE72F/qCfoN2YUtpP9DnqBPkGMGcmILANcZI/jOylvqT/ulyZmlUuIdoX+S93/w4fY1O8fmozhuaA+LovZqLmh/i2f73fiZeuKX9rW8O9uOO9mO3NZC5A4cTcq773P7TwlkdQWyWlujC5QPvfmMEiQyYO3SIW+ozl4ep9rbnelgYntTzTjoL4jMaToK9dbZa0VbRTuPVV/9+G1DD8ZDOQVPd2JCQJGmlNYEjq2wTwVyw25DriMzQvXRRwGO0XPa9nVKgOOAl4x7tD1gJnKFxGM8on8thddK1y/9fZlHVGf1vw7ahfEE4ozvkEgQbOTba98O7qGMENf0wbtWel6P8//gJs6DxWb7Y2HOu/b0ptEd/bVGoezKF8qJX6PfeK55VNKfV/Km6PXI9Ar0ixVpXn17KQyT9j/m2kPqv7xP3Kf+/mf6xFYhX5MtIDKyxyuCcJhWRvMe5XMtBILZAPa4op8g9w9QAIgzDkLiyVPvhxUm79Pqj8gZEBhZdBje7nMOSZ9oG3RvNZLEZMGz0TH6HiSyhf5CFrwv8W5AfrYXSEff9Jyzqf5keWWf50sA2fIOSj8FmF8i7Vr1iqNQUCI+Pc/vz7f0hT5mx3bCIC2eHqwoJNK0QitpvU+8X2MjxB/vW8uP9MKVC35UmKXFOPSe0N4YvgiQH++WAwKCMZL2xR7yzoztZWxF59FF3ukhLSkb45a9O6zUzlv0nDvmTgz3+bnY2Xrdqc3iELD9lA87hI5BrOJRge23RQL0nZyUfWMc+rM6WciXgzE/H87niuGW/rH6A0Ejv00eF3dLLh0vOHlSzCdRNNeqLi7GQXBzD7KCyyD5sIHYetrhAkZjpYpk5zMJZBLIJJBJ4PKTQEZYXH5tmtUok0AmgUwCK0pAoHMigNZAQGLQAlqzASeTbYAVJjxMFCacfT/rirAAALUQToArTIpsEsREgnNMiLjGVotxHjAAcoL7uQdgizGHTybS5lUBMMGzAc1sAk75mNDzHCZegOw2aQT0YXJ/LgbNuecDPpgnhdUtvWptuWcFz2MyZyEu+E7+TAb5zr0AdkzIyN/iVxuIaESMfloKXUPZjTShDIAg/E89jUhJkyo2WSUvruV+rrVrkNVyIqQD/vFQHXY/eXOtTUptAk0ZqB8gFDKkbpy7T4mVxD/azQuwmzYCZOPZkFN/r/RRCAp0BZ3pPvOy/ijGwck/a78n/Eb71j0KZnKk4LarApxaApsAu+gX6MGLeSBn+p7ooQ6AjdfBzynZ6v70CukpnQdUQG8AQwkZAXD1vMJBraNSlJG+jl6hNxbKrUNsKaHDQphdsOOFBb+/ujWYoYzUhXA42AhIC8A7ykp9yctWNKOjawELLyiygchiHa2fkD/5djy7BGIeySfBqVLUFH7ivlEBPm4UWI1t+fDfbv7e2YP9u+f/8NGf4HrKRF9AntQHG0B/ox7mBbLUJyAkIEnSnxeTZ4/QW+TVFuCMfGjvH1CCHsQmIifK0ivOOfr4oCpTGM+fvmo4N/eFajRUlYfFovT3jNpgoxJt0imzAZWSE7YVfcG+AW7xfM6RH3UFmNqpBLhO+1Iu5AKhyypy7A3XQXDQrlNK2PsVV293iQvuCT/y+UOtVjt0gzBaPBO7Z54J8sOnQ+eZdiw75XploYAzKjGEFuQpbcF9dlCO+5XQQezxu5V+iB8BiVXvDjGBN4VCY3XO5b1zG5Frw3FH+1k4ktFfyfti8N657z1yy8BD943nz3xde1sA+llIptTjzn29SLg0frb2QWaQOMgHgI5xjzGQfAEtsfMAx5ADjDcQGsi2qgaiX2xRQ9gYC9FA/4rXATCbZx5jJAQM4zleHa/vludieztwHSl90A8ZN3rpHvrzx7E2I1kYGagq3Xf1vuPeQKWR98OIdgHgRK+oA2MpsoGYuVMJwpWDOpI3cljt+JwugMjjIGzTq7AxoZf7+ZZXvK7u9101XRh/XOd2iaRYHAoXD6h/n3pk5JWPb2sca19X3XtkIKyapwt5UDbqh71Jj8X222rlsd/JAx3FTuCxMaUyTKJr2jtGG4H0oXMvnw3G78h5wUI7KtKfkQ9ALJ5Z1B950Hb0R8hEIy7WUgYjOCgDwHL6XQg9oG78xrsUzwXgXvN+GmspwOV2jTZ3jm+98x7sC/qJR87SHkXac8FpVufkYdF5FUyTFUtiCAN/WCRDqW+4OeLlIvo/xGr64J2LvrBimDORFUcbi6WpJ/7x5ZsbC6XbZeOxD7ZnG++/5tWM3mGDLVQf9hnbYmXDNkG88O6AjpHQOfJADzrhqpT/aNjKObPHRpzBjZXBwYnKpjjy6tqAG30ib+yW6Q9jJu8nHLuk7xt03YT224hE1oxq8+2XD4zV2MC7T8TN7pkjo4V2XdtwqMclYdhqVuePtWoV7ECvAzKRMvI8FmU8r3eBFfLOTmcSyCSQSSCTwEtQAhlh8RJstKzImQQyCWQSuBQJCIDuAED6jARIA2IAbjDxAbwCaMD1m8nJtc6hX37E2f3rrHZi4sPE2ogC/mdizaSLyT+TGiZAnGOSw3VMPCx+LxMP8wgwMoHVWlxv4VUAjQBhWYFNHtwDSMbki8RED/CYscuIBfPmMFLAxjX7nzIYeaCvS0AFABtAvoVJoRzmOs/EkP8BnQAtmfQDRC2foBpoaWQMYAByMO8KymJkAuUwEoL7AGnJ08BQymZysXztf5u0cW163OY6nm3eHkbgANBSDg5AMwALJt9MAHPOvS4TcMAp5A4YDkBJHoQV4HME3eBm05VuXpflR5eQaSSfbXhfrr++KWeB5qi7ELTlWSGygjbqrIhdB3B4qXKiHwFCAID9ByXrT4QdQZfpHwAGrOqlz7Di37xA/qnIJXSSZCB+R126FQcMSQghxf//x7mT2BoAcQBQVvxTP1slir4a8PZCl5/8kOd+rb4+3HRL5aZXom+wivMT2qC5cqY4MacUPT14XfiXW3+g5/NXiy9vXhQXhHzqCmSNHzybPvoxpcNKDyphkyEx6PcARegjABh9F3Dn8wp/NPrN6m2nHqu85qTA+DPSWe4x7xDsaTutu93wM3URF5BwyGaymxcgKsAy7QGwyljAyl4ITvQMWwy4TNtxQGgAumJfpnmGPCncLjnRveTCjx98/e7O+KNrw33aSWLezwsv874Yuv6cIgkNSggAbowN6PSnVE5A+zRwRZnxRsBeIxfCor1W6c4o8XWhN7ytONV58Fw4hofFvEicg624nFeorA2S0T55AZ3eW7t59Inqt12l6x9ls/K19u8e3hXYaQA2SF9kxzgJ4cJ3fjNvCQBpZMwnuk/9OoSA6qytfJM+daBbVVEFrnKtT3B9mrC5UKDPnUFG3MeYhmywG/RJxhrGMcZiGxculo/91osow5toSonxBLKFPk19Wjf/4rMQd9xD/0ZfsFWUA53GJrBA4s+V3tw9x3iKft6lhCcjesW4RPv/Xvca9ICy0zdoZ+r2hPrytkpusLSYG6rV/P6pT098Z/OR4VsGh8LK6Vvnv/6PIiQP/93mt5efGbh2rJobdPvDamVj+2z1bac/Ffxf+38jWdZPL9Xm2GIBZP13Sj8nPcSzokOQPVm7VSTZ4LuG/bm/kB7Sf0nYb2TC2Et9GWN4z0Jm5vlxnqfcRWwQ5beQgpA5U0q8l9HetA86xLsOR0H621qrrnfvuRI/VgTKBbk7rdq84/m+kyv1t+ReeN57ociG4tlD43s2v+xM5OeilpuL8Q18u9JruoJcCmHXQ7CLMoZ/eebQ+AGl12lPiLfpGt7x6G+0IX0a/eGgr2GT6WPYQ/oh73uUnYVA3IdOYpvok7zPGknCe3/aa5Tfx0Q6OMef2jIssuIakQ5Pje2YG1BoKMgO9BJ7Rb8mKdqbOyjGcDFs59r1ufJAZbo/SRLvTGmwNaTwVdqA2xvXvTOlwebjTQWZVdHfqtIM+rn8K/183g1bF3Q7TvBOc79Sh8jt1qVb3ewjk0AmgUwCmQSuRAlkhMWV2OpZnTMJZBLIJPCcBFhN/9PdyQwAFoAGEyAmulucw++fEWFxr77fo2SrjW11q606BkibVDKPAgAaJkQ24Qb8ZzICSMPB2MO9JK6zyZiF0QBgoRxcbyuvmTBBVtgqWD4Be7ifvElGTthMiPy5j3LYymmbiHIOIAWAh0kez+K7eYEY2ANoZxM7W13NvUY+UB8DaiE6yMPCXtk1XG/lMzIDcIvVlFwP+MjzmViaDNPkhMnKSBwrB88mX+4xsoLfkB2TV+rMJBfwk5ABgEOAJLZ6mzamrKxkpo7Il8koOnElHv6vFt/v/m77Z5JTiigy7wwjG3SsQwgI6DHvl+e96fYahUpbQn7RLyDpzItol74DVnCOctFfbbPXcB1x0NdYjPMvW2VTbi5eC/Bn/Y9PswudB11qyLFVSIVO/+tubAwQwoE9w/NgrYDw85LbOm/CPkwp0U8BwigbmwOjC7Q5wC5tzu+QB8cer912+r65t79WgPwtWu3KbwCg9H+IZ8DK84BPK4/q3ZA8iOvPNeiVrbLHbkCWme2kDNgma19sIrYTe2ShbZa8KyAteMZKxIUB/u9/zm7bPkWUmXwInwKwhj1ihXMb0sJxfsyKTjm4h3Ly+3alT8il5/UHGte399VvvGFH6dC7tW9A44naq77Q59XHt5cOPS1vmq9VwpFXV6Khh2aCTSdEXOBZeL0SMljohuVZSVb27OWfBghCmEwqISv6LosAWPGOnbcxBDtLAhxk3AK45LqyMhlTpb6iz29TjJXtfUnYaot4CRR7xlEYH12z5CGzUkG65zvgtRI6jny4l+fR39AX2hhPAwOwV8lu6Wc1V0cnOBjv0T/GFNrLxjfCn1n/rom8SHtQoctcO6WEPaV90WX+R88oK+UE8EfXGDv5//eVAGUpN/JMRFJU7tt49+k/337PhsX8sF+KGo+LbFyo+IN7tNl6/W+2fv+2wM2PB14eDyN0+9RCbujqE6WtpceGbn76N655b+D80VKYsaUKXuKXWGHYTuh5f6QyvK2VlK/R/8nBxnXuQjgaiLgoixhTwKD4gLx/0AlIR8YX3hloC2RDfQG2Ce+H1xzttKLXT4/y2jsGYzhjFW1vYLrZkyAjK1Zv6a6XBfL7w277fH9Klo5CGskZzHfyYXii2D94St/RUWwJR6E2X36LPCQeKva3IX7RZfqKHYw72K/l5GHHE1GeDmePP7V5rHJmsKjvOcJM6YCE7nWQN8TxDUq8F9CXsP/YIJ7BeyWJ/zthmVIHz8eOY4fQyc6hcjun9k+MDC1Utmj/jIaIC/Lk4P3xd5VuVJmGorY/IGJiYfHs4Nl2rXBtoT/oV/in0Vwh2p4vt5P6XN/Trhs82zd8xp07vnkxiZwjYbvxymZtQXuBNDt7giw7mGfcrwQJjr72tMXLb8r+zySQSSCTQCaBy1sCGWFxebdvVrtMApkEMgmsJgEmCKz8ArwBEONg8sVEhpWidzufy3/EeVNgQAxkxWT3OvMgADAyEIlJkK3y5FqbNFtIJwP3yYIJO5O3q5VYXUnif4BMJvGAGvwP+JL2zmASjjcAk33KYKGamFiZZ4UB/kwCOccqYPPmID/qB0hiK2MplxEqlI3JEpN+QDny5zkW8oYy2XO4Nn1QZiMYKAPXkg/3M4H8mhKyYPUjq8j4jfJQX0J32JEmROwcMjb5peXIdyMfKDflBJziOyvvmPzxvL3Oo9/FxJSwAQbEM6FGNvxPWb6udH+qHFfMVwHmwV9/Kpg7HU988Wwy3lJoEWQKOAcAFL3YhMAyQdPWtCOJAz0GsGO1sRFWRuaZd8IltdUjR8E0LjhMl+0HIwcvuPCVV9EdVz6WERJrITcuqT69bu6CdfbsFVfRvuAPXl+G2A2AVmwA9hM7AbjLqllAKQhd6nC4Efc1H5z/TleruRcEluLVhj0jBIit3u88GZJgBUIH/QJMw1ZD3GJbsU/m/cIzCeljJBnX0tCshEV+Bop3wCVIChEW2BFXn/Fq3hZdsZhOkS/loL8B1hohjSzSJG33ts7zuY7xJhRAfO+x5q5t++uv6Bd58wl5UdQXwrFG4Be3+q0dwdlg87H5cGyj9rEgnBC2Frtuq5QZ82yMW6tuci95EO7JPLG4F8CZ8lI22sFCNGFnAaXpyxaahzwgAhhD86rQsKeY8PI52VFywqN1x9+6O663+pOoJhRvxZBbCGQZoRgrxJiNfejLV5QeUAL4XxNZIRk9Jhv4jD4PiAz6mNZMz0t21YLXsv1l2nrmirJKkRexyIs08A5Rz7gIuYaeIaeHlNBFC1+EXCyMocXpb8iLwvk3t/zh+Ini1puafgldH4xcv/MeorLmVFbakfrxSR7oE7oLWAsR9ldKT3U3oF53/78IaRt/z+f+lBCCjZH89IMFt3X1UG6hJZmFo7npGXk9HTnV3tZUBK0vREnn3YWy4YVjiz7oc/QhSDr0GVtPX2T8oQ7rOYy0svcwZE2y/9eT15V8Lfo4pfR/d2X3Bn3uQSBR0HKai3OEOdqVL5VPemIs5GmxJKsk8jbW5vpGtXk1NhlCgP5NfyRP2p82Qh/twAackHdGXWGUhkRUPCNvh7WESrP7IUDRHXuPRWd4jtkldIv80iQJ/Y73Pd5Z8XrqhEhVGZzGQtnpH633aTPuokiLZxXyiXzQH+YJui4ZiQK/1qyWZjwv2T60uTIWNnOF+ny5XBpohSI55nOFIA4ayZD2s9hQGijtO3s4jKIgcKJ2S8+IlM7rfrxrMZawuAZ7lZEVKeXIvmYSyCSQSeBKlkBGWFzJrZ/VPZNAJoErXgICEesK1cLMgfAiTKoAAQAKAGEAjopOHPYLrv2G45dYxdWZsOlgYmThnwD/AQQsnAGTNIAHwBzO2cTbiI3loDsTJiZ1PJdJFPkCrDNxAURjrDKPB55NfqxahfBYHiLJwiilwysxeWNCxGSNZ1Mu8uc75SMPABVbBWoTfANrjTxYHrIpTSBQLg6rm5EaRmxQN6631aN/oe8fUfrP3XJxvXlukI95TvDdAGnLe3loKH63iSi/AQhxLZNRwBtk+JgWn+admU9ZnHo+aWMmocgCUBAdiNEJq8yV9Amoe0+jo3tTSuivrVRG99YLGq1bdGvwEHhR2yVNOIi8QH86wHP308Ke8LkEJuietYK765bHS/GGHuGCrBppgtHOLZPdj6XP049t5TrfIQiwT8jfgMf4i/NvSbQfAzYMIBzykb4O8MO9EB3Y0xWBWQgclRkgDVuLtwJhaQhTg/5DdFoIkZ36bh4/t+s7K8Sxi+aZlm4us138fgHIjp4vkxPXYx8Bq3gOdgug1vZOwGZin3oB9nav89DCt08/XLlrl0D1LfsbN1aLbuNQKy6KBNEI5yTfHPAXD00Hm5sCtSFsbSyCgEFmPJe6Uo4Llv72IHxoT+rHfcgdIpp8KCsEPG1E2RhDAQ4BoC00FOf5bh59czqxoAwZA8ux6/Y3He+7807ySYWJqs24hV0jSf34j3/oydquqI4ditZCBEEmiLRAD5Adz2LMoZ0nlX5IqQNQ2sF+HyT9DbRB9KPagwFvhyNTzWueOFC/vnq8PZlUwuG2CIt23g2Sg99985r7fnd/l/TjKBeERZoQtfEUkic9tnbaePi7UMfO2I2MkRVjHsQEutqvslMf8uVdhHcD7CV9A72hHzDOEU6P+x9WmyKX9ewRslT+XpuuP1yZ8zfmTw4q7NjMluLRb1SikfKAv3DiquLBs0Pt+SfOBFuOqoyUi/pRmclumQCS0XVC70DasYDEQvhIdzv6c1GyioL1GD+MuMjA36WWW/sXeVlE2ssCHcIL6kNK2Ax7/xVp0XaCZtWJ47GrxVbYohkeUBWRMbB4ZvA1m/ZMH9JG1DPaeBsbgX5iW9BZ7MyBbnt3iF95LSwGzXyiDbbnFGYJr6/vXHtpOzYe3bJ3VAgwFhxB9tHPKB/9hD6D7qFn6BzvgNiuzylByHQ8cuLIdeaOD39FIZ2S4S2LR4p97VtcL6HfvEE986Q22d4rT4xdjUppi7ws8ro+UnioZGi86vnF8NkoTObCZstrVpJS2Ao3NBbOfk+rmlwVh1JJiB02tHjuwAazH9LfKGH7zQNyHdXPLs0kkEkgk0AmgctVAhlhcbm2bFavTAKZBDIJrF0CABPvUWI1LQAUkx8AASb7TIBuco7+1mecyV9isjWpxGSLiQ0TYSZhTLgBwA3EMSLDYu9bLFp+T4PtaRAPMIw8CZlBvqyKZDUXZWF1Vxp0A9wnbz457Hm2CtdmQ3ymQQxAG8oCoEFi8ka5eR6JZ3TCxHST5ZcOuWS/W3gsG0fTAIt5Z1h+lJG6MfllVeXHlVg5zcplACSek963w0CctBdH+hzPNBLDykPe5Ml5W60J8PisEhPV2Dn1ZxAZrCym3ky+AXAABi2eOgAOunClH8gQwMgm/4CE616N+89ZiN3wVhSxE+Yq7T0issKICiPuDChHT+i/Rr7Fuha5xBlxcc6LYdlhZI+RkfRLsy1ceq5fdnVrhc24uQ57Mi/w2V2+or300Q+Yjpq3G8Am/Z7CAERh3y6qu12vE4uBD2kJkIadwv6ThxHYgOymC9gQbDRgHnZ16RldLwv+z8nLwuxvsgrIzvWAa1wPGc3/PJdPvEuefe/BD0zp8wIyQefM9lImxoooiAq5utMPSDgtb4unK9HwMa1yRxaUF1KGEE7s5cMz+J86U18Lg3UBGJ9qX7PFlNXCpfCJneATcBDywjxl8BxkDxz6y9KYpz7D7yF7ClAO7Vsxpx83qMJjgeM1FcIqGUzCDUNJOJxL4j4/SY62XK9STOIK3ivUezXioqsvoXSHeuLFAPGFnCAvAMYJG/ZKhSn6nnZcqEtOroidV55qb58T8N4+3pqcP9rcrTBaI7XFcGRAgDsrwRmjN6ncFnYQ77NVyQuRFr2OdH/g904+XVmn8zSbhFx532C8A/gFdGWfCwgJ+gC6SOgaI+yp66QSK9BtfIRwo3/Q7rN6VnMt5bfCr9TPFfqpLI+nMXlXeGeCrY8149ImfT+xvTj1NZE/exfD0aPyVAH0NUKRkH70oV1Kb1ICRAZcpn6QarQx7zbmXWfedlaU7PNFlkCXtED3eE/DfqSORG5ddae5MJP3Riee9fMFCIIlj19tll2oL5RHB/PRnIB/9BVdZQzl3Yv3UHQW2xDIq2Hf6f0bv65Nr69eOD3EnhAsZlmTJ1S3QDYOWPnQf+wo/Z3+gGcVOk9/QJ+wPfauSD/CzkOS/IJlIPLkHWcPj+0VWfHopmvOPDy0sfpG9apAxEohaOY2yQNkVJ/FZqXUatcL8/0j9W2NarFy9vHNewc2TPfH0cL2di3e3Vh0t7SqoePLByoOLyArCH3250oQuniBIZeMYDtPz7J/MglkEsgkcGVLICMsruz2z2qfSSCTQCYBYsc/ojWoPypRsNKJCRXAtYXnAGybco7//oSz871FBe7lGiZCHEyKWEHKWMJ37gMYYEIOIQDgwOSI37mH77aq08AIJk1Mtux6wAQmT3htAI7ZyrXlEzKbeBl4zzOZhDEpBJyx/QfMq4IJI2CBlZvJINdTXpuImleIhXEywsAAsfSKc86lyQrytboYkWJEhxE51AcC4dZuWSAQACsog21e3i3iUjktT5MXZSbfNLHCOYAPwDK+G3iDrLn/tJbMVZ29P8X/U0q0BZNC5ARAQt60q48upAtwJX3vsUL1siIprC0FuKE75k1EP0FnqoCpM/N1v9Zo+77v+bXYzc0FSf9gzhsr+m77ZNsRIOeMnAmcmQHfWdxccBelRO3jzaTV3Rh5VdDyCtIn+jx92myO7T/BCl1sEUQhIDn9D8B61RXUabIiBZoic9qQ9sT+AnYaQYItNGJzLaI38Jjysc8An9gn6gHYi+3CZmEjKLMBrxd4HwlIjwWq80xbUX4eCNVrNXjX0+Ow7iG0CZvNAl4BaAHUQvZQv86q+B6VMZ3GhhMDHduMLNg7YN5JPABHVqFDzBiozViH7aVtaCfy7aww1mEeEj0e1RnruI6xBWKf50ASITNsM3aY9gUs7ACSSknKa6mTZzcEm7VPePvD8bQa4H8rHW277q2C+G4O5TVQTqL7j/rlnAiNES9KgpybtDbHLQv3tCZwr6s7gYgLSCHkSdn216P+tvZbmGpEfY+dbF+ViKwY9pzkzXtrt1x9Jtj8OoXUOiPignBj2+V50adPCCHaArKdukJwHUGm6wH9ewnVzi0jBJA1bYsOUmd0EtmTeE/gvIXWAZDlWs5TT3SBRRiQHICyyJo2RyfNa86Ipudru9Ll2y3vnjsDpzCpzbVr2pa4JtJp40K4AWKsHiY59ANvCQOLeSbPZ3U59WKFO9dQTvob9eU9iGuGuh4hPdt7Fe883Z4dlyABe7/6Y+XBgo+lvSAIa9SszI26vh/1j26adz1vHAcCERTV8lAzVNikYnW278jwpgp6iR5yoLPoL++dfysCYFKg/5FDX9s5KK+FnUnkvkfn1kNWkGd6wUy6qvT1tyrRZ7Hf6B+EaxR5AAAgAElEQVQ23Yhk6oYNs/cAe9/s5KHyv7wyPfDLW687xYIibGVDzhHH5k8Nf+7UvonXae+Ka+RdkXh+UgkaOTmGRfmoHd8Yh8GovCuuqZz1nOqMWI6myAp5bXQPxg3eUR9QYuyArMCzwvbaSZe/813E0QXnshOZBDIJZBLIJHBlSCAjLK6Mds5qmUkgk0AmgdUk8FFdQJgIACIAACZTTJSZXL3caU8fcebv/Yoz+h23dTNigsTkmd+Z9DDxAOQhsV8CE27GGCZmRlwwAbd9JsjGVqrynWsAlZjI4G0AaGV7WBiQliYArD5McngO4IQBG+TLs+x6ACm8CSgvIJN5U3BfGrw1oM9WRtsz0oSFnbPyG3iWrgv5Wx58mgcH5WEiyoo3wmsBUiArVtwBpED+8Dv3pPM1MMVIEn63MlG3KSXzFDEyA3nQJrTNGefMh1i9xmR7UonJKZNG7gGAAuBBFuhAdlzGEhDohe4APHRi9peS2Cs4cfvVfzkV7Ht2Oon9fF+lGg+FhfzwsbabG/S183guVpgav7i34WzeUnRzs6E7fbzlTMdO0lA8dudUOzk7lHPq/R+fr9eiTv+30DfnSfJSQbUeQKb1A/oCfdcIO55rfXypDJf6/HWoBX0QOwNItFMJgMtCweG5ABkM6A9JSP8HPDqh+tneABd91LJ6IAPuB8g3+wVw++nuOWRCm6znQJ604ZQSNhnbxOpb8sWeYFsAhM2+rkSKmL3qhMfrEhg9gWERHJTPgFpAcAvpA2DL85EfcuS5vQgL5AC5TTgmyo5dZBNcG5sgECykGmUgH+wegDb3ARYzVvE86sw4uNKzqDd9CCAae43syYN7kBEyp22nH7rNs7IaqW8hCDlvRE/nGl0byuuCjeEPi5y4W4Xc1HD9vqNe+bo+J/ryN7Vx9CG/r/HmYNrCVrFPSAcFXM3Tgms4umGimo9Xb2srlJg/G457Z4MtcZJ4B+UhMC5vgKMlv75wpr3lnfIOGKhGg3vkmVLSfiCMy8gVbxe8UyCTsCHo898qQb6tiTyxsqzx0wgB5M2zAF2RM+1K36IvAfJTPtrL3iMoH9fQnpTrTiU8bsyLAZ2k75Hvo10Sa0Vy7yK2w8Z0dBMS5waROoDET7mJbKTrvUpEz5RkCCDL+L78GRbe7R/0G/fZewCLCngH4uA9CC+SzyrxvnOBnC+yR003i+zjEiXA+yQk3/1KP5DOKw7bTrs6P54rlJ4tDoyUXc+pD26sfkmExc2FssJGtXLY+sllz7f3wyfkTfHQM5/fM9BcLP2E9r54w/nRktZc6iU2YNkd6BD9lAPdM2LWdI3z9CvIFIgzbC/v350D8iVXUKynxN2kJB41YauO3bl8uH9k8+K4vEIWKjN9dc8LN7SbQ+Jr2sVGJdx25oC/LZf3nIZ6YdSGrCDM1FLJ0Ge8KpAnBDihCzuhSkVMPF/icM2Cyi7MJJBJIJNAJoGXlgQywuKl1V5ZaTMJZBLIJPCiSEAr6x+QlwVgD5NuA/aZTLMCeEJBYyJn6jddZ+jOpx2/zKQfgIZJPxMfAwothAcgEIAd5w1MBOxIb8htHhJM0G3lJMA9AAJADiuR+W5khU1k0mA+z7OVvkzkbfUy5eN5Nik0bwtWHFt5kKN5UNiKTf43zwVb8QwgYd4dBpByr5UjHf4pfZ19N2LBVnRSLjZlBYDgHCvemCySD7JIkxHpVXPplW8AMZST9gGo+YNu3Vk5ByhD25AXXhd5p3nimPPke3gevwGs0Ka0DdcA4lHWr6EDVCw7LmsJoDf0A/poYyAJj18VN/I3uo0NR2cTX9BYn1+IB8+G/tWe504MF9wBuVVFCqxd0xLrsdmmF9a0nvKGPnfq3jmn5Lnunnbs4BV1VOGpjyrqQ0OfgMO2ufCLIUwj5ejX1Mc8ugCP+W42AdDY+uk/lbcMz8OeAJbTv7FR2CNAoU8oQeQS7gVQiHdwACTAVQhFwhUZadEr9FEvWfI8+jKAj4UuMbKSNlgJyFpLu5gXFmXCZpjnWGcfBaXVyojMuY76Uz7GitUAKa4HlKYtsU+MR8iMVcDIE1nhtZAGba2OlPGwErYOUvgLSlNKyNjICrws2LeDPKgPiXtgTADjIZL5jbKyqni5R4cRIwaWI2PkTf78Zl5rEBc2vlBu22PICAuea7HaeVZHpnhdyNOCZ35KgqLu24USbvETbzFw3elZN7/nH/MbZ8Zz7eidrZNr3dRc2Tx3QFoolBhlNRKNceM7lIb21m/a77kR4aia/X51TptIj3lOxD4gJ3w33J8keQB5SG7AcwB/yvgOpY9LpvS388KDpZ/7PAlD5GRhKgHxeUdBrsgOQhDZ3tc9R1sgf9Mzu+5enaNN/4USOovdeEv3WupCW0KCQHysN+wScqQcvKvQ5vy/KBnJDGqVfNI5xxgPMGvvMmmx8J1yMo6zYIC+gq4D4lIX2gY9RK7W13sSwsszzf5/YSQAiK69LIyopY2w3YRY6hyJGIag2XBq0yd3Jk7yuWK5pM2z41kRFm55uLF9IBdjW+gbRkDR3ngVnBQJMChPhdPzJ4ffpL0rIEBf6MPICvJlTOK9FjtJfRinrG+h9/SF8zyZIU/ajYIjz49pbbz9FW3A/e3ay2Jiw/b5HxYZc+zs4f7jYUsh7JqtUqumXXfiYCBsL463q5gz1wkhK2J5ZcROWckOwl3RZyFI6BMdW5l5UbzQTZ/ll0kgk0AmgctDAhlhcXm0Y1aLTAKZBDIJvBAS+LwyAez5htKrlSzMEsCG78x+9jqn9uisM3R7J4RMd8Jjk2ieDyBuoAGrqJikA9Scu/85MIHZDBMVJlMGLgKycy+TKMYmA3jIPw26GYhvgBnAFICBhX6yFYoG2jNNAlCyUFWAFWnSgnIb8GYrggGMAEJspTTX2HPTpIWtkk17gnAtRxpQs0kgMmBSyGaKRvQA+hjpka6nkS1MMA1Y43mUFfkw6QRg+aQSE2gL40W5kQl50h5PObOfhBChPWkz27fDyBnammtp++y4jCXQ9a5AdzZrM989io3/zE3Roi9F27ng5av1OOibiNr5QS8/Ouy1dxdz3nDZdfPTbXewEiWnhn13/nTb8wq+f9XZthcvhF6gpdnJjrJTKXtuVRlVDjeS9rQC8OsZ9EmzE2sBqtcqefoC9gTbAagNuMfKZQBjdBtQiHPYFWISAfrRh47ZKuoXKnRNjwLTZ812YWcMzAaMxP7QHzmPjcI+0W9ZAY6cLNQNcdDp21Pdcl8A8PeIoU/9qO+blF6uBGHE/9gBs1urEQW9Nu2limmQdb0r6I1kpb0sFn8PsV1wipXykBaAgsgMm0m9sHFGcNtqdSsjnzyD+wDmqD8ErBFI1XS7d0NDASICEJM393AwZtEm1h4QDORrdeH52FMIP+5jvMIjAzsOYY49ZpVyII8J0wcIQtof26wekwxrmTJ1Ylyir9BegHYdsB1PC5EWeLTkJfyrBXxvqLk+Y0YnPv5Zr3D8rFOovL/vGsJbdYvdc9Plpd/sS9cG0IcoD3tY8Em/ARgv6Fk5eQO01dD98rg4Ju+Ab2pV9bD2XlBfcs/od/O6hDxAhw3wRw549RjQfsGzVzvRQ68pJ/0cudJH6NskyC90G4IPnUAXeFcxID9NTqK/6ALgKP2K1fGQh1xLe9ieAvwGMUZeFxwr7FthYzREF7pwvxJ9EZlQPogwdOMIz0vvE9TjEZBo1JH6oG+0Cx5Ak0rI9sHuecpr70+9ipqdexEk0CUt0BnIL3Tl7Uo/a49KhMYH7YZTOfVssd1fnNl2QzQ/PrkwqNBQW+SRwCIRbAr6hT53iGqRAU80K8Xy3InhMI482h3doe0fUsIbdkoJXcJ+vFAHOo+3MR5RjDX0MWwQfZl+wfPt3VQEhKuwUN5M2MrlWvXChAgYxgCFiHMKfj4slQYW6kEjGYja4US7UR3D24R9PeIw0sCh7nFu1EFn7fiivmBbjShZKcTfC1XfLJ9MApkEMglkEniJSyAjLF7iDZgVP5NAJoFMAi+UBLTCfp+8LJhg4+nApH9KCbAAIIUJTcU58EtF5+bPTCtILxMvpiNMsm0VM8AH96VJBAAhJkS22pZ8uI5JEfnym3kXAPwzGQRw5BryT4cdsRW+RiwwgWTlISAT4CBlMsLDvDsMsOI6wEIOe6YRCUyeAMkAK7ie1ZhMFE0OBkwY+EddKL+FvEqDW7aq1oiNtKcFk0Xu4zlMGi3evO1fAfrENRY+xDxY+N3AQuTNxJdVl1NKTDoB6SAkOJ/2Lpl1Wse+7Oz7BYBMQB7b3wMZ4X1xXVcWJ2j7jmSy43KWAPpU0DrIUEo63HD83U/7g8VbosU92tA3mAmdgYG4PRj6/liUi7fMLDYGBvNe3Snmc1rhPR4l3vyYG0We2I4Zx7vq2lK072zbiV7R7+VPtJ3tBxrOdQoRBTgPEGyrztE19NT2SrkU+dKXAL8BLQEIsSUALxb+DQKA87aCFPKV/kLfoRzouN/dZHc174B1lbMLBNNPKRPlu6lbVmwDpCDn6YfmTYZ9snJN6jv9nj4qJxVFv9cK+51R49izfnlpQ+MeoKmVEbsEYG4eZEYm0948Y1WyYl2VXePF3c23eT71sjZai1cAbYMOYa8BbhmTbMNyAC7OnxuPnhsj+J3Eb1yDXQTwxR7SBr1kQNnQH2T3lBJEhJFLP9j9zTYhN7IXm419hiymbLQ59tf22GAcaol00MdSiEKuA+AvxnGnGLT9LhEXDREXGsOSfn0yZlJO6lr719vc8I+Oq5udA70ZS6iXefvxLPMyYrxZU/umdJRxkkT/IB8AUsYj6s93gMtRAY7aU6MDOqqMPmMF4yF15fe7uuWyfgR5yBhEuyB36nIpXk2Uy0hJnktbW8hJfoMwsr04OuEoVyEE2Nyc9wTCV5EX7x60KavaGQvJj3y+1P1ci0wt7BukGnqBzqHn5pnEOwXtii6v1d7YOwbvJOgZ+kA7QVhg2ygnbTSldCny1e3ZsR4JdDfgxrYgf/rjEmHRyUcMRBxFd7TqjWvPHgo/sPX65NCI3mRdv9NutCv3sX8ZulJvLJQ/c+ChXa3F04N7RAzwvkl7Yhve0C0X/ezFONArypQ+eC6Jd2r0trOHhshKeY/kx+LYLasGDe1p8SlPUe7CdnKT5wcHS4PtA1G78YY49sYgKqIwcOJgRVX/T8oS20A/w64xTq+XBH8x5JHlmUkgk0AmgUwC/4wlkBEW/4wbJytaJoFMApkEvgUS+JCe+VNKrAoEnLAY3Uxwvu7M3b/TqT/tO/03tBzPBwQ0MJ3JO4B5B4xRAhAAcAAMmFQCTOM3gAyANO7jevJgks/vjEk8DxAJIIFJnhEARjKYFwKzIgBIrgeU4nx6fwojDGz2RN48P00o6N/OwfMBWAEJAKJs1Wtn1amSkTIGJliYCltBTp2437xJmITZyjXziEiv0gV0QD62lwQTOMCTtEu+haaiHuRv5acM5I+8ADkBQe9XYiLIZBiZnotTHIdTzqkP3u5EVeqArJgIE56C32lbns9zafPsuAIk0J9EZe1ZcUQb63r6XpKSAVRep5j59WLOrSrO9Hi10d7pFOJNThgX22G4WIqEVmhT0ULJG+pTkGqdO9SIo7k78s78F9q5Dc9U3cHtZReSryXlHFTneZk6GeAiIDA6Pan0DwIM0fmeQODycDErrGimX0IGvK6r+4CLFtoHUJMV+fQ3QELbaBeQEsCYVdCAMVw3r/xZCd5Zkf0CeVzQT+lXALaQvIA+1JfVtfQxCEZsHmApQA22Be8WbBf9UG2RnJRwjueSZEvOSV6vxa33asNl1/nofPWuYKZyV31/snyvAtUDu8AzsM/mycD/HXKK+il9Kw9rcwPbzS5frEyUmfuwxdhGIzwIB0Tbpold7Dl2F7lDdBOejPsZQ3gWMuD+Cw4A7q7XDSH6aJ9/qYSeQDBxH+0I0YDt/LISukwIJPYjoHz8jw4ha55FWCH0DftMu3Q8IkRMbFSBJoVnDgjUHNd3z02SEf1fTNxELk4u4J3GnqQm4oL6xm8dc5siLPC84LkGXqPrkCs7lYyo67mnwYW17ZxhrAVUR45GZKGLjNH0C2wBZUFejA/IgcPCu1EO01/CQKHDjJ0GdgKsIy/0mXBctqfECsVZ8bT1JfozCYDXVqjTlxgPaWvKiszXRI5025v3Gu4xjx28QjgIBYadQL/QOwsJ2auQlI++TNkYfy2kI8QFgDb5oO+UD91Zr4eZvU+8UffyfkO7o0sQsoQXop0+oIQsvtX9u5d8LttzXdKCsY3+96dKP7K8skmUjJ054P3kU5/N/8dbv6/dVxpMtsvLIi8Lgc1AJ44pFNTZmSMbvlmb67ta3hV4a9CvsdsrHfQlnmsbd78YMsYmoPfoGu+zbZVzY7NarCycGtg3NLGQU6irTY6f5GSn+oOWM3LgS/F7FA5qIgpD7VXR6oTH0oENw9bY8YC+YKfpV9izjo1TynT3xWjFLM9MApkEMglcZhLICIvLrEGz6mQSyCSQSeBSJKCV9s/KywLAARDiDiUmzEw+ACoIm9HvnP5Q3dn160xuAFQAEyy0ApN0JmWAhuQBEMTKTP5n0s7vnGdSRAJgY2Jkq435zu/kyT0GBBkBAFBgifwAj5jcE/8dIBNghQkdgJYRIJTbyAx9XQrtYeQDkyeez8payg74RTkBHSiDERz8bhsWkp+5zXOdeVtwDfcDYnGfufJTRuqAnJCZbfbJfciW87aC1iZxNnEElLC8qBfnqRPlBjShjIAwAEXkQ36QEjmnfeqkc/g3kAcTYfLnPp5tbUq5+mlzfWbH5S8BdCsRWTE5HIe7xpJ2s+rmXhW43s6iGzZLscBxJ/FzYdSfz7n9+bxfduNYDhlRKxfFcSHMt9040CbdXt8t/X4h57kbhovxka80Yv+ZmtvYWnB933F3HW4m8/OBs11Ke3dXT+kH6N79XX29YGVwetPYi4RfMRIQ8AagH11/ixIkHX2OvgG4ByhkoW54z+X5gLQAveg8iT6AfaLPXgycXFUrUivXARLp/4CpAKzYIwBhWz379/oOoEnfncg78bAEDsmz20ucPSUn3ivSAuD9ulISBVrd/gqlG9QAh57IDd1HubXJcrSMtMAWQYACRHMv+VM/wC3k860GhSz0HG2HnNdaHq6jHthLvlMX5AhIzv8Q2ng/YLuQu5FZ2DvzJuMedGNFwLi7nwXtBBhPuJK30jZKEA+scMb+vlLp25TQMdoW3fprJewxQD8EBiA4BF2zGwqK+qILW+VUMSnPit0KELXL9dw+WfNAIWTCUC5LAvjG3Jy/QSuZVU53n+d1SIvc9qIz/z9v8OZ/9MkYMgGbzfiGrbd66msHDEeXOsTARTxwuNbCK1F2+oJ5+5Ef47qFJqSP8ExCKLG637wJyQPd4kC3/pcSfQ+5IF9+g/RBjuRP21ifXI8nAPpMHugzes13kpEBkCi8J5A3urHe/RzQQeqGbnAvYz6kA7pFftgK2u1iZAu/402CDqIr9DuIDu7B/lBf6k9Yr7V6VujSpYN3BfIy7x8jNXnPoZ3oA8iHTYsz4DctuRf5u/ay4Am0D+D7Xykxjnx3+rFg9kHTHTzyaO7dihQ1cO1d4WJ5OGn4+WTGz2kzds/ZJI8E9ZdwkJBQIgV434XsW37wHPqWhRBMkwDrrSn5mMeuhWiyd2DyQo/oG4ydPHdI5MSc3pwLUSs4ffir7nxtpnzw6tvbp4KmE1dn3VHV7/b5k63RsK2sz98p3MqJ7f1NJcZCxlkjoDOvivW2XnZ9JoFMApkErmAJZITFFdz4WdUzCWQSyCSwggR+Ued/RwlABvABMJwJDxPzhrP4kOs0D0875d2b5WUBoMN5JuZM3j+sBLjApJoJC9/xtGCyZMAFoATgAPdZyCQAFMAUQCrAIiZTgAeA8lzPYdfy3VYP8wlIReI711Bmm4CRr4WOArSnHPxvYB6fBmgxkbLVYQADeC0wmeS7Pd/KYitL+R/QA1CBUB2c5zt5kQAsAR9sxTPltP0x0gRM9xFLhIw9h7woE/cgY2QKkISsAXQA51gJjNxoC8iLa+VVcb/z5LvPOtEChBEHE2sr8yF9BwxB3rR1dlwhElBM+qTteACUr624uaGG6+frbm561GnGpTi+OnHdAd+J+5JWUHLyIisE3il+faxe1Wi2wiASiiECwxVZ0ac/xVE/ar21FB477HnT4yNlbzp0q1+ruGc+MZ3ovqUNk+kHkIsAoUaOrRXEtFXylAUd7pAuSvRxQFzOs4IToBCbYn0RUIY+R38DjLTV4YAmXAPg2CFVBfTSn2yVdk9AfZUNg7E52Cn6IfYC2weQjR27Vwl7w/MBgwBbk6uj2vG2621QG2wdcqJntRfIiYEk2jyRBMlJr+DKw6Kv4CTlipO7rp2414YKznHI73+66frkgT2wA/mY9xV9GntGvbhuxQ2QU/e/2F+RJ+1POS8KVCHjZaC7geWA6AC0yBC7hzwhE2hzyAb2YqDOJIAx7DY23TbbXk3XsKu0P0Qv5WW1fWcltBJAPJ4XnLNQY5QH/WN1PqQ+90N+MV5ydHQojGIv58uRCQ+LJCnIi0nbxsRFbcxbUS+qirEQN+GMuJHbGeO0yb3GL1efTkE/+ON5p/aqQbf1jUpCPdEp6g5hYuSDkdnmfdh9/Hkf/IbsIXXQT/6nnNgAiBbKjTyRHf/TP6gn8luJ6GEcQc6fVWJsp1z0Tfo4nkvIDu8DriNvnrdWooryMY6ix3zy/oC+kxf91kI7IpN163eXoKKtIZfw1MLTgvak3tgTnoeMP6+EbqUPkyVjMgAzMkVn8MpBxtgZygUhgq1bTe+WZX/ev9T5q0qM1YSX4x2MsR+Zv0vpXykh90e65y/lWRcrR/ZbbwnQPhCc2F7a+ufSl4Hfx6Fz17HHc870lO8Mbow/KqLiieq0257YEyfaYDvXqrXjKAjOuH7OFtj0epIt5qHPXwphYe/LZiv4TBMWnTEsjkJsioyQPx4Fzemw3dJ45bablea1+78UDz37SKkviZMb2EBbNkxeFeRyQdeGSGX+gGwgMdFjrmzKQyXT06xHZRLIJJBJIJPAuiSQERbrEld2cSaBTAKZBC5/CWjFfVteFkzGfkAJQAJQAwDu3OSpebzohDMtpyFIsny1J9KCyRQJAIHJPJMeVhxayCMDD21lF5MWxh/AdvuNCRPgBp+cAwRiJgTYTxlspa5NsgAIAHr43Tw4mBRZaCV+Y2UXoD73c3CveVRwP/9zD98hR4x0oQ6AIwBWAC8AF+TD9ZSDctr9gB+suLSVofxOHYwcIF/zlrAypydt6fpQRgvVQVkAjriX8kNEmIwBh3gm8qMslAHg9lxorDj8rHP0t+9QwJ5Pds9RRwP/qBPADJPfv6SteWh2XJ4SSAHA6ORQ5LgTAsMrSnUp3pZSEi94TryoVfwbE9/J6dyQVnz6npZ8CzQNdVPYDsIhL+e1BKorSlHiBZFTLoVxO1f0trba0ZlyyZ2/od9dSNr1Zzf09xenWi77MNiKY/QNIoFQJpNK2AhAe/rXeUfayyL1A30GXYc0RP8B8OgTgK/YF/ImmQcHICdgKvvEQMhhA2xVPKAvq6m5H/vA/eQDwAqoQqz5nqD6CmUDYKd85MNz6YOUkfwmu8/lfwAtbCdx9gN5SXCPJ7KiFeXzMwU3ZnPlZNotbC0m8ehoHCy0Em+HPC78Pi/Oz3jsIZJM1hN3uzxivvSOD+9/6tXhfLPraUF5kSf9mXoiB9oau7PeUDS65QU/sG+0eZp4XutDuNfCqDAeYYuRI3Km3uTLJ7bZPP6QN6SRPZPxIU3wXPDsbkgw9jgAOGQFv3l1AF5DjDBWURZsMMD2nUrYWvQLcM5IZPMgQf5eFInnc90RpX4F/4Lrk2dFZ4wZCMNY/Yv+5vo4L+U8r6wHFKMkmVZYtlPycBocyzt92sui/dN7E4go6m0eNHxnPGZlN543rLTvpbfIArmbNyD6j2woH3Wy/T0YMwnVwnWdUDBKqwGL/E69P9EtB2UDwEdOgPiA7PRZrqNs6OVqpIWNobQzhBD9irYmbw7akv/RiTWFgered95Hl7SgrSFPaWO8IbBXeNJQd0hOSLAHU8/p9NlumSAKkBMeFoylphvomRGj6N9q9e1VPDtnuo/ssGe0NWXD/lEWZPs2JchWysKzL+V5FytL9ltvCaCP6MiUEjbonenLwPG1B7VTm1UsqFn/+/XbbTo3V5n2TqulRvyCu314S1LO+x1PpeUHfRJ9Y+w7L1v9Y++YtDdjFn0cm2DvuSu1F3qTJj2wRbawRmGqkr6w3SzH2j08X+5/SmTFeLtWcYNmrRDH0W5tpL27SY2X1g/14io6RCCkHeXiExvRIS4zsmKlZsnOZxLIJJBJIJPAxSSQERaZfmQSyCSQSSCTQC8JfFQnmcADgrG61UJ6RI5fzjutE+NObrjsxJonJ8XQ8X2b/Lxe1wIWAggwkQJsAFRnMmVhnphoMeEGUGd1oxEHFoec3wAkOABV+N1WhHHOJuYWbgEgxrwnABuY0PF8ABTKwrMpC5N628zbiAIAEIiBSSVWMTKpAyBiZRigCxNB8k57h5CHhb6iDIylTDABCTlvIZtYcWmeEQBFNuYiy+WHlcfqah4nAB9M/qxOU/p+lxLgBbIDaKGNqNu4dn30ncrXb3EO/grlubtbHyalPBv50pbkByhHG2fHlSOBpC+J5gWUn1h0c1ODSdgvb4vjYheOKfRT2YvjlkISNfM5rQuXvgnA6JdyK4qNm+T8XC7vu/TJkkLbxIVCrq00KiBjoB1GjcH+QqneCOItRad596gb/fnJ5Cn1UgMgDXyjP7EaGUAToPUCsqxHWBv6LfpN6BnyAwChjxEjH7AQQgRSAuAOOIVrrK9yLwANgB8gM0QftgDbALBCPyUv7nmDEivMAaU5t1bwD4CSOpE3IDK2i/Kw0v3TXAgAACAASURBVByw2+wS/djIik64oLFcMuZ74aiA651atVodctq50HOvkqfLhob2B6q5/o7tbru62QkOz7q5TWfc/ESQeNv25wc/OO0VnhHxEb7/HECKbZxSwhYgD+pj9nat9dAtL/zR3XjbQOsL9uBYwxON8KC9sGnoELLGPuLdwLkvdT9v7coCQBl5oCPm9bCGR3XaHHuOHHkG9hVPHOw953iWeRcAqDO+EAoKYC5c2gvl6KKB2wPqRJvVf7aJ6AtE7/fJ62JIBEVZ5/pcx50RKShvCsdLXIXmS7RzTJLs1rWhVi9HnryWXjnY0UXGT8Ykxifqjf2HaMOu094A7unDiHG8BzggWbiPaznIE88fdBJPC4B79J7nrIWssGfxfMaSv1PCm4Vyoe8Wjo28aXvG0APq2wDrKxEhZitoO+RNWVkoQP+l7wIIM8ZRTsp9SUS72gqCCjtkHqLYGMrHuwBeDBCbPBeijOfRZ6kX6Y1KjO30dcZ87kG+9Hn0ZKp7jz7WfpgX1zIbSD0hxYyAYx8L2ptn8B3PH3TyGd1nizwueOgqHmJrL2R2ZVoC6DI6Q7v/JyXGm/PCQ3FxygEBcuwqvBM44ij+qvq+xiBZ/0RjV5LU5V6FnrMXBEx4Rb4O1+mfeX2i+0YI2iKbuq57VDZkRNdskfFq6DvjAX1GZUmkNy7PRDd74T1ap5AEyjsQmbo/Ctvzrcr8HSIodjrz0/uioPUyuYCodBTY1udcVAE+rl8h63l3xi7SL7Aptggn055MApkEMglkEsgksG4JZITFukWW3ZBJIJNAJoHLXwJaed+QlwVxur9PCaAb8IDJcehUHw+cxsFjTtzY6eQ2DDh+ThMS3za8BtRkQs3kbVIJEIgJkwEhABq2YhWA43NKAIfMiAgpAfDYAfSUAFaYfPE/v3OkAThmUuYZQf6AdEzsyY8yA/JMKQFGcp7JHNcxgbKQUEz2AVtYucj9XAO5QD0AogBQzMODZ3M99TFPDc4xaeUenkvdDNwwksGAJv3UOXrVxeplxAzlBJzlOTyftgCguz31bORDGSk/9XtUobpc54nvo+yAuazspvyUB3kQU5tJL2DQx2hjK1D2eUVIQAHy/UmREpsarjc2mDgN/T84k+Q3SiEXFIKoIsBjTAroa6V3v2iLJImcIHIVpyiK8onnjzTbkQgMZ7DWSDY7bjyn2BEb85671ff92bGR/JBi9Td3lZ3wt1/mnXjfwXhmNugAjeg0+kffANCjv5hX0sVWv9NPICxfq0QIFvoB+g4Q8g9dvbaQM4TuWb7K3MLIAFoDXvMs+gLgJH2LfgzZAMmJvaKvAFACtpDvRY+udwXANn0NLzTqSV4QF5SF/m9eZecA7Q8+3AkrUy7liwKLhgVc71IooMlc3mvk46Qs5Gqi4Hn9bW1vWo/j5kLib23GycRmL346ceIgH0ezIpw2BYX82aejgTl5yLhNVztgnAOzkQurvgGIkZOFYvqWkhZdOZj3wWpi7fU75ac9ppSwdcgYwpV60n60LcQ0bcv4QVvS5lyzIoi7QkHME418/rErR3QYe0z+jCnYeYBuiAB0efkz0Fs2phWhRzw1RxtsJ2NxHI8LmiScWqGQz21QaKhZ7WOh1cuJr53s1exeIEJjoFzM6XluVfdMK4857YnR/u5H1fDCDpUvgCAkCmWAaDBPIVthb6uyIcsAtCkLvzFOTilB7tMXGTu4hgMSwMI2ragrKwDq1B05Iw/awLwOKBdys36P/JAp/W55P6XMtCVtSx8kjCFjFKQMdoLfICP5TjlfEG8C1aepPgy5CInPuEhdkCt14Byf6Bp9G6ICkgL7ZSDslL5DalEe3o+QA2CteTa9EP0OfaRf017IB9tCmZEv55CRLRahDJCzF5BCK3mI6drsuDQJIGtsG23Cfg3IHz0ljNxFjzgM/t38icNO38h4mC/1J36htEEtpzUAQVN9f4OIgjM5rQNI4igXhUHFzxdanueLz47aGnfVlxJfO+FsD1r101wbh+1jxYFRRXPy2eBbhEh0FPshEmSHIswN6tM8lZbKxcM0DsXNyuwdjcVZbW0V6j5IikS2Ia2+F6gyZB+EKDaQMZMD4pL3aOwAungpNn818WW/ZxLIJJBJIJPAFSKBjLC4Qho6q2YmgUwCmQTWKwEB2l8WacFKUibEAG+20nDAmfu8YL/3RE44m3RCQoUDx5xciUk/oCIAIyAIkzmABoALAA0jHpiAM/lmYgOAwm+A6fzPb4CAPG9SiZkSCZDD7rfZkxEhjGWABgAfgPVcx/8PKeHxAeDBNYAllNHAUspnJAT15B7OcR2rJwEHuJ6DvCkn+QBIAFpwL6t7WcVGeQE1IEIoK9dzcI5yki/l4tO+dy/pfJCXES1MegEkmPCRKA+y4Tv5ImPAKgAU6sJEdMFpHF1wprTmunnSCBdWuJ7bd+RcMhDvado2/fDs+xUhgZKi5l+rsENajem+WphGYVvcPKlVngtaZXlSvhRbFAsqUKyasgCLvjBM8sW8Py1tXhCoMSQFzWnD7kTAqgLaOF67LYS9lCsW8t64gJGzuZzXp5Wi9IuWVobHf3+LV7/94XhK/wOaAuZNKtF3ACXp9/yGTq+06tqINvoFq4whLQygpR+gw/S1XmSFNaj1N/oLtoX+8p1K2CT6Jf2OPk3/oP9TNrw5iA3//7P3JmCWHVedZ9zlrblW1r4vkkqyFluW8W7ZxhvG0GAwYPja0/ABhoFpoBsYTw/jHjDtoT/gAxpoGmjbjMGmjZuhvbSNLW+SbEm25UWytZekUu1LVu7Ly7fde+f/e/lO6WXWy6qsqqxFVXG/L/K9vO/euBEnTkTc+P/jnMNY0hV0FABoICvjBjv7qQ9gNvW0WBv8D6CzwNd+f08+ryEzL5dBvZJXP3KTS6CtArQHZe2yXoGX8/pxvOSCCYHbg2MuKK7TBtt1QfNEU9vwH0qjV8jaopSVB78eNDPGNkBUxgfcUgH2UmYjfpe1NdaEdYE+bfxOZRXS9RGyxGidP81OcIJKozu4P7IYPrQnhBbjJXWn/QC6DRA/W7LCymaWFuQLGYJOMA8w/tO+WHsg16WA6azeSJrqV/w+JUJiVkzEqigKq7l8OKl2H6w1RADKvdrcXKMpwoq+NVHIh7PqXi2roCTNCnrAqjgOmE+qO4pBbayRUTfbZQ1YzbwAYUM5NSG35loj3NkYgHxwbcRcxv9YNKLzEBnMS1hHQM7NSO5L9UGTyek+kTfPZvMB7YD+Q5CYZY2RkpQVwgVQ0/oVfY97IAioK32Z/k55saahn7GDnbkLAr7reHEeFgS0EeQe4Ku5GuOTg7ECMhJZM+fS5vRp5EYZcSPHZgjaBFdiF6J8lANZUU7IMZ6BTOjzyApZs4kB4gT9+Hi7vO0q+I+VlIDcGnXLrtU+CsjN4MaYw7st755/fKZnJ/Wqq06Ni5BoDuUKamIGjcpMmV0BSaN+W6l/NcFtCCpRT+o1OQmMIrlsKoW5fFOBMMYrEyM765Wpa0VYHNNFm0U6HA7j3Cc0fx9Om7UXiQRZX+ofCuJ8qRYXy2XN0633UnEULdMPWVSURXi46vS4SAp1Y50TWWJWR0sVnzmeut6lZEQf1hXMx/zmrSrO1PD+dy8BLwEvAS+BZUvAExbLFpW/0EvAS8BL4KqUAMAdwD2gG4tlwI6iK6yfc3FP3iXTDddIq/LGrZ2IRRZDgBQAEAAY7DbErZQtYlp+3JUAJljwm993FniAA4BRLPjIg92fXEc+gO58N9t0awieB7gAyAO4yP9mkQCwASjDp+2sNlcilo+RHMyFgDtcDzAAwENe5u8XQMYWYTwb0Ip7ACMBCtixTd4c5g6EZ5AHZeMAfDWQhms662LfzX0M4CMADuXjfgCyn1ZCDiTy3dH+HbAKAOhbCob+Nnf0b1lIGkFj91MvZEsdkS9t6o+rSwLoTKzAv3MiK56uuWCLfEEMXJtWn5JiPhUGaU+apXO1JGvk8xGWFiAXAwJZKw3tumwk6VDYDOQZKmwWC7H6QqDY3FmPFDkan54bGZ2uTg71Fcd7yvmJfK5En3MiKwxoM/dm9Cv6EuMJff7rbd0GiFtMDNBHbLxA/wFGzMUaIDW/AdhyXwtsPQNombRd0gDGfE4Jay76FvfTp8iDMgGG05/5n35yihVSm6xgvGIMYHyivuSBZRnn2fXMb/RFdt4uAIMLYoFkWRHKz1ZO7oFyuVyYk9eNIYViXSUio6x4FYDO+jlI1oTpbElsRiGINjfCeM1IEhcV+GKqoRAJs0FuVOyRgqC3QGBAVHOlQ3kYE6jr+QDRiPW8j45YG+ebF23FOAz5ZNZsAOOcNxd9Rl4vSTadRSGMuGC8R9c6ZWlkd7fssnwuaoqkQK8JqP6Evk9pZtgUBuEGgYmNSrWRCptch0mFXKvFxVxUEhEoewwZNaVZvpkmAzLRQM97RWhN3aZv355u1RNynPYlb3Nx9jp9N0Afspq+gmUAgDZlZ45CZnxHXyH/2FBAHvy/2OLhtCJaop+l6hfsqv6sEkQ5cyekIGWhP0AK0DbM6+amCz1nTNimdL0S8xW7tFue8tvlhCig/6Pjp/Sl0xZ0GT92xLP4si5Hl5ANfYf5mvLvUHqrEu8yn26Xk7HJXFUxZwNOt8Y8HV0JzmUU5eQlp5EvYxHvHFh+QLAQ+4DymdUPsuW9gd3vZ+Pa62yK569dQgIiM+ZEWnxTP6OzvMO9Wwm3YhDkXQ+RA65enXWQBnAJsqJQCDLNzCIpRGDLpk5OG3VOczHvytobFGOCIcO65GbFmxhNGw31L03V6K7y0r3Xudrcb9rDFES7lZ8sM1xxYLUTcaHLEpEieKKaV9fG3IyTBeV8LvP+q06xxGjnx7sj/dNIM/oDfRbdp4/y3bt/8j3ES8BLwEvAS2BFJeAJixUVp8/MS8BLwEvgypKAduI/IisLALyfVwL4ALj5lpu8b7UbfFXocutEWjT7XC7Iu/qkwvb2ndDqCPCIBRvXA0gALhrpwOIGYIOVEaAT1wGmA3Kw4GahzTX4kzdXTNwPSGA7IAFfSeRhO4h5DiCSgZksqngm9wJCAjCw6GPRD8jAec7xPPICrCQvEkCKuXTR15NBenkeCSCDxRkgDCAHz7RymBsWs7Agf7OwIC+uY+Fnv3POvpuFBwCP7coGdGQHJXlQZg7ASWQ0b8WSpaHb9563uL2/C1BBPVg8AgJxAL7wHflS7/fTpu3f/MfVI4EWeaCg24fVSSqCRQqNINw9mDWOrEvrSezkdiKUlYULtgdp0BR20tQNuSRJSo1mqg3/cgCVc9V8oFChmSuKwBgV2FKo1OpR0szSfDGOy8Vcuqq/hC6bJZFJF30HaGbsoM8DTtKHsMSy2BOLgT6zYACAZVygb5v1EqAiYOxJsmI5zdgRXJn+A6BN3oxt9CW+A6QayUkZIQMBA63fW5BtiA6upy8zpjAO0Dc7y8R9gKxmiXWyiNo8GwqE7purNbeEgXyPZ8FgkiY9ekii6MuTkqt20SaDwqz6FVuk2puTq6DMrRacXZKnqMnBODs6mWQvqLpwIB+4AzmXjkwL6dYDzLLMxiPkfjlYWCyneZZ7jbUFsmYNgz4x5hpQZkTCWQPHp7PuaOvIssr4wq396QMHp5qKUTErPmIqTbIZkRRz0qL8bLXRk4iNEIkRxdpGnctFjTwh1V1QbjSaDVlbKH5Fy5pJPmKColqvRZr/3KYgff9h5TEPFkI8MLdB/EFaQE6wMYCxH4sA5kLmDa5Fz81VEOfQR/QaUqClmydjbyyrdqe9CJmzy5+2Ye6GkCTYMCA6ZeI8/Z5ND1gmoZuQJliBUBfeBZhPjaxkvKBf8T5hfXZBu56HZcXJimBd0iZbAGCZrxkDkBVy5aA8zKGUkfJh+cEcynsLfZw6c/0CSypuXInynSzos8Qc4x+WoxZbi3Iyjj6sxLjEeb7TNy45YdlR/qvhK/pD/zKLPdqBWGFY4dFOEOX2bjYvj3mrBpexR6DGMKGD2VdHXWSDq2okaf03P5TP8wytv2b9u6RciT/RsszQZDI3cUKECJ4IeWWct7AQ+YElx7zFxdIHVsT0vz9UQt8pPzdA4vFp804q0uasx93TPdj/5iXgJeAl4CXgJeAJC68DXgJeAl4CXgKnlYAA7i+ItCB+hfmZ3ulmH5129eGq67leru+zAVc7OuriwXXCPcsKwt2juBYAjoARtgMLgIXFHHmwExhSAMCEz1cosXuS8wBPLMQA3cw/sxEI5Dm/dnuWrOA75wAdyZ8D03TbgQsgCeDBYtGeDwhkwJdZUVi+tuva8jXwxKw5IA5YjFJOgBcDVYw8YfHGc5hf7R7yMgsLI146gURb5JmlBWAnIAjncf0AsEt+RvoAmrCrs+ya43U3uyfvDv4JwCmExeuVPtOWA/Kk3pQZkOurtGX7N/9xdUnAdCuVW6g5YSMEdV5zMCwdkYuowSDLqiIxZqWUjbpIClFqPdoBHsnqok9+9iPhHVUhKjVBHdVaI8W1RE0gS6XeaNZ6SrlaXzk3lmQuqYkSKeSjxbss0WOsewDSGEc4ANgA/MzN2WLEhL6D7uIGCnCTPsz96DHg4NkExl7Q0u1d1YCngLZ80p/4DuBLPzJXKz+s73e1/58UqMkzbfwyayfGKSMgd+g75abvAhZ387WfyWolFgnUJzML7ZRt9WnFOQ+Tej3oazbToixccLvVcg8U5sKysKsgSJqFQZdUGmG+FEXJdZUgqo02s2IziihrVG26qJG15AXpgmwBqa+o3a6LwF8jKczd0II2vgz+Eb+UyXYi7M3lgnIUBauFD5bzsas3FGhbSlJrNJIJuYaSX3odamztsBZhIVunRBaLgavoHpsXGPuZK+krgKHoGTprQCHn+I25ztwq8TnvKnC+v2CdtLOtF+hG9TzdQC0lYtrFgHLmuC8pMZ9jEQBZwe9YYWDxges16oLLLQ7mL8pKXSA49inhdgmAnjxPEodLPfxcz0sWWGBZv4ew4D2A/wFrkau5uGJupw4QRYC4lBH5Q/xcDHIAGfC8v1fC2uIHlXg/Is4G/R/CijGSMYj3FHsnOlfR+PvOXgK0EXMFpBa6S1/EVRfE3Efbn7Qb8xoHbbe2HTj71KdBZrTOnhsX0CIoklZwDNesYRw5/whIErOyWPRQ3MsxtjAf/rkSLtnQf8Yg7uZ/dN029bRc4y3hLuvU+vgzXgJeAl4CXgJeAmchAU9YnIWw/KVeAl4CXgJXqwQEdP+pSAvAD0gEAIaNbuKLRVe+od8V1gWK1KeNvjOyPc/LVQzguhZDUc7iJhjYbpYE5taIRT+gOoAfQKEB/IBQLPJYHAEcAGJwnQEWRi7Yblr+Z4FlRAQ7IdnhycE13MuiCsCTg3zMQsOa1PK2HWOdv5vLDAMAbQc59QLcMPKBe60OncRKpzUFeRh5YSQH11JHwEYAURaGlB/3H7h/QF48CzkBogBGbHKJfAlMfjVy+/7giGtMs0A2l1fsAGWBCbDBjjh2rj6tNvygVdZ/XnUSQMfQp++Xk4lMsRC2NIWDPxb1Tg9kjRPlJGlo1+WGLHDTUSoQLnSKu50JJ89mI7ET+JGQ7/1j1XqzpADRrpCLp4V37BPoPtJouEm5uJkWsdGcq9br2zYOJtplvhhdaQgQRA8hIOiHgH30i1crAeyYSwkaxkg99Jky0x8A5wx8A7ykv5wbgkOGBMBWf1KZsI64u/0MiFPGOMgVYkHQF9kdTh/C/z59zFzZ0b+wAgMEhmDEkgkAlj7Md/qpuYmhTq3juu2rAwHV8q2leCBCqev1RMYqWVmyZ4xSQNW01yX6QYC2ON857czvS5uJPAy5eiEKa3NEUVXfrmukkfegpjDt7TqlAM6tMY7xB+IFcJqd9RcDQD1ZN/9lgQRSuf1iHhtTex+R1cQuxaPIKyLunKwuCkqyoAniYj4ek+uvqjY8xyIoxvW9UWlkdfW9Zi4nolAza2u2eHaOsTgd6Be7tQEP0VP6BoA/Yz9gP32HHdD0M/obeo4ec196gcF1+hb6Z9aN9JvtShAXgOkWA4S5Despc/1mlkG8N1Bu+jz9kXFjJS1BWgLtctBfeRb9f58SGx+wWOB9AlIAAJffcPvDBgtkD/lj7yFL5bvS53ke7XmXEuMQJDAWNsgYN3ToAmMRpCmy9qTFSrfAmfOjDxipahtlIN/YPEIsGYgASDyu4731J9tZsuHE3Iue+Slnc0WL+DCSotWvmMt4f/2v7XKgL/YuSrkYNyAX0XEO+gfvoFei5d7ZSNJf6yXgJeAl4CVwESXgCYuLKGz/KC8BLwEvgee4BFi8/EcldkqOuJE79rjc+oZb92M9LjckYqGv4SpPh668TbbmpWkXrQY4YbEDqMdCzeJTAFAYkQBoCaDBwgmQw1w28TsJgAawgIUUwKWREvxv5AJitR3ktqAycB+wH/DfglgD/3RaO3SSBuTBM8yHLws0rrUghEZMMHcCrrAgpWw8ywL4UhYjKDhv5EZneW0xa6QI//Nc6ooMsNrADRS/Iw+exye/2Y70Q27uyZo79mERR3dj6cFiE3DX3EoBaLBQRvbI+y8omD+uWgmgQ/RHwGx0Y1yERW0miMNjYWFqZzLXEEg6LPB7Su6gZhRlQZv904pA1SQXRbMCOrYLNReFIUojzWrNZlLvLeWPiOUY01ZxBe1WXIssmNuzf6T5wy9R/+9+oI/s/geQoa9BAlAuvgME4uLMyETGA4A4+hD6CxAPQcAOYrNeOO/G7LC2IF4F/Z4+ZkGdzQUPu8GRG/0MEBiglTGFPg/RSh04zxhDObn+lNgXFHb3jjXZ4eNTNbmDkuFEJo8faS2Rw45m0gIeBYgGxVqzFbA5yeXiRiLDC+3SnxWpoc34mWJyNyeDJBjPh/HamVDb96OgNJkEgL7ICiKZ8jDmMu50WnGdt6x8BmclgUTtpvgvaU3trLjpbr/acJUslkRkSOGDYJ0IilwgskqERjkWNaH/e/kpitwxuWBLWm6kFMhCT+3sT3xHt9BV9JR5A50FXKRfQVIzD1ifgjzDSq/ltmgF3T+dSRg2d9N/2VWOL38Afw6IC+oF6M/c/xIli/XENfQ15j7qRh0vpqVQJ8hscVF452DsZM6H0CDANnJmzLqYZeuUOXKlfLTvK9sypd+jG+9ol+/z+jTXPa1d8J0Z+O8rL4ElrAxa75WKb0Eb2HuguU3l/RELnr9rtxVkhr0Lv7H925f1ybj+GiWIvNe1Pzn/pnaevPdBrHFgucjcau+h/6DvvFPSz7jf3pU5hw5DdPLdSG7Ib+YwdJ13X3RtsQWF16W2sP2Hl4CXgJeAl8CFlYAnLC6sfH3uXgJeAl4CV4wEtEP/mKws/lIV+g0lFlkVN/PgKjfwclxDyev9ZMHF5VlXGyu4wtrdrjEqQmM14IO5UGKhBMjHIo0FEsAFwBpzkQXNNhdNyI3FnZEVZm1hCz4WTPN7T+cPA/95Bq4RcJm0o50397CjDDCk8x4jDuwc/1M+OygXgIQBFZSNurR2Z7efaeVikWn5cM6sPmxhx/+2gLTv/G+LRwuYyzPYJQsxAYhJGQBHyJ86ADbvcdV917qn393nRj5J+djhzU5wdnwCqgJgcg75suj8S9quo17+69UnAXNV1nKnpODbrUDXDcVTGA4LjYkwHh5IGvIdkQ1q97cUPBjUhkylrJDIj7Z2++cVE1jYujuh33G0PysDjZx+bzQEugt0rU6m1aQdYHkp6QLY4CKDPsS4QBkA2unj5u4MkNLcQQESAuyYdQifAJgGYp58zvn4im/7sKefAPDR3+g3lAFSAuAHwoSYFpSVHdcW7waLDIuhQF/dpwRYtKS7KixPPvXNQwpZkY6r41eifNwbpWHdBcm4gO0cgLXcAuXUDmUXKKg5njwygc1Cr2OFPB9S4IOoqcjbUXLs0Sy3Xu69ktks2KLCRrpXAdVb45cB2exKX6ot/PkLKAHamTgWOZFNIv2m1T+eoC/Vasl6PNWLoCCEdqTGxf1XqL5USWTTFCnurkxvptWYw+IwJvSd8d3mEysx59BX5lD0FKJihxJEBQAk4CU77XE1w7yKPlYuIllh5bR5EquKTyixo/zH2uUFEKUeAO70ISwE+E5d+aR+3NfNrdoFbLmTWXeWnfmXedlIFLNculRkhRWScRRrD94dGKcYm5j7eV9hrOX371eiLhCq3tLiYmjOEs8QmZGKtLBf0R36JfMd+g9pwNiNnjHv0Kd5Z+M3I8xxT0ZcGDahMJ/T7ncpMT/RV5i77L2Td2D6G+cZC3gOn9uUmB8gMJl/0W1SK56Nkr2P8tkiKpT84SXgJeAl4CXgJXDJJOAJi0smev9gLwEvAS+B554EBHzfL9Ligyr59yn1u5nH1ruGCIqpB3OuvCsWsKYYFkI4qwdmXWn7ZtdkzRw97eI8i2kWZOwEZbEFuMInCzcWXOb3mhsA/0gsmADubRc2izkDC2znqS2ojLBgsY7rCxZqtgAEYLSYEjyv00WTkQZ8WuIZdo0tLNkByg5GFozsVON30EDzad+5E9asNszCopNk6Xye1YXFIotSsyYxn/rkTx4cLGgfkRuo9a7yaK+b+W4qsoLd3MiV6wB8WaCSJ+ctmPEdtFk7D/9xdUsA3YAogAiA0HpMirpxOCjkTwSFse1ublL7udfL5XVPM0sEmLqn0iy4VoB5UQ6hpmR9UUnS9CjRQcMsmBRRMVJvJieazeZMvR7Wa42m6erppGyBf9ldzQFZAThDUFL0n75Lf6G/0rfMTQx94kElgpiSx4oebR/2uHOin1Me+g/AkLmvM6ssygGYSj8GMOJgjAJcgkw0AmPJ8uVyYbNQiKcl63G50arXa4k8A2VTQabQ52nar532/Y1Glq/WmkUCdOtBg/IXVC3mYtDtSj0KJxtpNNFoBqvVoBP6XbyFO8x1iiMCEIUrm9lLAFCvaJtcAZnR39CHo2pX4o/CrAAAIABJREFUXKgFxL5N06CgMLrTjTRdI74iyInQEB8VEAMmjV1VxNRhWTBNQGKof5qlTvDVF4dBh6u11twhl2Z8cI1Z1FkMCPQAQJQ+ZVZ3l0qkzKHMcYDm/1MJ0NSsgBgzcP0EsQLBgssqK/elBkyZx0nIz8D+zg0IlwOYi9yIOcC4+Vol23HPGMWufIhWfjtCjI4L7ArsUunXc+a5iywwjBSzebMuQgPdp1Njbcg8yMFcAznJOyDtzdzJuzBzEu+4jAVmCWHvsMyrEO8233ItFopcb2NEK3+VyVyePmfk6AvqJeAl4CXgJXD1SMATFldPW/uaegl4CXgJrIgEBIB/RqQFYOL3ao/2YTdx35gbfHXRzR3c7vJrcy4nzyTNkZyr7K270m65kKkNuGD9kPaOWiBsFv+AFwDsABkAfxAZ5jsaUJXzWBqwwAIQtMWbkQH2yXkLcs3CjWsBcNhpyILNiBKu5zdzKWU7yTplYu5nLB9+I38WkDxjnxILR64DuDQ3FiwiLWC4uWJhEWi+fjvdWhlJYc+lXOQPMAqxYoEyWXiaeyiuedw1p/Ou+nTZjX0xc0+9C1ICogI5AkAD9HxBCVdSLFb5/U7aqrOC/vtVKQEjANBRdA1QBPBfJhXB09Ug2Dcc5luWQ9rxLTwc6wqhp0mQhJHTv0EqpLWs3xRo2x3TuVQuoyYEsE6mSXJMRMawyIq5M1hXmODpE5QBMA1QFd3+F0oQEy9Won8CqFBmykRZ2QlKf4OsAKxZDjFyLg1t4CTkA+OOkRfkRZwNnovbJXNrRT2wqABIor91jRux2MpBO+mb2mHfqNWbsyIsjgm0Xqcd+LE8PB0LsohxtTeMsin93lAA7qIMKxJJo1FvEuciqa4q5I/cVs72zlTT/QcbYXZLT/CYCIv6oarr1aAD+Gtj1LnIwN+zshKgPylORUSQ+jXqSwfVVgU5VgtlfRGL8MvLbqkeiK2S5YV4jfRYFMW1MFLQdZdN4ylKxekk2BeUrk200T/QP/qTgZtm1Wig/wUH189gzZMJMKd/QJ4zZ1E+dJ36MddjKWC7uqnjBS/v4mY+U/kXXX/Jytcmqaw4lAO5YpXCOxRxTdihzzsH4xefRmLcoXsnPZG5sh18JXNrExqL3xF5RKd1jBGASz5axAd9infCkxtplHem80ZSXHT9XUk5+by8BLwEvAS8BK4eCXjC4uppa19TLwEvAS+BFZOAgPBPiLQAGPsJN/rpm9yaN29zhc0DCufZcBN3pq60q+jCOC+yoiJri34XlbV4EiYf5dgJCtAOkYAVhLl9gczANB2XRoAugBkGtrDotsCcgIQszFmU8zu/GZnBd37boUScDQgKgEez4uA6AFDOWRwNuxfZdLqLYoHI/Sz8AFf3KQGksjvUrEGoC88hD57BsykTiUWn7cC2T9uxaQAUoI3F7DAXDpSLw4IKU9+HXXNm2NWeeZ479pGc2/8H7L57qxLEBH6LKQ/kzI+0ywy4+t/VRrgQ8IeXgIET9Bn0Df2BHDR3Y2PfjgeSt9TZlOtqQk3Z/Uz8ikkRFLpWbp/qSQ8RgKXp8gaVRdoRPqvPipKsBFIAs+UelIX8+UTnGUMoE/0KsgKdpi9hcQQRAAjLdfSzrj7jV9jtEf2WPkef4tnIDMGYlRd9HXCVvk69CWpLX60DHi9HCNOztSyfi1tkZD4OBDSGG+XQqVfEz6xcQYm0THtzcdSQn6BCLh/iMoi4IfIOldVyUZwr5IJCfy6be2tf9uiDc0E6lHPDw82gMq5gzfVmazxselByOS1xUa5pEQ6FfDSjoPVPyFoJK6YtIi7K6gA5KVsjC9NKHMelNMkiWdcck4JNidAa1zUW5JbPrEsg+1YF2m0NIcC/6C9ApR2XGzBp/cvIwZOWkivcjy9K416Kh3SREzKtq/0f0ufHlAjczFjJOwFEFu8vkBe8h8zpOsaqy00vLoUor9hnQk60K7egnTvOX7F19xXzEvAS8BLwEriyJOAJiyurPX1tvAS8BLwELpoEAMRFWgDoPe6e+JW3ud1/tk1ERdkVdxZcmK+6xkjiwgN5F5VCV9ufunjDlIs2AMgDqgFIXqOEaxrcQwHiY1mBn12APwLbstjC6sD8cPM7i3O7lwU4C3FICMBOiAgW6Jy3nankYb6nOc93ACCeQTk4x+5ELDIsiDYAKXnxSb7sYOUZuIrheYCqRjQAqkLAmOsq5lXuAYixneDd4maYiyrqZn7z2UXO7m6sLQAZKBfPjt3kPdvc8f9WdEc/BNhMkE1AUn7jWdSZ/5HtPynt92SFpOCPTgmYxQ86TT9iJy4IJ3oO8VaVhQR9q7XL+b0f/oY81qSz2hl+XBYABcBVRX3OCTsXjhpoR3hYl6VAQ2QF/aDZvne5EqcsPNti19AHsLCgn6D7lAlSA8KA8xYHx/rVcp9zrteZqw5AP8rJmEE9IQCJwQGJSVkZP+iDRlAu63lvv31X+on7D9RmZuvjcS4+JjnvkcXKNZHiFYigOCLCqCaLlr5qtVFV0OZSHLWe3yzkotl8IXdU7rn2FUI30pcPp24vBFNPVoPKzb2ufnNvUP/PLx3otjt3WeXyF10QCbTAZFIkqxoF2YbokgsvBbfX/FaIo6q4qP3qVD1ZEPYq4P0RkRVcD2GGnpGYW87Yrm0g+7IFojuA9k4w9bIt7wXRhgubKXpD7C7GpmuVeIe4S+l5SuYyiPGUMQ2d8oeXgJeAl4CXgJeAl4CXwGUtAU9YXNbN4wvnJeAl4CVw2UvAglvf4/b86vXuxr+5xsVDspqoV11hU78sLoouLsjK4mjgilHJ1ct5l+/HpQrgPAts/C+/XQlQjp2hxIdgMc3OZcAa/ocsYPENaGggvQGeFhcDEJTvEBB82s5Ns9KAaAAYJU8W7xANBNEFgGRxb8G2yYdrDUjh2RAU+LOHGJi3eJjf8c1BfjwLSxHmVJJZUlieBjaZZYWVjbwAEFpBUdtlALCFtEA2uL+ZdUc+OOue/q2cqx+F2OG67e1y2+5JrjP3UORNm/jjKpdAh+sQsyLaJ5GYX32sBl6mRL8CRMW66eQhAiIRaZHWG4rAPa+L5BFgXSH1TrRbnPP0lfQsyQp7hrln49n0E/oAz6F/8z8xLe5RgqTgObg64rcFVgwXYVe2kTjmGo4+17krvDOWwLI17odfsq3xl596ZCyuJ66nlKsV8znYn765WmOmRRTF0XpZVPRKzhP95TxWFmWB2uO5WO6f4vyEduJPyQqjXo7D7KWih18Kbazj5w5SvIWHduYvu1z+wpWTQDvwtgVmbvVBEX6M+Y8pMX/0xnFYVUyLY5ow1mtySGV9wfUAzha/6VIFnV45QficLqYEILqwsGR85T3H/ue9gvcc3rv2aG7Y7+NZXMxm8c/yEvAS8BLwEvAS8BI4Fwl4wuJcpObv8RLwEvAS8BJoSUA7+SdkZfERff0VpYp79J33uev/7I2C7CtuYChw0SoF4q4VXX7djEsb8tZ9WOD/nEiN1YflMgqw/7VK7PAG0MG3NUQCwCTg/HolAnES64LFN8gbrmO4ht9YlAPusBubXdgcgJ0QBnyaOyiLX8H/WCjwifUCC3uCUu5uP9+sMTp3fUJWAO5i6cF3XFlZzAjAXspkVhXtIpwENA3shKgwt1Gt3dJKfOKygV3cgLZcC9rI/xAzYy5tFt2xv7nO7XnXCZdMAnKx4xyygvofVgKEsKCq5j//I7SJFWQlPuV7XRuCA33I8/rCWCKL69v5OAN1O11uGZGzoFjKeyWK6fNYWgImd3SLvgQoSn+BJHhGqdOFTGcu3Me1RhLQUOgt51tA/TLjVixVMnSXvvhlJcqGlRMWVvRtdgXTNyEu9ymh3604GxeqoZfpw76r26dzIU6GBkppPhdNyooCw5Xv9PbltlSq9fXVelotFKLjPUGwTdYtxYG+4kit1sw302w6H8dH8oVwuJTPT8hRFOOnEUeXOkDxhWqW53S+bdICnbXYRrQZOgQ5xzxSU+MbKWhWUIDMjOHLtq54TgvJF34lJYAu8Y5j71BYY35RiXcHxk9cSPLewftDZ1yElSyDz8tLwEvAS8BLwEvAS8BLYEUk4FGCFRGjz8RLwEvAS+C5JQGBzycDeQowPqO7iTPVTqQFYP5vKeVcPPg8t/nnmm7w9vUu7L1OwaKbrvfGXjf7xEEXNCNXvDaUV++mizflXL4XN0YkrC4stgRADVYGkAEsqnHFhAUB1hMGclJ+doUTBBewjt8MUDWXT+zOtuPkrmidAKCFhAAYgoCAcIA0gADoPMw1DIt/nsd1PJ/ycC8EgxEWFoC704rC8kK+9vzO/M0nvwUX5jfAhhOuPnyNG7tjxD3yrwjqC5CLHCBrzGoD9zTUj12T7D6nzr8nsoK8VuRoExSLyRZ7Ps8AYOsEsTtdfXTW9yTA3SEHu3bxe0gnqdH6DbJkRSp0lWWyyMKCnbXEPSGwtfm5/7S+Q4TNLTf+wvmIcFGwWMsKIJc+hLXHRqV727oOsQKwRtvfqcSYcCksLM6nyme89wN3PB71lvO53nJhIArdZsW32Fxtpj3FXDQn64ptcg21Rr+Pqg9Ua9XGdC4XPT7QX5woErE5Dhl/IJ1oz4bA8WXF0DhjofwFKyqBBw7i/WneQkkJfTeCm3kEIo6xmzmQsZXvzC18MubTtkvGr1jRgvrMntMSWDS+ok8Qvm9W4t3M3l14Z8KlJlaYUz6WxXO6yX3hvQS8BLwEvAS8BK54CXgLiyu+iX0FvQS8BLwEnpVAB1FhMRQU5zVr+WA/H+KiDZT/exEX3+eaE5nb/0cDrjG2xq16Q93l15ddc1bAS1Z1SWO1qx2IXG5NUfBNzjWG6i4cPOaiGMIBkAYywXagYlUByENgXsAcFt4APgB1EAR8J1kgbu7nerOuMKDcYlgYkWEEh7mQ4tlmDYGwOneRk39nMGCcr3At57C6gOjg4JyRFd0AdjtnO6KNqAE84ByuqSKXzHxXsSpe5E58Mu9GPs0zAJjJl98ppwUfxyoEwoPzd0n+d7TLcd4fbR0xosJigyA7krnc4rz5wbY6GdkA4MZ3kyskj71vWJtQDwPxzAIGWdt36sHv2mR+Upwt8G5xBb2FxrKaHHljUYRVEFY6FodhZ1uHLjjYjRVCF9LC4lncrXLgJoe+bTt/6ePoDsfkxSBVliXJFbzo577vhuSjX9mbNZNkbKbSrNXqica8rJxGYU3ut4R0Z321WjIii4ugjOuoYu5EqZDLFAC91TeUGMu8dcUKtslKZ9UOlt0at0Re2PjXimvRHuP4NELc4qHYdZ6sWOkGuTryQ6cgo5mncbnJuI+1Ku9XvMOwOYOxl3csf3gJeAl4CXgJeAl4CXgJXJYS8ITFZdksvlBeAl4CXgIrK4EOEBpgBOCfxMEO3Za7Il3TAu3Pk7i4Q6QFO6Nvdkf+3yddbt2QK25PXXHbqCvtWO/SWq+be2bE5TeErj6h5+VmXFSVm4I1cy4qGugP4M2CGkAcQJ7vlBErDOYtFtyAmezMxqIAtzE8k8U39QLkNCLBXDBZwF7yxh0C1gpcR/64n7Hfbce/+RInT7O8sLw641xYme0+A+0XW1RwHbtpzTUU33FlRfwJ8jvhKo/3uNHP/IB7+j2flAuol+schAQ743GRQ72+rUSwZPNP3YqnsVJkRYeOKNvWczkgEZA1CbDDyCB2B1MmyoAcjeCgnhbYE6sY5IrMzXUVv0P0INNWwOZ2PsiZvHke3813e2fAciOkOi02KKO3wGg31hIf6JxZK+F2jbbCkof2oS89ffrbV+7XJVwn0X4VkRm4p0LP6A/sAKZPW9D787YCW7larGxOBOFWjgTinp2p1I5kLsgnSSMWUzdVKsQFDcsKch7JEqOA76g5kRUtiwpLbUB8ZQvlc7sgElBbpSItbMxi/Ot0nWcEcGsO8e16QZrgasqUuZV4W4ypWKx9rv2JxSbvR6HG3KrGZK7zh5eAl4CXgJeAl4CXgJfAZScBT1hcdk3iC+Ql4CXgJXDBJMDC1YB8c5cEaAJ4DAjW8pmNxcX5kBbK4x+UfkjpeW7/78du08/e7KIBrAeOu9rRqvC4XpcfyrtmRc8TNhP1RS6cy1xuY8HFZeF1IbvBWUQDkOMqhrmKcwCsWFtAsgDmA2gCfl/Tlhh1oj6A3NQFYLYziKm5frpZ5yEt8CHOTkTy4x4LkMqzuNcIEANL+SQP2+lv7qkWA+adbqGM0OAZZlXA9ZQP9zcVl6WTbuQT693+P4zc5Fe5jvgdtBPursyCBHlwjjIhA0BmdlB+sl33lfowWSNXiAaeD2HCDk1c9hA/A7KFulBOzuFei7KRaDMLIM59yBQ3FMiZ661tAU0A6PYq8Szy4TqzzKAd+R/5AapTLnN3RV7c2wJ620SLEUXeAkNC6XKYfiM3swyirb7Zlnn3uy7uWXTcSD0j5ehLfL/iSSkCcSvQebJt40CtkI+jZpIGhULODfQWMsU4zyZnqtnGtX02RrXk4UHti6ug5/O0NlFBFp3km+n14k+sMRY8zgdPPx/pX7X38p5xvxLvFbi/ZN5lXmbjA3NvVaTFKAG4az/fklGnleiCMbfw/qtWhr7iXgJeAl4CXgJeAl4Cl0gCnrC4RIL3j/US8BLwElhpCXS4zunM2naoA+azKx7wF+AXENAAcK5nBzZgGOfj8yEttOM/lZUFu/nIb5M78jffcUf/tux2/J+r3dAbyy5rntDevnWufqDp8nIN1TjacElFC+rHR2WNUXKFXTnFuJhwUQ6XQuzgN+sJK98OnTO3TFYXcwVFXVikcx/1NcsHyBquRQ4sykGDyOPrSt/TvofnIC9+x18+3w0k53pAe/KmXCzmycuAcp5ru2UhMrjXfJKTB9/Jk2dCOtznaocedNPf2uAe+enQNSfNRQ+AvpWDOB7Ep7DYHhBLnAPUZefkF5E1D16hg3rzDHQB3bB63qjvWFzwuxEoXMP/1JXyEDidXZyQQZz/khIACfnwrsF9L1Ui2DMyR1YEALXgsnw3Cxprb7PMgFiiLEfb+aAHXEse5M1npysV/buiciG/5/ph+ovc0FnaE9IOS4vLaYet6XOnpdMVT1agXG2AukXCKdlue9O7zlgvJ+XRCWp7QPvy7qJd2ueq0OvLu1Uun9LpnanTStO+2zsFumIuFE+Z8/Ue4JZwuUcFIfifUnphe2yBqIbA4H1k/SvH7p3+558/6Z7MLNyYE4wcvXyE5EviJeAl4CXgJeAl4CVwVUnAExZXVXP7ynoJeAlcRRJYHOQT0JvFKCC7xXBgDgCgZkELsMzvuCkChMbSonqulhZaQFfapAXg/EtclpTcM+9dI3dQDTfwmhtcOllzQTFwjfFDrnZsS8tF1NwTgYiKaZdWe2R1URKpMedKO7GkAMzHXcwtSpTZ3AcBlFssC3MvZC6vqBcLcqwUWHizyDfLCdTgBW054M+fZ+BuCYIDsBywECCdPNiNDljAJy6QOt14kA+/Acab1QXPR8aA6w8ovULJAgabq6O73YNv2SP3T8icMlE+/PdTH/LCTRXWCJSdvACWzX0Vz2fH5H2Ssfn3pxzndbStFCAFqDMypizUycgDAA92ZyIHEmXaoWSkAoQD9wKEcx49Qude0k7mxgv5sKsf10SUHxKI5xE8nOfjngt5AKRzP1YWHBZjwXxvo7Ncb4GH7X3GAF/z8c+9Fx0Y1K5Vnm/kl5XJytK1PEu4S2pX/7w/LIgvO2shuyxeyAWPXbHcki+q/0Vvs+WW80JddwbC4ZLL4z9950cWV72TRFkAtv6bF3xsJYnUCyXys8pX89lS9e+0qFvsCtCAZpsflhyPAJ39ceVKoEN/OvsN47DNVViQMn+aG0r0yshL5lPbJMFYzjvF2YwJ5Mk7Du9Rm8Ms3RRnzfWr66Px9w3fEU7kBicHGxNYbpr+2nx6OZHZV65y+Jp5CXgJeAl4CXgJeAl0lYAnLLxieAl4CXgJXHkSYNFpMQUsMLVZHVBbQGZzbwT4zGKYxSqA/TYlwHquYbFqAXDPWkptQP1OLdQBSP+tUskd+/tjblyb7zf+7JAbeNluF5ZWu7i34KJC6ApbM1cfWe1m9+Rd322ZyItjbuqbO1zvTVOuuOtaF+bzchf1UeXzDiVzQQRhYcG6Abg5+I1zgO0A/BANBhzxuwEEBjRBCgCY71PC1dJ1SuzqB8xFBoAI5MOzIBgA2vlupBB5I092LVIGwHbcJJEnMFfTpcmsy+ZKrvLUJnf8Q7eKrIBMweIAEgBQHoID8J58IS/4xOVTy9e0EnXg2X8hudJWK33wDOoBsIHceBb1gZggUY7nK+1sP5id+lzLdRBJ1IXrKSf1uEkJUgLdItgz7cEOTyOFaEMAGrPqoP7k/TolZL1fCWsN5IA8ISY4T9kgcminQ0ro1o52/ugt+UG20EatwLYWm0XfnQi4swF5uGXZRwdJAZFC3dAhym2BpNEXZNYVbGq75Oj2vBbAJZccrbKzE7cup2vRzS5QalWL06T0oAvDrfPfk4cHW9ZVP7bpo/k7w9f218ICuna7ErLGtRd6je5fNqTFsoV9AS5sA/Imy04AvvU0gfDn9dQugHdn21neiwHvk8+8DABtkwl9zPotRCQH/Z5+13LXJlmi54yd6CBrDc4vcGe1WJjnK1/1HyMJzarQ5gPGAhurzSKLx5tVFuWye20stzyMjE4ashkMBlQfRVsK1ioNujBY4/JBTu7sFJFJeWD9ZvMtz2RsJJk1GmPh2HA8mH5k1fe2gGDV+YKNR+elrP7mCyEB6zfomsXg4hNdYI5gDmWDA+8D9r7BWE3fImA235lbmGeZT08hE05Demean2ZFUPRoHsinQVjaNbt39xtPfKFSSGub9T9zPHkz15obyyuOdLwQjerz9BLwEvAS8BLwEvASuHAS6NzlceGe4nP2EvAS8BLwErjgEuhwCWWuewBPACVZiHKOT8ATQBQWqBYHAhcBACxYG+CyB7AYQL3l7udcrSw6KyywDr/JgKXsuAfIzVzfTTvd2h8ruvym1UKS6y4eXCuLi+OuvLsgF1GysCjHgpEyN/mViut/Wc0Vr1GA7uKsK2xiwQ6pwBxmFgAs/A0I5juLbcBxrgVsN9dNBlyx4Lfg3JAzAGwATsiJfABycWkEwIUMuc+sO8jP4leQD/cAWPHM/6KE/Aia/SKlh1ztyHZXeWLYjX1R5FB9mzvyt/tdfZj7aB8AAkgjwGR8SvMsaxcACp5LubCq+IpAS4iCFT+kO9QN/aBuECYcPBe5IUegccgsiwPyz/pOnV+rhLxeqYQVBrpFHQABIRZoC8gbftvRzo/zEBo8C9IB0JPg4zwPSw3ajLgkEBCQH1hkoKPIxe5DHsgL4gI5z7vZmicKaBtAH/KhTWhfA+UJKn9eIKGAH2U374KDo01UAI5SH0iXV3FaCVnQhhBPtBu6ynnIAsDLBUTBYrBJACx6NW8ZVXBpuNGlgXqFvrd23mbjbiDcJfk0ZdnSVH6hK2VV1xNIq7KaAK2G2iF11W9veVHt/3Lv2Xg025Dbn9v+WgWTiXqbM/fWw/zx3ubsY+/7zjuHXzV6T6drs65A1ZXkw1yAupG6NCF1N1nTZvyPngMIAhx2ukZZUneWAtzbrl5sTDYrLwPGydtcphlpaNZinbvy3cUiLLpYUiAj5GU6juJTNuLOYKlGH4bMpI8zrqHjd3KTDvoxdWRnNwekhllvtU/Nf5yJsOhC6HW2IVkA7DJWMY4xJjGuIFOezXiO7CnfDiXmum8pMW5wHfcyLjGmMV70qsbUMRf0uFkREydUi1S5rQnKrhhuFvk6b+t1TH1yu355UlrzbUnoNfpEb9bpflzk9Sgo0zfU2C2Lpsmo596ZqNQciQYOP1zaMZFPG9Fk1BvNhXnK22mJNS+UjuNM8jnlBn/ikkug3feNoEAHbf7cre/0H7OaQBdfo4QZE3MdJP8OJeYK3sXQye8oMecZWcE81xqPGBtOQ3i3LuHZj/Td1PupDT9YOlZYv219bXjX86Yfa1w3++T4htqxx4bqY+RlgVPoswuI9Stp/L/kiuEL4CXgJeAl4CXgJeAlsCwJeAuLZYnJX+Ql4CXgJfCckgBju4FfACUASIBNLEL5BBQGpGGnPr9Z8OmTu0l1DtAFgMeAlPMSAEB720UU4O3blba56UcmXX3iy67nljeLhAhc+ZpxF8QKxj22WoC+Fs/JnOJZ5PV7Ue6hYpeKxKg+k7jm1IDLb87rXKY4F8ROAKBiUc+inDqaH2YW9ABRnQeLcq6hrkY8ACQAFmERYcAcIBzXch1gAXJDFhA+fHIdMrJnAiJ8WgkAb7VLGje7dEK7cZ/Zocv6RFpErjHWdMc+ctglE5SXNoKogBwAzKb8lIfnPKoEscPzIT+wKjkoGS6MwqqTK3hQf+pK2cx1FecoH2QK9aOMAC3IF1lBJAA+WnBsYoHwncRuUfQH2WKBAREGkcEBqI/OAeZzfkc7X3OFgTwguDi4hmfSjoA6AKOAoMie+35YCTl+tn091wI6QpLwfHQdUoi8AYLDNrF33sRF+3l88ByA0uvbZUEHkNv3dVxDX0OGECz/Q0k2Eu6ESIoWadHaHf7zratbbqS0k5salrOG25qFwZawlJX1S2+WBS5oZgNpEsRBKXu5KJlNenp/cjj4pIDVmSCf3SYNjSSBp6XR16WNYO556WOjvxr+RTI11pt9NXzZzkdKN/VcW3kyv3Xu0NfWVY4P3zL1kAVJR47IDmIIWRmobiD9eRE9HbK4JF87SArqgQ5TX/SMfgULRVsAIkJU0seRC8Qu5w3As2DvnQTPKfXpACoZh3mW7aiGgLPxBLdv/N/yJa+E3tP/cQlnO50t4Li5tbskstNDqQeAPv2LTwg3+i79m379c0roLiQhskTfGX9/UIm+99dKjC3UGTD2JNhqFVoCcLWNVXx2EmmMnzybsiA/nkGfI39W8OB0AAAgAElEQVT6H67leM4dSpDHRrYwfjCeAQozRnE9B+5y+F5QT7xf6WbV5togdGPBardH6WCQVxtFIgQhKiL3VllWrM/mRLQWVYZQ+QftzQCLtoIlQfiOmi5uiEnUTvYjIjC+urE59sXybPX+h0o7t4Qu7ctnDYHRweF6EE+KmPAWT6YUHZ9LEGlcgW7aPGz/nzJmXUzCp93/bY5nXofst40Tr9Z3xh7aGXIbnWTMpc/f2q7yD+kTEp8DPUa/uYexiXGCsWm5h5EkG26afiRcXzvelEuo9J7Vrxp+vPeGue+Z+Oa2YjJHf6B/8r5BH7bYXct9hr/OS8BLwEvAS8BLwEvAS2DFJeAJixUXqc/QS8BLwEvg4kqgDcDablMW7wA5LD4BHwHgzK3Q/NbweTDJgkIDpBm5waKYhTPgjs0PBOAG3D1v9wBtwP0RLeb/WPkD5v6gqx1e59K5b7tK7zVu8t4nXSoLhMKmxK1/e49rTsgtVA+WF7HLVJXhf5px/betcbPfnXazD866eMOw679ZwFRRYFFxv4tiA6WoHzJg4U39LZaA1Yn6toKLK9mOaj7NnQdgB6AWwCKy4zwAHcAmwDmyMHCdBT75jIhfabi5pze7qHyTa5wYdmk66GoHGi5r5OXaqihXWEdFVlBG7qe9APbJj/sBsgHxIXQAzmirzyjdIblZu+nfC3PQvmpnZEKd0R2AVP438sB2KyMnAMJ9ShYgHDAGAIXyQ0YAZJrMqCdgCPkiU4BZ8ubgPjsgiACJIUKMrOA32o/EQfBvO16vL8iStuSgPcxFFW3/oJIRLoCa+5QIYE6dWlY29JsVsLYwixIjKQCccHfF+c4DmXBQN8qGe6xHrvv7h4b/6ru/JPuIe1ruQrRbu1c1uj4rBrmwnJVcLdgwly/0pBujNbmh5PnNanhrnCaDYS5bFdZTqbyQp6EwbOSj57np7GAhaazPDaaJ7EzeIukUoiRr1IKwdv3MnqceH9i9MQ7TQk9jdjjK0sHr0z2bbio9OloqV7cEDbdGXawmie1VouzonLlCa1kZCFA2q6SuYP2l3oG7RIwF2trAS/SCdoBcAvzDKghgG72gvox9L1Ni9z2/Y7GDWzPGAMBD3I8xBqCnjC3mLu8kkdNhTYHszBUSljVYhPFcc7WGThvID9lmVhb8jrwZw9ihTz70tyPKmz5i1h6njMcXyAIDvaRMyIAx4PuV0GHGCMoCSYAcFx//UScgC63vMgbIF6CD1CQv5Eq96hbv4pfmCTs7jDi2MdtAfMYVG3cYKygHRCayhRiFIKFMjBVvUoLcBBDGuo/d6ciN9kPGL+543o+2vrdGBvc69cNttIgslpz6hsugxTWKhHqK3K45WTu1WiZYdXIsW1B4/sEcox7Gbjosu2PxqtZ3jTibRF68rZjV3ybXUAfqQW5GfXGqnNbev7Y58bnj8apMekz5aldiHJBThHTuJ+x9h0/0iY0EkNvoKO3PXGDWiJDbuCnLLqQLLvVP+gr6ypzOWGPkGVaBjBFY+jA/shkBfew8mBNtXrTzzFuMO9QRgg9dZwxGd08h/BblN6/J8wnZMC8xBhXX1EcGkiDq/96RO6uvGLvvWF9zepfcQjEOQs7aO+CZ8l/0OP+vl4CXgJeAl4CXgJeAl8DKS8ATFisvU5+jl4CXgJfAxZaALUwBcEkG6LCANuCMBTQLe0A2wHcWxyxK2dUH2GzuaswlBgAz9zdXgqzoFAgAvBb3H2/nv1qWByTKAiDXIyuKSZEXLMzZTdgQgaHl/4ZNLl4zI183VbmLGnB9tzZd7cE1Lp1+WhYYNyi2xTqXFHpcOHDCxQrWPS8HFvgswpGP7YI365OWi452AiACZDBw0+RpIKJZbQBAcA8ACJ/ISKTE0a+46r6Xy/Kj7NJZ5ZMddPmNCiw+M+OSGZVxbsyNfEZkxh4AevNzjmwhLCgn+QHgAYJyjvYhfXwlA2t3tsES32l79IWEfgCWANUhBwgCgCBkZe6vOA+AixzMBRLtxj343AYQROcIPs796Bj7k7sdyAAAkgPgmHw6iYvF96DPnQcuq9AX8gEcRZfIw9xaYP2A1QUgKTJH3xKRFtly9dtcQdlD9T9lANymjrjyoI4AUqc70LtfUfplBT1992/v+91/en76UI+sI1Lt1t4srRpKV0dvqK7L9+YLTfFwbvdsvbT9mbUbc8lgVOrPKkEua4oNytyq5rSba+bDXC5xjS1xpJ3cO/KzdbcunpSD/XQerQqz3GTanzvRt/bWm/ofd9uyw+6z9TcNrm0cF2P4+Rf2lCtvCUJhuJl7Optw30rHBJQ3JJ/M3a1EO9Je9CGLBwCxhuw4TLZmiXGGql/Un1sEkJK5YYGAAMRGRyDOANOxzqHfW90WFxDyovPAJcvfK2EBBbBHf6U/A4w224Cl7YImT87zHFyW/ZQS/QHwcPEBoLn4gCxh3IG4QOb0sY8oIXvqhI5bnIgFrqO65LWsU10IH+THGIrMKDt97Dc7MuO5RhgufgYAaCep8p/1P+MJcmGMI7YPlmOP6LmVtlWBuc0yIhnXU+ZiijYzMpQ+DBHx5vY5xp6ljv+t4wfysIPxdeHB01U6WVJsC4CK0Wo9SdYVre8RtiXqvZFRj6d5aJqFbjIuu9G4382GJXcot8aNR72t/zuOk4Rt6LLb1jQnf7sa5veLwIhjl9wpuQxLLuccQ+o0xXsu/2REFvM5YxOkHvMEcwaJGBA/rcRGgv+qZBsT6D8VyZTP8yYuFsWjoUxGpEGcQZAxNjJ+2LvIz+g7ZTbL1eW0AfMm9cDiigPCw+JbnGkDCdrMWEQfgsRBi+nHkBYjUZY8X24BC+WgMiHmnrkS11Pkz5jf1WXbcgrsr/ES8BLwEvAS8BLwEvASWEkJeMJiJaXp8/IS8BLwErg0EugkLFicAnKYiwTzf0zJbGcxi2Z2FQO0chggb8GWAcKYH07rU/t8qtoG4gHgCCLM7j+AX0CxfUos+A0EPyF3So1WYkE99jnKBfjMbkq+zwMV/S/pcRt+aosrXVNxhe0VV9pxSNYZ610olGgeqAbks12ZAPIADEZQAKJZUFgAOuptLljYeW0WJ5zjnrpLmlrUZzlXffKES2uvccmsogxUBEgUIpcf7JN1iDbYluWk5+G6G7tjn8gKgH0AN8sP8sMAQcB9ygSIt1+yYQf+pTjQC8AKdMasLZAxZUNf+ARkAwhBz/ikrZAZwC+AjJEeACPUl/OArOiegTqddSMWBr937nYG6EXW3QgLQGIAY4AY02fyo1wkygmkyO51QF9IEPSZA33Hzz7/A/y0rDLmOYuzjmtBXdBZdsryCWFB/znlUBgW2nWXdld3AqZRKZ175/7y9huSJB6sN3JzjTBsNotxfm5r6YXDm1ftauajaCCadQPprKsWC25KO7Vrad4JbHJjAj61I9uNRX1uKJl2mxsjMsbIuaf7Ff93br/rDyut/+X6Q0qWuFqi+/S5Ohh1m+IjLt4s8caRiA2VSpqYDgsATtw1obQ7k4SzivuFk7TcfI3Yxf5lpa8pAeUCfiFLdq0Dcs3KAqNFAMrS4kxgWjcxrdQ52+Vs1iHoKSAm4Dbn7lVCJyEQzvYdGCsakh24arlbAPPfbW8cf6YSFnq0U/42nfteJcBGXKb9r0o/rrR49/SZ6kuZFx/o2eeVsM6BsKA96Av0uYa0zKwvuuZ9lhYYRvIiM+rz20pmLWH5L0VW8Hs3YtLcL2GJBfkxHIqm65mdO3bg3UNT7tgYbUW/hi4wUgxC/SeUcKMD4YQMVuLgWc8e1FbagLunQDNFqJEnMBsz9fSMWYYev4wjUY+TLrjpqOwO5ta6/fn1TrErTnun6MX8Y8VtWKW4OEuODzWn/vVE1Pvw+x74/gOzYXHuQloGLKNKF/WS08RQob8yj7ftW1r6gKUm8wRjzz8pQZS9rV1gSK33KZmLSIg/yFfmENOvZddtEUnBfW2taY0rlAnikXcZe5/ptAi051B+dLrTutB+453H3CYyN0EgMB9DWlBue0dZyjUf5eHgGWgvczNzIfli2fSu9u8tF46al+7SXMJcy/sG4wrzP0TeKeP3pbaeMwH5Ty8BLwEvAS8BLwEvgatLAme7WLu6pONr6yXgJeAlcBlJoCOodmepbJEKWAxwDBDDrr753f/zO3yBW8zdji34bSc/eYGmAASxm5fryAswmnxwFbTiVhYLKjAP0D8oQMBibQAK3q1kO20pF1tT2U1JvdgNaBYiLK5zbur+p+SOqeSG3lh1Ay/pd9XtsStur7nCtmkXD42LuGDhbmQB8uB/ZMczeQ6khO3atx3L5ioLqApZTMjNU7+IiRE3t3fM5QYFiDT75eap7rJmzuXXVV1jKnKzj4240TumnXbKuhMfE6ibAdAB8M7nMW+pwK5G6vgvlL6u1BCg+IlOuVzs7223UIA5Zt0C4QAIj5zQFwBaQA3OIzMAGcBfQBY+uY/7kRfEAe0GMEm9zQKDHenIgwNZPNTOBz3lO+0M6GQH+ti5g9osgNB1dHTxYTvmAThpT0Aryk+56BtfVMJfPefQewCh08Yj6PIM7uXZAMcAT3wuRVYc6W8qSERYXt8IF27kn476dv2H7e/ete3IgeTF4ddr0+X8oYHqzGBjR27tvr71gdzFiJSYdPflb9Qu7WLLxUzncTg3/8gDwncfLFHN+ePJ8ma3rT7sCi0PXypYfdY9Xd/q4rThbgoed8WkqpzkbU34NjHtOWSf1IKJM9FqqTQzBR4TpIdLnFaLz1sJkOxAF0gQABBD6AekHK6jkHUikGspYK0jm7P/ehpAE71DVwDLaSP6McA/fuIhiwDeAb9X6gCg3CIZ5gaTmc+qDWZfUnnikABnxq/XKGFRgAslpLkSByQciQPiiL71d+3/ARoBOOlT5yt3ZGcubdDtn1VaTFasRH1+T1ThTym9Jw2DB/R5o3Z7o7Q8m3bExRNK/kvLfBg6CIm5nGN+/WOzp7pWoFEs1CiERUWgUSjAJZRGrgwri4X0RkvCqShzrmsRHSqtqD95/wtcoxC70aosK7Kim5LR35nIisWFbQbR+qO51f9YTOufVNyLD+az5t3S+fGribTo0oC0F2M+eoElG9YLjPHMRXbgAowxiBGL67GgItnxZ/oCifio5AnRVz1HmdoGEfSUuYyy0D/QEghsxpvTHcyLXL/YsuuvdA4CmPGLvCGCmUeZo+gXid4RuvbtVgyk+TqjkbwbURbuY376VSVGeDvoI8y1WLli2WnvWYwh86O9P7wEvAS8BLwEvAS8BLwELgMJeMLiMmgEXwQvAS8BL4FzlACLVEA6Fr6AxuywBRwzdyjs0uMaFtWA9CzSWdCzA9D8LHMt1wEkm7skgB9IC1sEX5RFrBbjHxVpQRmwiACMw2e87Y6kLOxMBKAwKxLbCQiQcatrjD7mjv9Dv9Kk670ldVt+da3L7i263hf0u3ht6KLSAaXQ5TcAVLNDmUU8cmCRD0AA2GfEj4ESDVcf2yNrjd1CrmJXPTYiVLfk4tU73PQDMy4qllxYAtoadzOPKv5AMXXJdNNN3Dvh6keRG2WlPpASgAc81/zg017vVfqS6n5RZKxnnelAppSFT9oC8AP9AOQALKE9TDboHrs/2cmJVYZZZmAxAqCP1QF1BIRBvvjuBsTFtQ47YyHU3trOm3IBUC4+0E9AFaxqOMgXsKeT1Oi8B+IDgsRAYsAfC7CMjgPi8GmEBf0CUi5crmsoXY9c2C1OOQCVAMo4AOpPbqVeVxv+f7bOHRx9zeiXjxwqb5744po3rBnNDW28sfbo3KOFG9G71vGuDb8f/XbP75SKfSO7CvFsrJgVbkq7sznk576zbsv6LsDT7S08iy8H8nHzWPMWN5KuaTVgTVvIy4GsNkLFs1cQb8gLOwBgI9FQ0mYXiFYDrE2RFnDZwn23gPUkCADGlX+vBAgGwIwchgWi0Z/qF4q46BCGjVM8Gz2jzbGsoX//gFInaLksGS66CNoGvcVqaPExIHm/cyQauHVVMnNIxNJwb1p9FZYtgq8ZwzggKFf6ACQlvUPpz5XQQ8bHO5TQaY5zJS7MnQx9njGrm8uqzvrwTK5lXoFAgVT8xeVUWOp3S7WYf+uDt113/OX3PPzU4MQMY/GvK719Ofcvuma5ZMX8bZAU7VlOsSieVFyKjfrMazbNMwIqpkumkSOAjIDMaB3Es2B0bNm06DsaLmIvqQeuvlqe1GqBiEG5aNM089D2ne54sRunqj4mKynFEThtFdU/f0jk181hlr0/55rvF8jOvLxkm17MoNLn0Dbncwv6yEDImMl35gzmj25HN5drdh1jAfMGGx4+qNQiLc6yYDzf3hGYA5gLsPCgbdCSM5EVPI7xEYs1+i+WovuU2MDwKSU0Cw2jXC1Xc+3rm0ZWdAlO33Zm1nrPYwxkHkbxsFrk/aLbQRkoP2MG1/OOckqgbW9ZsYT0/GkvAS8BLwEvAS8BL4GLIgFPWFwUMfuHeAl4CXgJrLgEOv19A5KymGfhyUIXaBHgDnCDhSi7+/nOjmjbU2qwC2AaoDqLYxa55MMneQCs188CyD3vSraB+8+JuGAn5A4l6kZ5ACLYWWm7Epm/AMLZAcxCm52IWF+waM/czEORe/ydgl3j1W7odU+51W/aqngSm1xhS+SKW+qu8tQet+5HGi7sW68YFMcVI2O3Yk7URUzgpVzggXx61I9oK3ph0DXHr1F8CgUkrlf0f+wqjxdc8dpQW3ABRkOXJoEsL+ZcffSEm7o350Y+hbsJysaubuROmWkDgD1kCmkBYLBP9TVw8bxltxIZtK0s0A0AUBA19IyyWmwUgoJzDmAFImGHEpA2gA3tBGACcAlYC3nAdcgJkgIzAM5BctgBsdDNXQ47yAF0AIeMrLB70NdvKFlQ4o7sWl/RYfS6EyjGCuArSgBf7H6nn1AO6kkZzwjuVn900CluhVnlQK4AVOEjv0/g9CPaYX0S2N01u/cD73rqD3Obq4du2FV55qbRgaHnr86NHr+v7xV93ym8YIG7nPFwlfsv7heCV0afi7cWnnblEHGvzMGu75m46Or5zD0ZbXaV7OUun4bu5uhhNxIP6HvN9Up15dZowQNjoC5JHvdQgbgTSIvMIiacKiksbXDHAjgGAAZZgFwhHI8KYAOMM7/oS1qznCM4ZmQFOvFaJXSFtsWagjai3y33QEfRCQg3CAr0hF3c0DXdyIqT+R7Ir3uxLF1ejFXLzvpRWcZMtUDpMxyMW+gqsDf9CpZKOhssAbwvqaLERMHtGHkhh88oMcbQYmcsxKIyIk/6On0HywrIuG7+jABX6fP0q08rQSS/TgnlZTxAfpxjfEOOkJVdj2YcvWP9sfFNxWqd/ryc9lpsddWZL3U3aznGYOYF5jbGsuerO8TS67sVVLsscqIs10+368wxfW/KoOnHNbKtllXRmM7FsrCY1PXzu93FQei3kiwupjRSzInA2KS4MxnXZWmQJcNRMLplwFVmNO2OZO6zNy1Z3VZZt47L02FvXn2zpKDcJ7nLU+QjMmyXyvB7haQRxmHyAf1/oh3vYylxPmfPL2E5xVzD3P/Stg5hndBp6XU29YV8Yw56oxJzzof1zK/qc2qZlhaUBX1AR8kHQpR3qh9SYrw508F7Abr5fiXmN6wreWe7X4k+ZhtHzKLCLD1bY2YXosI2DjBHQpZQLvInz99X4t2o28HYfJeSuXCENKlcBGL5TPLxv3sJeAl4CXgJeAl4CXgJLJCAJyy8QngJeAl4CTz3JMBC1XbVsai1wKQsiFmEWqBFcw/CAhYgHzCORTbAEKA0wRyZBwDIuI/FLotlyA6IDiM/LrqE2kD+STC/HdAW11GA2JQfwIB6Ul5AcuqKSxTQH85xaKHfHFbci2uVxlwQbZB1RdGF8biLBl/gDn9g2kVlgWvpKhEVz7jVrx9yM0+ccIVVFbf2J3e72qF+WUnU3bQ2jufX5F1xa8E1xnOutGXOzT6syMflkiusi93ElyruyN98wtVHKBckBc+nbLQLfrPZ0QlA8ajqdSn9+y+rHdukBSA+4BBAH3oAOM8nu1LRM36zWBDmwgWdQo8AX/DhD1AN2ASRwW5OAM4dSp27Y/kd91yLD9p5qQNghmTtvJx6EVuA6+k3X2qXj/ssLgnfz0hatO/v1w76nWkQvkX/t/Zed5IVN04/9s+vGL/X3Tr74Mt2Jc/0F/rrlQ2549f+YvWvc7tKexslxYT/WrawenvmbnK5sOrySttEWoStoNltd03yLab/FvqDOk2NtSN7Lg0EybaPgvLcXnzSHa7tEJI85AqxkOE0qU0G5b5avMHtEsDeIzdRUadq0oo6BMq6UDBfKmchgTQai4uWVneXFO1KOQ1Q/Ed9B4gHEANQ526A9HOyJloiKDTPo/8zHuB+if8hUGjv5RwA7tQGfYVQRLfJD6sh9PqLGmylv9mY2vgaWaNU1BZLgur3l6+XFMVfgnyLtJA7n5Pt2C7Mf9cnfeceJfqPxcfBJGYoCyKNE8GLBIFDzu7MgpYfsbkgS0UCGdfcVfhvaOf/Sn1CEECw7FNiHIfIPe24I9la5swHkB4QNT/fRYCQOrQnYxoyY1yjHpBTkI+MF2iIWV00c43mP8jVk9okuK0RR2+TLdMp/vv379jwunXHx92akQlXqDacru/y6JOnsJiCmGBOA5SlD39Y6YPt5wNGM97IHV9rzoNYOCpLiX/W6DQot081xae4TYTEDRAP+u0mibamFCnlFMfCCNRTduvLAulZMkmaBiFYj+JgdGu/e7SwzR3uXeOmN89bRy11rJmYdNccOuxy+cTNrCq7kcGBFmlxWIG5lzo01vx6vtY4rrJ+qm1pkSwTZD9tWS7zH9FJ5g7YH/QRiz3IUA50rlucFNp7uxJ6iZ519tVOF0z/Ur/RzhYTqRWEvUucChMRek1ZmOPpI+T1b5UgRS1GUjdxQtyhi3+sRJ9nbGLTAnMhBDrzLMQaCs/3TpKiW352zohFykE9kQ2bBMwCsTPWzuJ8IGnoq7hG5NmMy5f9e8nphOF/8xLwEvAS8BLwEvASuDIl4AmLK7Ndfa28BLwErg4JAM4B/rFTFxCMxSuoB2AVC2IW5HwHQGLnM9cDDrOIZ6HOIpndsNzPb4B13EeeLMKXDZJeaHG3gf6HBSgAQgFIkNjRDgAAMM6CG/CYOgA0AqqxSxj0iPptc1mi6MOHAe8kp/1cYwA7ANgJN/4FFu4QOrGbenBEAbz7Xc8tOdd7feaqB5uKTVGUk/IZWWRoy/qxOTf+pYddYwR5kw/5cT+AHmUB2Gf3JQAKgbTP1vXEhRbpafPviGdh/q2NFDMiBoAVHWEXNUQAu5jZzcx1uAZC/uy4Zsc7IApA9eeUAAEBWJAb4BPBQDkAIAGcz+Y4PTI4nxNgJmAT1/K8LyvtU0Lv0Q/KQfkrcgvV8hO+uACSxclTcvGUG8mvGZRZzeRs1AOoveDYWXnmA289/rFD24MDx7YPHHhxsbd+jRxOjUz19/Snm9LopvA7k7OlyD02tdtNNhcaljwy+yJXUrDs4uCcWx0Pi7xQCJak8Uw9jNf1pNUTSRD2NYK4R0TGiGJljyZB0CvAFNBuHLBV31tWACIrqANk31CaKQBw0iuyYrubTfoc5EXF9eQfye8cmYzyT7gwWSc3RoM3Vg/096eVrlYB2n3ucmpJ4lqkojgz9aBWbItTIS50gb5oB8GmOegXWKKgH4w/jDFGfZwrUGaAHeSYuQHbp+//9+I26fI/4Drk5l1KuGYBULQxlMsZS5+UO55EQbRrsUtKkvtr9f+1q5LpooIh36xg59ignHKU06r7Znm3eya/wb1q9hG3ScHQc1ny62qzHbqYfkAfgFzFisMsIBg/imlQKtXzOwmDfjhM5z4TpxPyMZS8TFzVmjCd/a6+A0r+1DyRtaShCmW6u533u/UJycs4BCDblQUQAG5ubujbtCHA57/rVj+dY+f2v1JinCVfxlPKz/985+A5wTVPHZ5o5OJ4y4HhUTVWWCvkBg5sX//kTG+pVOkpLiApj20ccv/zra90b/rM/W7rgeMuX1+S00JuyA8imLmAeY3+/VElSBSIVfQMC71xEROzIt2g74LoJo09Oc0b0BdhK3j6NvUbAGdz+LRElZc+rT7ppA9ub35ji3Ag0PZSx8ajo42h0am5NAr6ygergfq0WxeMaxAadsFuER/rc+5jA69skSCLj0YYDTWK0ftkhfLOtcMTH5dVivWfsy7zc+QGs2TjXYWBEhK0M05QJ1lhsUsgAD6kBN3KPAwx8GtKWAp1O5hvIFRj9QGsHCrBCz52Sh/RO4dtEEFP0BcambgqkKQc3YgTzn9SCVIAUg0SkHEZyyTmQiP/mXNIbqn4FFbwtoUFZTE3oIx7O5SwaMTt3enMeuiff61E/6bvMO4hI1z2nROBbOXyn14CXgJeAl4CXgJeAl4CF0oCnrC4UJL1+XoJeAl4Cay8BMwFADlDTgCAWUBjgF8W2yzSAeBZtAMqA+AAjJE4B4BuFhhcx/8AtiyoAZzIr7VoF1DbWkhfTkcb+McVEQnXUYAI7C5+sxIAMu4OkI3FLeB/FunUjTqamyMD1wARuJ4d6ciXeTFx43fOKqn+ofLXBvd5sAGQiOfxbIAU8gKYR048G/Dsn5W+oHJa/peT+M6qLLS/QHzqDqDBTlH0B2KGAx0xX96QX4C8AEsW2Jzgo8gHcARgBWsegFTAndcqQRSQB+Dix9oyRFeXuzN+uXXpdBRvliEA1BAnkF60t1kB0Ma2w/WU/L/+G7fm/nz862uf6L3++sncwNbZ0qmecnZV9j7vdVN3Dt0y9HBffk1j1XShFNequca+nRszrBVmk7BUUZiT7fWn3HdnTsWXDtV2unoqXkyI6kBj9u519YmPH8qv2SoSYq8AzmfyrlGJ0uzoifxAOXEKJB84ERjuoHb1o2/IFpIIufL5hiSLc79nuA8AACAASURBVPWs4KaTQdcTTbshESETzdVuLFs91RtPXhsH9UEFi36m7uJv3FJ75pZVyey6pVwZhdA7NXc4HRPZecJNy0XUixbRO7Rpt23i9DvbAQ+xRZ/8vJK5RzsXSy7abYcS4CEkIzuw/5czKAXgIfdAqLGzGKCT8Q5rAMqAfkTrmhNBfzKb3VLdV1bQ81Vyl9U7F+Z7psLykADqF48rWPrx3CBEhHu4SHbPHjXFBeEYjfvdfT03fvz5c3trG5tjs0PN6a+LaOCZjBE8k0S/Muah8t3dx4Nc80ihZ+4b41E6EZWqD+byjYPjYVbdESUTtWa89nejZPR9hfrePwqzuRfKCkP1ybB7wapr8YEuAJQyTjH+3amx8pDGpW4uopAlrUs+gLjsHO92UGZIMdqQcY76tKM5uLQzhkJHEGDy3iDi4sUTg73lKEl2Hty2fm0ahq5aapvxdDxp/84NsrKYdHGzIiuL9AGxN5QJkgciDKD3s0oAxYzXANS0G2WHvGDsoU1bVlORaBclns+YzTjAPMHOevSRsYb589RCdK/7KWchFrCmmYmKijUzUBFZ0ZWtKDbqe9YdHX9ycGzGlSvVh+r5+JnCTH1//9jM7VGavrOUD9elYaTQSIF763X3uW+VrnMnFLtGOnfKMxXv46+vOXj4wFhf34EvfugFzzz0/F31K8zSwt5x7P3GLMUYz5Y6eIehX6EPWM8xhjO+oweQaugOc1C3g3gpP6r0m0ro1kl/fG2igveIebdg8/Pb7ygx3pzuYHz5gBJjIfr4V0qUcZ8S+gpBuOQ8Q8ancf+EjkH2kQ9xXujjTESnIysg+f5ECZn+DyWsKyAwGe/OlTA+gwj8z14CXgJeAl4CXgJeAl4C5y8BT1icvwx9Dl4CXgJeAhdUAgKNyd921rFwNjdOEA+A6PzGIpZd/SxEAXn4n+v4nZ2nLJIBafidRTzAMLvfyQPgDLDHdtoBwD8nFrJtYuBjAhcAHdn9+MvtelB+AEoABwBSPgEwWOgDvBlRgXD3KQFw8B1gAUCL7yJ55OB/HhxjsY9cyAtZsUMfIMNk9jv6/pDKczZuinTL5X2ItEjapAX1MmseAH7QNANdAVHQMSwY0EVkYy47IHTYGYsuAgYBLqJzgI+AnRAhAIqc36e0Q8lMD3ge7XjOoKLuRf9tdyugJm6caEN0g/bju+145VmqsmDS9iHgKCTp3+IDLijePP3IlvHcqlc/2nfjO+0aPnuS2dnbJ+555pdH/zJ7Qfzd6+Read1IeaDn4I51+aiR7ti/an18PAYfdfkBRbT+nr6vyPAidHurN7QsIOwYaWxI7xl985dvKj9weFXxK1+Iw7HvpHFYbsh3fZJFI7msWZ3NFQGaOFpkjAqLLlNmyom8Acogij4isuInZQ0SCiwX0JxdU03LrpL2uMF4dEPokpaLFPnF33k8v+qvBSLfv6t29NC2xvBvC6TvCsqFu9yGcKu7Q1j9J5KvulI6IuuEpAUgEwj3TMfPtC+grzI+AXjTJpBZI5LzaUG8v5y/Gf1iDETXsDhAl7j//zjNw3GL9B4lrE4Y8wDwGCs5jyxbwN2vnYA3OylH8n15O//pfNJ4e39SoczrtgYn3Fyt4DJZ3ojccCJ8nCwuWo9POozSTsQDbxVp8ZRIj4+9evahT8tFFGNPsngn9QMHhVS369aINxUn+n64WG8oLk7pX0oeQTMO5g4U0uNh3ZVzhWzqxPrxP/mj3sq91+SS4UcEmfcHWeNdKrZc1ZyyOfwdyhYdob6Mb3+vcZKxK7UytK0rKDwkHuTGUmQFJYSURNeIWQEIjNxOcRCmdqSvGyG4W99fL7dQz1s9Ovmq8lzNlWerTqSFe2r3qRjy8Q1DrpGLnID5TxVq9cejJMWFFmML5ab90G8IY8ZzxhPGEAiUVh8wP/xt1z7IlU6HrjAnQiqjq6eLk2FznxGz1PuUw6wgCHCvgOvuUH5d10AUKsB4PY6/dWjL2kdlZfVVWZsc23pg+LgsSKajJvZKbjyspe8Jj2Y91GZdz5h7ycbH3dHcandvT9dY5+Hw1lX/rnekcl89zP3j99z/+BOSN7vknxPzdVdhLjzJGIY+ohxY+hAf4qdOc9+f6jfeZ5grcFGGfrSIRyWAfHSVuQs3ad+rxDvQ4mOHTvyB0oz6A7GRxjUW2DiDBSdEF66gmMdOR1aQB/qIrmJJwRhCn0E/6x39vmtcmS4khZUTmdg7CPoLAUln/xkls/LoUq3WKebXv1FCBlg2MjfTd1txm3zciqXE5s97CXgJeAl4CXgJeAlcDhLwhMXl0Aq+DF4CXgJeAqeXAAtWFuAsWlnM2+52xnDAXXPdxKIUEBkElOsB5Gz3LKAyYB1AJotYDn4DzAWANtCWvE7rQPwybSzqDVjxR0oAsQATAB4s7gHsABwAr5AJgBWANecAyjmPiwQOXL0A/kBcAJRB7ABqA1QgI84B7uFSBtcygBGAXIAUlOGKOwDwdQBwAAoB5AC8AugBvOByBoCc+huwiOxoA9x4oGvIGn0EYARg4XdctrDDHtnuUEIP2eGKD347TveOwi5R2u5MB88AGOd69Jz/Kc9dSugG7Ue7LtD59g5xykwZeuaiUvFrq16aFtLabY0wf2sSLPT90pdOH35zcMc3bxv89kviJOk5sHb9/upAPmnmY3ewZygWeH2ynFHQdFuKzzgsHxpZ3j1RedazVDOLw4eqt7121pU/3AzDR1/bd8fjpbSe1qKepB6ESnFnORcAX9ppnf7hnb97IiwOj7ss3psrj5VHGhsnnp67/qa9czcc2pg/eGRrce/tvbK06I8nBjt4GScy5TdUxo/tz69/+A3T337vlvrILSI6AIgXEwGRWvYtwuoflauozwWzblKWFsSB+KASMSxoyzO59uI6Em1vlhfIGZILHTmdixLahPENPQGEBIxe6FvrpKRbwNxHlBjzvq7Ebmd2YENinbIz/de+0BpH0WVzkQTYTh7sYr6pHVNkNMqy1T3yiYU7IOJUkCpBoVkN1diLjrmwcO2h/NrNH86/PnvN0N+26vWAjb4Lr6VehWYzHUrStL9SbWSNRjIbhmEpzsVRHG4ZCBRopxKuOd4Y/PWn1+Rv2BvV9o8281vTdZPv25pLjr9HFhfKYoEam3URCvaflABQAS+HBeg3/nRtK24FcwrkAmOaufBaXA3+p52whsJKCsLglFgk6jPmqgaCEQsrCB6eAVB8bZhmLbJi+77jrjRXbxE+chHlGh1ikxWG+9IbXjR6w2MHJodGJ59RXIvPC9znWfRbxmUjtdAVq2zrc1HQdmtD6s7u87uUfkypG1nBvMkYTlkZIzheqvQhJfKBuKJujBV3iKzIi0DcoPaeFlH1yuHc4HoVYAkSJPu84k/sUc73qm7fUP2rt9/9HSMXALM/p1qccNUskSO37wkeTP9N73jFXXd91eEy6nN9p8aXPrRu3atK5eqta45P7l5Vnf7Q2Or+Jyf/dfWw3EV1yqRdjWc/zjGo/Sn5XOAT9CHIKObSH1Baiqxgnseq7L8pUW9ICvq1jYl8MmehO7wX8A4AuYErJ1yaLT4gtH5ZffwPNjTG98hNHvKnvzD/8y7Be0FXBqmdEWPgPygxVlAe9BV96UpSdnl+t1P23sfkAXHCeIQuUyd0uZtl1eJ8LGYOcx5kDGWqeaJimS3gL/MS8BLwEvAS8BLwErikEvCExSUVv3+4l4CXgJfAsxJoW1IsFgmLVpK5LWLXIICHBWtlMcsCn91/r1AioCLgOwt2Fs/8BsnB4p3z+9r/AxpbnAuAtE43Bc85wqK9exG3ECSCZyKfzyhBRnSSF7ZLGCCSegK0A0zgHogDOJFzgByAm4BzgFWAb50kBaBBrOdedm6z2vVY0Y82adGyQGjLDUCJ7+iOxU/hHIAI8kKf+M7v6B8y5XpziYNe8jufRhjwToKO0hbIFUKJdgT0Wex/6R6dA2A1sq6zvtamnAOIJfEc/JQDKlFOQG58eHMAUgN40Ucs1ghl5dmA46vrYb7Q35y+Zibu2ayA26f4grq9dk99Z/++LWGcNUaSgZk9G7esahaioQP5dcQk6Cxb6zuxKnYoEPZEbe1jT1Zuvk5Bmhe8j+2vXbtxuLGp9u3ZVzQe/f6XtoDu934YvKnrwb3xez/8W6l8ycQ00kBvIc3XZhv7K+7xh9KhfpWhMOLivWtyY9+8tvS1Vyo+xktwaNNxrFUZfmEmLDa/0nPL5293D+3Z1Bh9SHEbkBGg4MIjdr8Z3epuV1yAd6bD6jOpqzS/JlAwaQG3f670M0o/oQR4ByDcbWcy18o6wP3vSn+mBOgH6WWxUAygtmfTHhAU6MWblF6/hDwgJSETCXQLUctYR55zkDqL72m7foGAYxwgTyKis/sdoP2NSgb8c2vLjz7khWQjX0fj7rrw8KdmwtKxQrPRuy+//icX5y+3QYCrg3eP/TRyGVMZFhBNsrBwc9VGLEO6eK7WcI0kHZieqQ3ILCYKRYrUms3RciG3KY7CchRHPbV4a2Gq8IsjYaEZ5qO5qag58rWh2U/+cj45ekuQNQXIdh2+UUKsTAA+ac+vvXDuqekHStfiNpA5hLoDEHc7cHFDfwTMb1lPqQ4tnWwTe3ylH9Kn2BlPe+NXn34PeUGbtQ6CaRfqDdc/NSvSwgyFFj5ydM3A6m+/aLdiPYSTPbNzI7ueOjL5qnc+trjdlpyj2u0JCcP8B3kGaUF5Xr1E/dARiNc7lb7cLj96YNZ37OAHDG+RXiKqdoiw3PVEYcuN+/Mbjh3OreY5Cw7pB+TrP6rffUGfkHCMK5WfeMtXOss9I/mR9zH1n/VZzY0GSerKxerPCi/vv2ZbzT1fVlnfLS3EpStxIVcZLKyaLZZ+fN3w+K6nr9/84d2PHvyqCAt0nufwjOeixQU6RP9iXEAvsRDqdvx/OsncQeIe9O10geUhD7C+wMIA8hoSsxsRgjXHXbJiC0VY5IpZ/YgszdANdIgxp9uB4Rc6g6s09Jw+AkHKnHaKNdUSeXQ7zVhHn6QdcfeJ26p9SkZcLIgB0yUD5lnmOnMBxRzdslj0ZMVZtIK/1EvAS8BLwEvAS8BL4JJKwBMWl1T8/uFeAl4CXgKnlQAgkxEWLJwBSlkUA74CoLBIZ5c5i3xzgQAwA7DCgpnrAQwBC1n8sqMZlAgQlh3nABu2cxUQzawrtPn1Wbc4l3sbiegxssXAaxb5AGz8P6a6sFO8tXNWYBZyuk5EA8Dol/Q/ZMakBcXW/8h2QP8DhnA9QMWTS/h+vyrICmv/tk5gbXHShY1+47u5wUK2kAF8ch75AJJABNAmAJjorREBgHWQZsgaUgFgGXAUnUZ/f5AmUEJXuYf70WVAZNoN3/bELll8PGvO8OwvADi2tx1LIwgrANYd7WfSN1ogX4f/fUAhngnptUZcxKZH+m6uPDB46wJfNrJESF5fusvt7nny/2fvPeAku8oz75sqdk4zPVEThHJAAkSSiDZgjJe89oexzYLtD3vXBhvnsNhrFgdgjdPnBBivwWCTM8YCRBYKSEJCaVJP7OkcKlfd8D3/23Va1dXVPUEz0ox0z+93uqpvPOc97zm37vO8oaeR9dyg4R4bjeYG99mbO5IV9EkJrv+tx6oc6rMXv7glc/BHD9d2vqW1E8o98fxi0Lu1WOklZFIMDv/eazHyXV1EZJhcImWB3BkFteoOoyjt17rdSwOvL+Vlf1C27bsWwk3RwdKTvVLQ++mn9X/xuSm79j/bryaA9YUzXs+XZNldu754T/2S2mEskyEVCHfSXp6qUfm8clv8ilp4h/IFLAb3aQzrywmZscYnTJsBw9dKboyuvEkVjxfGAbCXfjNmpVufeql123WXoFMQS5CyVzev21Ee2gg4+f+pAq4jO65T7hTrv7kesB6iT3j/XK8K6cC6uZYHjwGd36mx/95oYza60j5QvDe7fbeA6n7JsJNO/n6zPZ9S2JlJtWXF2uGHUT4Mw4FiuTGqtDHbwjAaKdYamwI/DOt+UCunG1vyuVSQct2a49qFdMo9LjJjv7wujtnZn3gw9KsTo+UPHXctX+uVLaJlTTz/x9WOPoWuym+rT92zJ7PFF9mCXMnt0Kn8tjYC5AO6s45Smc9mnjAukAPMOTwRIJJYQ7lPx+IIlO8uVix5T9wpcmLb+Oah1mTK8TmVfAZr9oNK1H3D7HW9X333XZdAkpwskc67DSQFXji4KKxFVJj2wQRCUN+kCtjMejamyrwyOTG4d6nsZJy7crvrymeyb19m08VKxo6n0KoiHYCEM2Q3z6HaL/zVJ6Jf+NlVh7LmIFOe5YeZR/JZ+nZ02HqjNRk+7/JtY1ZqZ2DdngcPX1kUNsv6xg1XP2nD/FyPI6+ci+85FMkbZU+63ojzsZzLYaI0B9q7gx5BVPyY6nNUAegpjAv6ZUhi5jRhLdFBCE7+Z7xORNDwu4fnyCdV0Xf0cxXZrXH7P3Nez03KU3OoO6zck49qPIPWIivwVqJCKHxZFZITsvzhEBWtXhV4d/BMfJ4qZEqncFZNMS1/GKICnWYNYz1FRjFJmpAV7eJK/k8kkEggkUAigUQCiQTOZQkkhMW5PDpJ2xIJJBJ4PEsAEM+E2DDWvwB/rNuAwlgRA6jwgkzlWABgXux5mceaEJJjTJUXeuIwQ2YACHNtrgNIYsDn5fAa5yFZgZ4gC/Oyb8DAGMTAc0V9ir83iQfIirgYYqLlf8AeY2XP/uVjzTGP988W/Yh1RvKNk9yqGnKC7Ya84Dv7DYmBLkIcoH/oNaAK5wFQo7cQCeguBAbgCzoK8E14L0BRrgP5hG5/QxXS4VJVA4bjBQMAzSdWulwHnWduAAxyfwgIgMgdzfO4v7FMbg0zgz4xt+ZmU4Ppf93ymtqx7OYnLXh9o9oWF9cK6qq1+9MXeU9K3bqpkEr1j3cNbJIwnL6wVFsM855ATsiWSJa735cmhumo8YmKnT7iO17DStfn5xcGAOU6lTdo4/3Zj88fqL6ifwUgJ5LCEJl8xoC76ziB6zoAc72Vqt/leU5fLgwHc6FXKkducS5Khwvh9r79la2KvF//yLMHPz0lgB0yAhmZslttfIcsjD9yU8/Vey9oTB7MhbV/005k/jZVyILWAnnztxrNt7oXW990dlr7Gp+MZcn43KTKOsX4M1ZYNUMIrFUA5ShYEXNPiNejCqNjwtzRTuY5zM1qBPehqwLWIRNkg65Byq4Au5tW+FwL/WFdhCyBTGOdRM86kV7mDiS7wHqZcZvqCStH5Y2Svz+zTXpmM9YAqp0IgNdoO4D4AwJsaVeoMFHW2NG5dI9cKKoNv0dhoDbKDWHQD8LeSqU+GspzxbHtlMZTXkeRn82kG06g+RKFA/lctkvpTfLV9MWTY/2/Vyxmn3zfjsI7357yx9/nhBWFjgl/6SGRrPj2Io17KRM1akocnnas6HJ5gSzrdMuRzBfmxpgq32OPFwHvloD3OFSaKt5QkAKAyhAWkAPMu3WL1wjGd+4fx9r9wPRw36UKC9UOCnMtxhjyiXUBcnJdwkJjauYEawTtQo9YNzoV1hX6hkfXp1RZfwibY9Z/4wVjvMoshdDi/rHHlSr6ATnTycML8pFj0Vd0ahGvmjevLRHuFYgoZe4WooL1ObvHusfpjX44k6rXLjx65Ff9re5Fd7V5WpjLTfYPXLQlNfWHynXzm3Y9gixDrmldL87ncC6B1B2ICrrBswNdYs3gNw6kpPFqatclyDPWEuYPXgPLZEVr0vcOog51b0g3SAXk/HlVyKY4j09rKTi550jWJREWL5IX1YZ0FPPFnEdIJlP4XYBXGNfE2w+ZV/V7YV3i5AR5KmgL88joOZ47eHlBfp2ooM94lDFXGHfWGYgKM4fbQ6ad6HrJ/kQCiQQSCSQSSCSQSCCRwKMugYSweNSHIGlAIoFEAokEVkmAF3hDWGCtyss7scYBB/nkZZ0XUwA3QF1eSnnJByDBA4OXVawIAW0A4jgO6zyuAyjDtQGoeAawj2sBCgbnIVkBYEQfTNJT5GWSwZo41oDqofq2Xmz8VYOQbDg5CUiuHIjnRfzZ1K8YhGt+5wC+mzBSBpAB7GHsAAENicYn+gyhAPDCPj4Bi9BrAExCfQFEEgIFsOi/qWIVjx4DJnMvgCzAL7wkDBAJkYXOMyfQF4gMQ36gN3EMeAA+AUvoCv/TnsKNIz9Umshs7ImIR99SAstNX+Tu+drOrge7x3IjvZO57q6Cm3MHgmJNILDfJCs4w1YomUJkOfdXbQewS9eJFucawwvlsIcE0CSHbQ/Jgxny76g6Ii0ikRbtgC19ib2JNAS9kn9aIYP2pVzbFdA9oP9TURgKBAs2Tlqp3mJkz6kzyubsLMyWLyzX+rr+I+sWsSA2hIVZUwCKh2t2auPneq87/qr5bzAWhrD4SGv/m99Za/5S0O277Kz1mfRPWDfXPxzLDlmNqZpwUCSiJb4NltTrFUBv6v2+536+q1S9XyGE+ord+Q1KH/4ybV+LrECGtPOm5idExSrr6yawzfjvUMWLgpAvgHuAhXhZtBe8feQFZEOk3ScdECHh+r47cm/KP4r8q31Kui6vGRKMmPBJgK+MnyHruCYW/5A2jP8/qEKGRYVSLVwsVjVkdrZRFzTtuVs0m4Y1r4ZTKXs2CMKKPGZsRYtKR1bDTbn49ITZMKx15zPeNpEb6Vw2f3im+9WFRteT7tm88O47+gqfudkNF5H3K1V/vr1DShb9Sunmi/Jh9baqnS5UnDTPivaC/JbX0md/9U73snsOME+QE/1DbyB4AFWNh0qHy6zYhJX7lxQa6lbP9++Sp4Uvdz4II8iVdnIBvTJhnch5gx7GpZlUu/XCBvQG4GZdQdarwnM1T2A8WTcAiPnEUn9Mlf4yXu3zzPzPWoUOYPnO8atCQWkb7USW5BogHNSCCZ+1Tkg3mmW/4yHjgcqv3/SU+91N0UyPVX2W24ju3lE4foFCUGWUN6O1z8vfj+0YsXbMT+S7jlT/U6pyi92I0DHCXH1Ea9nMOextwbjRKeYdBDZzYi3Ppq9o33+oQg5AbLPGnMizYllGTQ+diogLzn2vKuQHv5fIa7GijKcGuw6kR7vIU7OpMWOJ2GslK/jNBSnKPIA04Xok1T5VssIYixjvWNYkcqdACnOPN6p2mpftzcUjjWci7YAg4znJXGEenKxXUvs1k/8TCSQSSCSQSCCRQCKBRAKPugQSwuJRH4KkAYkEEgkkElghAV5ijacAL/IARACJgK18pwL4YRnMiy6W5bzoA54AwJjYx4QCYD8v9ZxrQipwLC+zgLmAO3zHqhRA/7x5uW2GgTKEC31CLsYqFpCS/rId2SGHks6hn77xttD3pJxBCTSJC67YqkeGyECv2wEdxgVAFHKA7yaXCsChsRRF1zkXAM6E9QAoZXzRdXT7ZqPD+gTUguQw3kiAXxB9ADmchw6wn7kF8GWSPHcCm7BazU5mNrhfH7rh+FRmJKq5mbI8Ko7KC6FPn1aPXfBfnPlcuZ4Pwsl0z2JGgegboTsiK11bnhR4ecQgrCzalVvG/qgEs1/nAiQCkIefn/lxZGVCm3TKIYAO0892so01wvyGU1/shu3YXWnPkVNFuKPhh7scxy7VZaFvRUFUtJ0eNWKHa4UH06F9vF7dGBQq2+rZ7vtF8EQmrE0rGkr8+H8/mhq2b+66tPq00n2QRsjjN1X/lD61FcYPbw3Wm7tFWvBJaJSyAFPAN9YZ+sn4QFpASPxih+ssb1IOg0uKPblLpkf6vtfwvC6RFYTyWquQUJccJcgJAsjEbF9xfDMEFGsnFv0A5YB86BdESCcvA86XNbbzdY3bsywlPg/t/H/Ylv9gLb1rsZS7Lhp4qslJcUfj3XftwGKfvgPMQ1gYS3HTjp9p7mf8P3NX4Y8XAv9nbCXb9mp+4MoPbLtVD6+MrKgrCqMBecwM1vywLoC/WyGg/Fo9iHw3iORNs7FUbVTKaa/c25Xxu/MpWx41Rd+7uF5oPLfWX/gUugFZh44Tcm05nIxylWgRdOW6ke3a6M9dpzE2ZG+rrCAXIToOdxUrlZ/+py9yPeRGZe4BMNO3F6t2Au5XyL35D/H0GRss5G9XEu7C5MaBjMaZeQ3A38kbAtKCXCh1Ac3C9K0pgGfp1YrSzFmE5xTeVpApq0ialhNYSz6jivcPnlfoZ6OZByk+bI2QRawpkG9cH2+ZToWcL6wlcYJjQ1ZwYGtIN5EXBqw24QyRr1kDrXc859bwGWP/OP3U7IduzGaKc6OLswvPz9zxU/fkdqQOpldHBproH7DuvOYJ1uWjBzKjD8zckJpo3KCV8fvkxtB1v9jMlcFady7mMED/mNsQScbLql22rD+QkQdV0Wm8mMzzfo2hWHMzcoCs2Kt1eZ/m9f+r76s8ZQjDVajlLOUssjYp77sbBeTBQVdMO/iNBbmO/p7ObyfWdfSA5xFEGPOUdfFXT7JDtIV1D9kgD9rF8w05JsYZJynE5LBEAokEEgkkEkgkkEjg3JVAQlicu2OTtCyRQCKBx58EjGcFPecFmJdoQ0zwHRAutvhWBYAlbAYACkAsgD0vsLwEs5/vgL5YfAK0mFA6Y/rOyyzX50U7BhZVT9pS8RwaFvoEyEr7eZ4BOCIX+gYZA5lD/+inkS1AXByDPSmPjATaPDBab4oeMi6QDgbAYz/jR0UnAYQAtAD/2cb4AhjyP0APeg9QY3KWQHYQOx7LWfSCYziee2G9y/UAizmOfcwVAB50Yhl0aoZRqQnoa7x3+xu8b224vlZxcnXHDq/XUeiVu8MZm7oidU+0NXXoCWmrsj+0nbFcWCfUzuZJr/+Shp2qCxADXGMO/qUs6PEO4R51k3g5+/F/Mt4nkCqATu3x/LGyJR/DfQI5WwE6QwDRfwBk6ki17rNeXCYAvL8RhkqN4G7Ih/X0bqc0ftzJDmStoK9PSWVzQsNrk9cfCtPHb3NSmfAAEAAAIABJREFUC+9VpCrCT7UWZEbs9OPfzV+yR4QF8wYw7B+bbQRU6/Qb8nXaDpAHOYGlbx3rbskRkJAKcUFeDKzPP636J6oQByuKYltZ1Vy6MjXSn/P84FqFDOLctQr3YxwhKrk2clwF2DVBbUB8wHHC+eCpgZU0/1NYKzoVkRDhscjOvkeEBffZ54Slcnf5G51i1aNjhBeClOnkNcP10Tv2XzdX23+LW5+rWkF3Xt4wWeWnkENFlFUMu7rjWFXHjlKikTMiLtxMWjm41RB5VCiJjL1RihRpjNONhvwuGmHddcNh37KLM9kXzmYGf3lsw8yfF5yoYohqE3LpdWKmhc57qgoMZqc6kRUkx/7J/rnid556873eyOQ8OmYSauOdxLgTeghCplNIpHYZEtqLOfk1VQBngF/k2Ljm9gcbNz/j8jF95xieZ4Rxai+s67/WPO+fRSYwf5bcuW5cXteZD+gW68CqBAnNCzL/0GMICzwr8FSsrJGfqL0NEIfoDusE7QHkbi+0CW8uAOQDauOJnjM8v5AtbWa+8d3k+LG+vePnykfSTyq+qv83bs1FC6ltlal6Jmy89OLakU3KMbPq5gcUqW67O2mN2AtWKiVNmIiuisrK5RHJSj+y/k4nMB/PJTAb3aHP6CDjAvGFZ0x7AcgfU0WH0B3G+XTJCgvdkQ4VlHtmn2tFucCy3308NdiRJOgKq9a8220NBgUrG4V/rfBpPGsgunh+8ByptRJdHdreaZMxSuF3GesPv9luUIXIJj/TyRRIP+ZMJbTdYmCn7jnee/nktvnbIaTOx99yJ9Pn5JhEAokEEgkkEkgkkEjgcSaBhLB4nA140t1EAokEznkJAGKYEAGATcTK5sWeF2Qqlq28kLJ+89IOMcF2Xvy/pYqFKWAQABNgPlarWJlzDtsAXQD0AC7YFgO154PXQTPkkBlAZASIRAUApG/m5d/EbTbx8wEvqbHcdJ3Ey8JI8RH8bPHAaL2rIQmMJ0b7PkDo2ANIlXlgQkaZvAbMAfYzHwCAsCjmOzoAEAiYzX72QTQQpojrYAGPTpjrx+Gr2ucB4E/2478Z7Xb2Z3bZ+xvHos2ZYtTVm7Wrhd3evmije7w26h0NCyn3wqrjZAp2DovtexVKJCfLXULy3KRPADlDIAatyYMJ86RwT8ab5AM6juTTreWNauwXRsIaxAdtRe+RgdF/zu2WN0XDc+xFWeBfo53bldd4KIgsT4Ccm4sCf1tYZd5TUhkr7C3a3vBCbdPYxtK2Sbuv/AnbrrUTFhxLOCrWnz9S/P7JN019gjFgbSHmP3MN0LaVaGId2qH6TtV3qf69AOU5AXp+M8wW1zShwmi3vE6UsHspJwU285AIs6HjDBZ6c9bUyEDu/ssusI5uHWaBMsB7sxvLH4Rg+roq8kH2R9uB4pZ8FXjrALhD8vK9zU4/XkdaC+sHwCBr5f2Rk52K7LTv+ZOA3GuBgmyHtCBGPiHLIFBIXN1efl8bXmvbwcaaXzrsBLm0vGM2KKqaKz6iohwVw47nSrZ2w3XtnOOKX4isYiOIyr4f9ElTs9mM5/hiLKqNRrZS9+qaSF5k+1E+0+UcH/ot7jcxOv12dP2DqpAyAPSvq9gZ67g3YIlUsx7MwJOtLIon9i89C6Xqs266c9vo+MyoPCEA05EV8wi94/vJeFX8p477a1XOhzQeU2XeMTcDk1vh3b8UE0VfbsoLvYG46FT+uzYCun9LgHOtZR6hg8x5PCz+XLU1fE/rdQCbWQ8gTpiP5XawuYNnBdcGUIakwBOpYwih5k24LveIQwSt0Qer6V1hvANZkwxhQfvNvGaeZA7Vrw0+MPt31Zf1/+43B92x/Rqb+6R5PyMA/dpZd3UOewHv1tDoouUNi+X6QdUKkXbR+hllGZrTee/U7MuIPDRk8COahLlNtmYNY21kbaa/r1Btn4Nj2ga5RE/QEUiCFWTFCXJXrBqGeD2Y+gTyz8y53elpr++T33CvnK7aqT/Suu3igWTKHbkLrWsre6y5oOeBDdF8xYl8vLji0IHUUyQrjNEEfaZiVAFpyiT8n6qQMVeupTfxdtvlmZIN3dRXq17PxyvpocJc1wX1o4NPrtwy8rK44W97zjLhv+JSrR4+694j2ZlIIJFAIoFEAokEEgkkEjhHJJAQFufIQCTNSCSQSODxK4EmEG+s7kx4I8gGwC/ADwA2gFjMKnnJBTiCdDBAHYAQVsqAUgB7vPTz8jqmal6SeclmGyE2AGAAbgBAKacTzuDRHDATMotnGJX2Y4UJaYMlNp4oALStFvQA3CYZ96PZ9uTea0igA6ERA1OaHwYUZz7wHb0FADXeNBwGcI1uUwDOscI1ZBbgIboBMAZoy3aAQfSBukyadGray1OfUg7c4uixaNNlk9GGuE3VKNvz/eCqBc9tfHMmk7vEc6sDDTudC2x30bcUfd6y71UFYOPeANjUFWRFy72M9wd6u6qocb2zTgp0kn4bzyvmPCRdPKflMLHBj6zBMAovFHkh6317QA2tK/eBowmSkqdHPW1F+ZrlHPUth/+tSpS9rTH5zAXbrdzh9ez7S3lZ/HKH2xMqiVA+xmuBtmJFjhw/qQrhYEJKQWJQkDMgPYD91wUQLnSwYqcfkB+EzoFoAOB/ucI+XVfLpHZObRi4Ynaw1yp25yArOomFbdVUw/9reWPcqfNYzwjBs2KON8kKwEFkdYHqk1UBxIkV315YIw1g+jF95388QYibP+8G88ZrI+qQQ8EiTFETRCd8kSGEAe2frUqOofbyRGU2OWZ375mO5ocV8clWTChnVpH5ZkNZfrtKmh4G0UbHVainRuAt1qubvZRXchynqhwW4jSiUI4olh9EfaWyv7FU8afkkeFnhnsapUo9EmkRiLBAX5ENxMuwANkHF938RQJprX3plfmMlVzYV/ibhd3Hj01v/cHEdRsnZq8QWYG3CDH1eQbh/QBwT2U9NR5urf0i5BPPKqzhyXfCs4ZrsD6jQ9V2C3C8jSQvCATWbkLcrEVYXKV9WMKPqR7/zncurVml+5jXtI1nI3kwDFmBHrQmVCZUlwlJdkxjtZ7HTmt/eL4QrgcLeKzfO4Wt4njmCJ5UeFdQO4bkaZIVxiABXYOkYIyYD8xxnluGaEWO1Un/wuP/MP1v4jZ/e9/mru982ImixY2NuVeIsPix1obyXXkurHFv0Hp28fvW1oumxH4pPzuaWLHerKv2qlX/S3QY48C64Yu8WDUe7dc8S/8jV8YNTyOMLMjtAnHZXszvnHjNKd79O+YZEB8nEP6Ufrs089cYAiqlXENPU/4Zb9hf7DmSGna/0X2lYmOubML+9KYgE/pH5G1xrD8osp6Hp0hUWJIz96TP6CsksAnJyZoJyUYxnl6rpWA7k1oHPxGmuz4S2un+Sm5k4vu7fmZmcvjJdsEd8CpWyss0AnG9dlipNoyMolOVz1ka6+SyiQQSCSQSSCSQSCCRQCKB05JAQlicltiSkxIJJBJIJHBWJGBIC17CAV0hHwDbADH4DujCyz0eE4AcvAQ/V5WXaF78OcZYjXMOIB1WwoC5fHJ8DBqpAjjhaXDaoRXOigRO7qImZBBH852+AFQBpNFHZAcgADiAHAizg2UmQBBAVVUgeP188Co5OXE8to8yuVVaXDDQWRNOyhByjC+kAL9rTExxjjEANnoPKMq5gP3oiQmFxjHkcFllNS/vB6fX+pfBDc5U/buNp1wjEmJ0wJ7bU7S6R7u9+UMXd3+vkbHroa0458oLMKD9JPol5MwfqEIwMDexCi8bi3Bds33A0GHjEUKoK7wAlovCkLzajazCzd7AjU/z54x3Ff0E4ES3N0s2O3URgNUryX1ODgR9H1VoH4URcvyU4O1RJWku2G6/kEo7HwYL/VHjwjAYuC8sbytZPfvJLUHbARFbC2sN8fr3ysviMH0Q6EefIISQJ9b7hrBoPQ8ZYzENiOvqHOYkiWlbAUa+lwTmMX9Lpa7sV0rduVAkxZGDF2zcGXhu1/xAu8H1Q7fYfHT6Lh2zwQ7D4vFNQytyVrSECmKc6RNWzICDr1ddKxcGN4M8wVPtfaroB/2MPQLa8ya0yWnFv82wM3E+D1U8UjoRFgpzZLtO15752vS1YuXSQTbrKT+FXW3UA1+5SCpyssh5jjtje06/r9g1aU/JvoPQq9R8V9TdQFcmrRQXYa0RBBcql8WiAMtavRHEeYu69ORoypsxm1WSbamS9da67T1FFvq/KoJC8ZAeSrEhEst7evneIYG3r8qkauPiifAOQY/e2qGvHUNJNcebOUkbCP/ENfjOMycG5jXeq8tffcL/2196OXMUYuUnVclBwbOuXR/JmXGzOvKFtEBkETC9bhQyroD7kAqmtJIV/6qNjCcEmglNtqoNa3hXoBPXqjLvWCdWu6Qs5XQh8THzHU+A5bneoacQBciO9sIYMU8MkM0zCzIVeTG3WccoGC8c+/j8H5de67xxdlPm+5++oD6xV4SFP+d1v1BhvbjGchEhZd2b3W4pCbzVd2XJUkg1K5rQijBjvT48IhnVpd+hiMIotui/TeMBcbjs8dKhzWd6EzJg3WLdgASCCIOMai94E8zKSey7YXXD3sbsNcgfhTVryOmEPuI3AbInVwbyHZUu/VqfpowS0CurfcP6Yu9K3kTh0w7fkdt97IHs1kV5X4Svu/ZLp0SSSL7MB0gK+olnEmPMukBOlsvXES5z5oOR48IxK/hb/lBp9Jrx6dGnHRgffWa62rujJ6jYeVcrR79jz8/Lv67hB0E65XpaA7hnXQRZ7FmaEBdnWoWT6yUSSCSQSCCRQCKBRAKPhAQSwuKRkHJyj0QCiQQSCZycBHgBNwQCL5q85BICCtAQ4ASrZixXeXHH8wKLcixLQUABljgfEJHzAD0BBuJQN6qAQbysUzjehEg6uZadW0eZcBL0GRnEoK0qwA4v+YRZAJQAGEAmAFoGMDNhdc6tHiWtOVUJGNKq1R6WsTUEBr9vGHuOi8N/NOeC8aoAdI8B1PVIu9/N/KlXjnI7f9T74oV3B1f6PwgvtbZ7B28JvOiaTZnDF0Up/9Ij7ka7y13kPnh8AILhLUB8cazK43nWGgaqQ0eNtwHJw9HdZUgXhFlhna7MW0F/2XbRd5NLgusCvu5QHdIFNju2vVXERY++pxQOKqfO5+RRwZxXAvDQT4uTUdJtcO9sRgkTFBuN+eI25i8tp4Zv/rLtlQEPSRrcXvBKoEJ6VgmHJACc+cR6BJgPMfGHqu3hTH5K22jzv6niSWEIoxXXx+JeYHGQqTVmc+VaadP4TPXArs2en3oITG89oatUtS6+75A1OLOQOrhz0/euve2BcHAmlr/MyJfzGgBYsyYAhBIXHwCY9q6XuJs4/4Da6AVW8uiTyfHTQSzrbyLhsvrFWqvE5jFI/QerzoisX7HTM/N2bvxLYX1bVKn4m+RRsSEMIyf0o65QjEXaC4dEUmhco2y5UkeP69pf9xtRKgBhlc4p8cViuVqfFpFRzKa9+qaRHrPux3Kpf9gK73zeroXsQOPuRsp78kRmYC4VBQMokyk1O2UVnLw10Ffc1jVc2+bko+tEMx05Sf875PUeVcgBvAboN+Mdh3Mz4Z/Wldh7YnkxZ0iITeg2Qk+RuwJFAMw35c2ZsH7XBn9uWAByTTrNmP5Vcyfgu4mVBFGIXqILXJfxLJ2kdTzPTmSN/CBDydmxyqOheU9DiuLJUtG4dwTSBR5zzZTykXRr/CAXR7VYZbX+KNeM2CPaHUXMZWRm9NV4XLL/qMJDMWRzP7n9JbcqV86fi3Q6JI+L11SdtAn5FjdpX2azdU1ln1V0claPV7a8zSItNCpRLc539aKoIOIiij1O0BNIlhkB6+Z3QYuoH/qqMTxThfWY3yfMTXSlE1mBX8gHtDqr4fZsUBltNGafaOS6LgDfyftJ1+K5wG8oCAJkhaGHacNyXDvW23xYU0J6xL5USk52hz52iM7gN8UbpaNj663nTYKCUxlv9AdCCU+1lzS3oUeQRaz1axUI2DcpZ862yMuW/d7Nhwrbrp8av+a/1aZS271i1R+qB3ZezQyzocJ/pbx8PQjr1Zq9qHVhgfVDa4Z5NrZ6Ea5zy2RXIoFEAokEEgkkEkgkkEjg3JJAQlicW+ORtCaRQCKBx68EeLkEXDR5GABXeOHlxR3ABuLCWJZjmQlQzwu8yV8BSQGYwT6+A7J8tXkMIAVgKpXjz0evilbNMC/iyAUQAhkBtgB+GBkCHANyARgAOhr5AlYgA2TXite1Xj/5fg5K4AQ5MAgdZfSasTY5LwBrmEdUtpvwK4bMWLenH2682n6R96XLD4bbR/vs+XsDy+k7Gm5+hmDiwZxbchph5lg+qt7WG5aOCRw8Ii8LQDDICnTTN8m1W2+i2C5WBy8L2gX4P2aONUougmGnyIWF4pI1PH+MdwiHQAiwZuTV/17lNhD2aWWk9F1yGcl42iDnCp0QiTlRBuco0rbIEwGibSEeWKNRo69R2f/acm73P4sTqRHCCOKitRASCGv3r5vcAYC+AgZNiCpIDpKDf0gVILa1QGbQTtajSc7pkDcA4mSDQkE9U/XVC/3dO2U0/BBi2HK1wdlF66o791l988VweGr+CTv3j/+uGwQArpAN38NbI9Jst7vjdZD+MfchKgC+CQm1VvmCdkAsAHgDDrNGQAh1DO2zznXadzGueBoQMugPVp2nxBSWW31lZviO7/vHRwtRmF50bXvGkVtFox6m5WWRVoptcFTh0nZF/1va19CP92NS4EKl1lAkKUvBYCJIDF9jH+RzoqfQgiVvhthrb2a4L1u0c1v25Ta/XITF8wvpPGvlirK7Nm5dWj0UW+a7G0MrvEAXu1ceBVxp7SfG17T3X1RZgwFhzVochxA7KaKipRXN8FCMGZ4ZEGSMB3kwWstgxcl86r7s9s/3l0qXeVGwgxBnzWLIChIYv1YVHWCu75Penex6j8wgmHhu7lAlfFinPCTcEgMCiBEIm9gTp62t8b+tZIX+HRAPBbFI23K6Wa+j5ChBFHny0JKxvDWr0StrPvMcp/+0nzkfj6Vq9MFDn62PXv7798i7Yndo2XjvrCAsuOcX5ClwbXlPnDB6W2Packkv3aPc0RPyRORqvn5TBBak4p+pEvYMUgddZV6fjvdCp663bzPEAfLlXu05e8zx5LeZ15J1l2X7s6nBO/xff+7/PCXPhuaFDIFtSC+8MCEyCb+0HBMN/ZEeWRv8eevppXutL/d0TNHCGoZuWh28cQgHR+gnxsd4zGBogqT55L4YlxgPHcgKdKedQMXDjvUMndqqgH4PhunuB+cveO7EsSe+IVPp2zFSLza6Ko3GoLwpvJ4upVQSoy2Pit5qJbCU7ybo6U3XZheCQIQF9+Z3kCf9C+Rlcb7/7jsZ/UqOSSSQSCCRQCKBRAKJBB5DEkgIi8fQYCZdSSSQSOC8lYABIgDueMkEhI8tMFV5QeYF1uRgAFTgxROvAkASwELergE3DFgDQMcLL6AD2wBSOM94cMSfJtTOeSY1A0DQbGNlTv+QFWQF3wGakBFgD8QO/wPqGk8UZErybRmlrw4DdLryaEsKbi5jcOf2yy6DL2sA8afbjOS8JZKK8Tegm7E2Rzatcl8XACOs0NNLxexxpRH4d/+VOx4ILrratYKR2WB0a8quL2Sd8h1pr9wrL4ueRTu/ILARAI45ub+ph2uCfpAWbUXJveeZ5wBWKwoKpNhtT5Mx7W2zdqoyGDUAxQyIaUhMtvUueVjYeVXBWAokwmFCPwXIyX6esFdCvLVWpKPoSl2X/nNeLQryx3QQtyIHQTthQXsARQkbFYd2YkPT0wJwEyCPbYRTaicsOPTlqlgMMx/3SK7LVu4C/ljzWMsgZJm/V4msWJ1NWDs2Hp+1du89ZuFhkavUHIW66VGOBRNq6WqtnD9m5xWz5QErdK8QWZnS2unE9ySh+HpkBV4BjB3yB3BnfaA+bNC2GRrK5CQgVj05P1YUReW7KsoefqGXP/bRsLyT8Rd2HYfqG9BoZZSz4rjtRBvCeiTrfLuuAVOaFEdUVDTo+1FZFvtBPuNku3LpoVzWm+rz6unRG9/qb/v+e5c8aFJe19xAz+aJjQOXFvO5GxRGa4Vlt/JWWJv8WWujP6fM3qK4pBZURyMZjukKuqEs8luh+Jv0HyFtGK//q0qb6WMcZtDUUyUrjFBaZIZeAaTzjIM0W1GUMPx5mxsz2Z31iTicT0vBOwMCC3CYNZ/5uGYS7PbrNvsFqI0VPu9JncJ5cRrXRBZfb96nupbl/VB/3hHAnBOxNKBgX5vlRbNRsb0UYs5yFbYtazm274R2VQC9BtZqaEgqUj5kOqU5zfwg5COjgEwovghSDBBu1FjNqf61Rm1FuCp5Bljf7L7C2iH5EP4LMN7bLdJCPQoV6EzEhZBuXSFQ7o8ofk6i/xA9GDowD850YX1BJ2nns1X/R4cbmLBaX9Y+km0bUvSEbengWcH9+D0FOcLz//mq/BYg10krwYPe5uSpY/UGZYVXKn5K5MVTRD6jA60FPbhelbBlyH5FvhyRFSZMH+cRyux5qsw1yBL6204qtXtYoLfInnG+LfIyt9aGL5499oy3RLMbnpKZs3t6nFqwVTqS1VLdJT1JFYr1LX4YlEVcRBmtAfVG1KccFkUt+bWU501l0s54sVynf7ZIiyQ01Am1KDkgkUAigUQCiQQSCSQSOJckkBAW59JoJG1JJJBI4DEtgXUAbWMBbhL0EkJghyohJoihDggECQGIRfgEABxewHnx52XchL/hBZqXfHJdGEtGXlYB3+JkkU0Bn69kBc1v9a7ACjuO1a8KQMA+wE7AF5OUGSQL+VCRGcCpAbDXIhOaYnrYH4aIMu0242Ss+814nI7l6MNu3GPtAh2In1a5nrKMP9Z4mfN896veN4JnCOrrv2Q8Gr0wayv9CW4MlhN0eYuHqlF+SF4XmqcRcxVgEdAJy9n14tjHom/zskBX0FVCEsUAGsewMMTKo7sOh/WsXCBKIizYZMKf8Q96vVlG9QKx7Jw6mlIE84zyXqhZ5NZQFgsRGK48UERUKIAIhGjE3IFcoN17Iz+fCiuj427XQazZsW7+R9VW4oA59eOqBwjbY4DZpqcF7QUYJvTThaqdQp2Qk+BzqgCucUgp5cSgzxCtWDqzlgHwdSQr+ueKH91+cGKhu1h+Q+9CyeoulMVMtAypbV0kIPZddp/1LYGwC4rVP+HsiPtnEto2Jbnig7X1/ar3qeIdAKkbJ0dHcp1OOJ1tLfksPtDs56tXXke3csrPtbKHPtIobJ71/fSo57l1DXpJPNPRqsI8SbezOmrAkfeMclbYYi66U2mnaltuzbbCosDWo2mrXu4uTdR33/ceq//+f9upe7AuIt+unkK5a8uRqZn9uzeH9UyKNXO5DE8tWBdVj1h9fWWrO6zgyhHvk5eK5SrqfiRoVrbac3qCvE7ExS49RfAMuEWV5xDALXqLN8XDJnhMo1pIC7ws/l6K8kK16qWt7RagnN2T2RKD8Tvrx5UoRb4GS8MGuE84KeYh4aVo48m0jekGuIwOQnABlhMKivxIeNu0yg3yDhlAVqA3PF876gyJtjUFM7btdCuvereU60K5wFwu0Jl569murTwN8Zz0NO5FEYwK4BTm1Z2jGgp0mHtDJgCE8yyHNLQJPcVc1Hp0u/r9ToHsz5NMyM2wXKCeJrwBa0HR5JRcWmSFQszJJ8ORdvhKYw0tpvHNqb5eWs+z8Z9VGc+bmjKrnS7x1NoOtdOQFegkIdqo6FFroW/vasqSsXs485D7MZbIDO8wQkFBXLKOUSn0E9KNSnis6zSAby+6uWOSZU8HwoK17S9V/7cqa9kR9LTpxWTWMojXHaqEgOI7BMnK7PYP9dgs72yBAPwTVQgjdGlm+vq3lOav+Wl3Lsz1lv3Ulkqpvl0Dtknh34Yq9UZKxESfYzsjarPtuY05KVk5nbL7u3PpGdtxZup1XxPCLvV0p2siNriXn5AWDwk/+ZZIIJFAIoFEAokEEgmc+xJICItzf4ySFiYSSCTw2JeAsZhuDf0A+AEASuHFG9AFwOQGVcgLclgARj1RFdCRwvGQGwCIgAGs8Ybo4Hts/XqeelYYLYhhWFVe6gFt6atJUA7QhKwAY5EX4Cj/c7wJh4D1IvtN0mZz3TP52RqGArkbsIbvgE8ULD/jZM8ishh3kj6fyTYk13qYErgvvCT6rP/iTePRhsu2pg5P99lzAJPOkDNVLYdd1Xl/cC7vFpTnOESXTE4HvAxOSFbQtDYvi6hJYOChgQXvC1BaFKPpYZE97OQ290XiTpb0Br1Gp5kH3HsSC2vYFHkoxNCtLPBjW3lKE0nlPB+DeVVjDWzCqLn+/OVFERbMD0DSduKAECqsL+9VpQ3LJu1N0gK9Jrk0683bVJ/eQfxEwSdE1L2yDqdJtAFAD3CdkFKAmJ3K3ZV85tuTGweObTs0GfYslja7Qfij8YFNG2qblSBvvSSqWD8sGPjzav02SahTXBdkwNwbU/2YKgnSISwYN/pwtsKmoCOsR4RPAjwlAe9S0TjZjn9xlD8wYmd3lMPylmPiJOIwWVoaKkFgy9o9VCQox/HSgrxDZSJQdC8px1Tare/1GmW7b2EsHIpmy12V8Vr+/i/sdBplEqhfHTq2pzBbV6kWtx6eOnT31buf1S7gzcemrc3jU1ZwiWd5Sn3REl7JEukTF6eoHEg1a2twwPqGvC4qWj0PCMg+2RBL7bc8qf+bpEVJhMQXcmFtouakt1TtFLlUlstBpRXAk0D5OKwtjWk/FfkQHHgJMYduUuXZ2DhR3goB6oaoAMxG93m+kn35aaoQW01JxLeGVDTeVHxCjhP+bVW/ICv6erJerRZ0yW2mJ5Nyhup+sFVj2ZvOeMdrNX+jkqyzr0uh2jKuJ8LRV3g32x6R74Wn0F7T8rKZkprv1YOCduF92ZphM0wqAAAgAElEQVRXBb3Cu+vOZji6VW0gH4NCR0ldbEsyXPJGYQGQJCP5I1ID0ayaOyMa1zdosSAZNuQjIPotAuSnNNanPS+aZAXPXBNi65X6jrdDe8E7kvWFXDgQFqfiFWOuZYwEMPqAiDCGDMxzwi+1PmRNTi+2vV/1g/riD/mLD2SjxvuVs4IcLK9raySEC54S6ZHJeU+yYYmOiSdVCA0MSnhOQNqu0NXmddqJL9b7f1dF//iOvi5OPee3rdKO653F9IgzM1u0G/VqerHcEOcc5rWyD1RrwXDgR+nQDvqDyA49T2ogrwqdm1GDhlMpt6aQUJ68eBRazCoqEbcycgfmd2a73JP/EwkkEkgkkEggkUAigUQC56QEEsLinByWpFGJBBIJPI4kYF6weWEFpKKatZmXXl7yAQEBKkxYFYgKXugBFK5Q5QUZwO1HVAFcABwBBLEQ5cUdUMMk1DxjlsOP4hghK0oc6qDZfyy0AXTuUAUoIOYO8gGwQKaEyNqhCkALMIIczhZDYKw7kT2V+3M/xgHAlPHFgp52sC0Gn5vEhSFkml1UIxMiY1kWj+SXf4x+2qtaXaP9qVn/4u47Zm4vPbNQ8nuGtmYPzFejbHRNz82X9bgLgPiEL8HaGkCapLsnNcc6eFgAoKEXJN9+gekrKFPdcl446WRuioICoJTRe9YEiIMZgZFzgporunFNx8fOFQCUpLCI6QtxF0v/Rb4+AQ+Jq44eQmzG+qmktkFmy+dNUm9IQIC41oLFMCVDLgvOMTv/Qt/fNPUJSEIslf+XKjkh2gtA398o7NAfTqT6jyhp8Ia67e0S2Pqr2o5Fuylj+gJYiVX5H6sqrJEbbT46fbvCQhHeh5AuB9S9ncwcZXhYYna02skrYNwZtl7uMOs7F8gKPB0AtfEkIdcC9yueCNRe84onsaOZmwEw/Wuqf6gKINwszdHKTPxCZuj7/xBGI8fsICX/Ebs/UA4Lz4n8hh8u+FZ0xPLDjJJxCz0Oq07dn+izJjbn/MXClslvXTI8c+fu3tn7i+lGoVtj/kyB3pcoHNTAkW0b7L0XbR0+tmVoR6em+p5rHesZsgaPFSx3m3Dp2LdnZZFcLxRd/tNen1WMLrI+2/h8DI6e9SKdCsdTgxUlBLcPp0fu+V7uCatA4Gk1SsdYPWFZfEvl75SH3DwfWfNXxIrq1GDpMjqBxkAkISPIJAg6SDd0uj3fB88YwGx0fa/qunlO0inHKcltRrkpugUi79Z03KKx3BjUGluCUM0OlcjeDvs1m7LKQjKu9d4TO4WH1KiYxX2+TOoJJaX9KApzddkyv8V7h3ZAvL1P9fXt/byp+yoROxnFECvYFzQmLRFA8SG2Zj81ZBbQ05o1EJXV38i6RP/9jmqcQ0vAPLrbGmZvlSg7JeWWbGkrz0BCenFN5m8nsoLrAdbjjcBn7Im16ibrb+C5y5rG/VgbWcMglzDqIAdJp+c9awwh4W5VnYasy4X1GZE85FBBjyBYW9dBrv9m1X9wwjBbT6dS6XoDnUSgEK4QhTwT2sNJmZajaxRkCRH2LdXPq0JWoFMFPJXueOtv09Zo/MisXa400gonltEa0CfzBvnHiJtUGDGRW9UgkP5EwWCtHvm5lEfC9uONul9VrMvBXCY1ZaW9SiMIArdhz0ivpmt1/+Hm5DH9SD4TCSQSSCSQSCCRQCKBRAJnXQIJYXHWRZzcIJFAIoFEAutKwBhSA1biQQHJYMIZ8eJuwkGwXgMrAMLzAg6shBXoRlXAel5EOQ9AHHCBF3ZAvzhGvSphoE4VADhXh85YwwIkAYJC6gDAIhM+KWwDSECGJrwH2zkHwNaEhjrTfTQE1JLN9xLYgUUscBCFbRArjCfbGH8zVowPYxZ7XpzphiXXO3kJiEzQOB5LC+XP9aZmiwOZqe3D9ePzc/5wTzXKFfu96S3VMNcQqPwdgVxY7wI+nZRnhWlFh+Tb6AQWusugEh4SoVSkbjvblIE2FHFhQDf0Az05LjpihHS6DZvcFVZKB+SZ9MZSfomZExSKF89DRB2HQE5QuZYJv8J6Qxgd1poPdpAYIZb+SJXE4ivA4KanBWvNbaqQp7+p+pzWa6itV/m28y9VO/02JWK4XP0DFG4lKzgcwA+w+auqY6ql0HEseVgAQBKG6K1a1fqVr+KJgm/foiTbl8PLOJrxzoXWDkV3X6/gBYJnhQLixGNG32tnk6xoaQz3Yu1i3WYdx5J8qcSj2ni2wkJ9ws4c3+sXL2i4jqMwQtFQ1rM3pMIG5EU258NrRo3Ay1b6w0JqcOGB9MjsXVs3zN99ba5weCjVKOYhqERWWAr9ZJW6stZCf5clUNUKXMPzPtQikpiXc1krmrKL3bPlKWVPALbH42V1sZV82rVukwfLnemf0Jr2ntOygF93cFp3KmwYOpqWxbt003Zk9b59xF+0/qOH3MVScoHueA9QFt08iT2mRYTVBvziRxTaCv1ZleDdXL9p9Y/Uee5CbtNnLvYa1We3tAPQurVAdJFXg/HDu2JFHoNOUpuaLac0ljnPc4bkTbFBMzjPtJalfJ/rRP2am5ONIFoC2pVoW2DznDwr9CyLBjX1BeDbaZ1XUEQ3kqozX9HbZe+DJmkB4A0R96XmPjyWVpRb8xfbF9aOycXStS6pHY6TTJviKa14IBpGQcjiItICYP0duj/kDPMZgg0Q3+RuOCEp25QxY8jz7lpViAoIu7UK4D1jwDN7Xe+dtnwVZk3kmcvvAeYZ5zN25M8Rn7qmcQJrFCE0Y+JXtdbzvIpCbXkIByMQ9j23rcGDIit+S7lgPqX5FWluQcaw7pGfxoSbWquPrGmEn2O8IZluUkVXSyIqlnXpmm290Y13H7d9P3SrddGTYrbkypdW7hOvXo+y0o+SvC1yjSAUOSmvCq3ucnvqkU5pUzjnuW4hnXYXXcftU8+n9X+QVqBAERZrSz/Zk0ggkUAigUQCiQQSCSQSOMckkBAW59iAJM1JJJBI4HEpAQMY8pIMUMBbJS+xAFvE4wZ8BywA/N6hCsACMA9ocUCVl3RICwA9gHhAGK4DsMGLdBxfW0WchWytz/9CH3i5N4QMPTLEDCEbTBgmvkNQIDcsaJGp8ayI5dwUypmUiSEsaJMJe8N32gqhwtjhWQF6SJsgKxhvLD053qCKa8ZEP/+H7/zogWMFXo+3kJpsbHr6rYvPssbr2wRqRQfLQdficOr4gVqY/ZZrA/PFHlCLJ+tZsU7vGXtANkjIuBhPCcciP4Xl1ZfcbQD14lBQIipqNdspar+ClEe1iuX2KviLcjTHQaFilK6p8IoHogVgaV0wOVRMgmTWCBN9ik+sm4mljpcExENrAXT8W9VWkm15f5O0APjDe+FPVfESi0lEQW6KzeMKZM7mR/25tw8GhTumvD7WNzzEAProPxbdtAEwmLUNEBLCb2bfhVsaxNMP/kmx/Wc1/3M61rY+E81bx51B6/mO8f9oa3D8b82aDies98ua/Ad2RnlGQs3BTExUnHaom063OcE2+kXILfoFuHnjQ8drlFiavbmftzd8dj5f/5HvDSzY/bbfcBXeZSAK/UE/1RV1O0HVKc9FlcVa44pjn3lhX/nQRV5QszJB0Ur5ZV1iqTsQFpVsOv5UcnILL4r2svXQZPXSew9OuGFYHphZ/ESm2ijJor8ajltTzqY4mfbqYsdg/idVH2wSCsvEqmT5sEobCE2D0bFehYTCi3D3sL9ww4BfsK729ll35XYvkxXc9P7MNmtvenNPj3JwKGzUYi6qL8664OQrwzQ1Lf55VrAWQ4zxrOQ+0FyvUm0lK9r7A2jP2AE0G2OCNZ8dhIPSccy3HoHNQ9LVUUX16pbAFKnLnpfnha8E3Hl5T6Q0SUUVRZ6ICVe8Uk0W8wO2mI1Myu0TRVVW5pmcQOp9QRSiP8hmhbdAM58Fxg54Uv6n6irCgs7szWy2qk7KGvEX4uq08OKOZmoA9aqnp3LBxL8coqrCqkVxaLXY6EGVZyjrw4mIGm5HG5m/XI1144dVV+QhaQoYkgVPKrwrMLbgN8wqwr5DUm1OZyx53jOGxruU+0Iy4FXRqUA4cSxhw1hnOJ41iPUgvq/kWZeu4DVHTh/G+HmtFxKB+mavEeyqZdOLGszXrsins8ZNtZnQTzwvIH2QI9I2+U9WnTUzX7YUxilVrTVcLft98sEclB6lAimBfG56tZqntH1CukH4p4zy27jyoatGoRNW6mGUEQumUFC9Oieby3hBuUYkwFhej+Sat7Y0kj2JBBIJJBJIJJBIIJFAIoETSCAhLBIVSSSQSCCRwKMvAQAIYxXICyVggEkGyf8AK4R5IrwB1sG8PANOAApiGQgggOU+L94ALwCakB2AGyZgCmzFmQTmHy2ptVqYA9pi8YqsdjRlAViKtSxWjIA3gAMQPoTQQkYQBsjGhGI6GyaHhjDBXhVSwoQUMda8jA9ALe3jWCokBoQTABeVsaJtcCqxrB8j4/do6c0p3fflI/+s9LTO4Hht23P2Vi57ksgKO+uUJ0fTh/fvyO25c1f2/gmRGXs8u2H07JSuv8bBDDSA6A3t+1H6gbAh3baN9w2bKlXbqU45GVlrRzXtP66k3Jd16SpEj1FM/DgIlBJtV3Qw64sBqwCsmDvGw4LPWMma1tqAk6wrALPtBUCR9WaH6nrJjLk+RA4W1Vit4+IVW3fjNQJxoUTAJsfEMkFDN1WxiGbu4E3BvIitummbQEvmRloUCHPoQl3sYsFvu4TT06fVqLw2CoAnsXAQLVoVu6LzSsrXLZgw/a5HFrgjx4FAUOMZ0zlolR1elvHnXnj1kb8tbZiwr2zY6cEg1TVqNaqbq6n+u7N2o6erMPYjTqPSn1c6E0gKT0kP4qU9ToUTo+ExQVHqzlmFnpz14MXbrPmB1bnMq/nMA/MD3R/Ll2t7u9Op77qFYqjLBDj0qP53DdPf6HIQqcZrjctDHpB83eQBAfBd1p9V2nLqG9BrKiTzBap4E/6G6qUk1VaiH+sp5QfjnBV35C6UTi1HR0K3MgUnl9W2p2uYeT7OSN60IM7dogqozfoPAcbzlGclwPVPqz5L1eSMam81OkgSej6ZEzyHmR8n4wXnuK5jOa5dUeL7SMhzXQ9i3GT65SwTaNQKIiy6SE8ii/mqtqW1zuc1hDKKd9LptNPT8KNCPQwGM2n3e9V6VBZx0fGZ1Zy7PFMIVfUO1V/vJP4jqRHrW92XW88o/UCkxaLixy3h1yRZJ68F84XZF0IdMneWRvd/6C9GEW9TZe4BtCPjjuB307sCWaMvJJknzBbP304F8ge6C68tnt8n+0w2ZAXjiJcDYfTQGYiP57TdyOS8YvPHVSFd0AO8KFj7lskKc57kWfqr770U75IfBK4DAbKCJFrszb+gnvYIC2Vlq2um22B+fLrZLrxyMDwZU2Wd56T1yIN4rRCJhWPVkMiLIceOBlOe2+VK7zVR0RXyl1TVATzrsmohBLGv5NtTypNi4W2hfZsWSsHhRiOsjwwqVUpCWLSpRvJvIoFEAokEEgkkEkgkcK5KICEsztWRSdqVSCCRwONJAsbi2YQMoe/G6lnpMGURvAQSGpDR5LQAgDEhpPgOIMAxvIxDVvAiHod6eQyC3YD/ACeAKMSLBngCwAAkoc+A/wAEgBKAX4CeY6qQGQYU6QhwniHFo30AZcbLgu+ghrT5IlW8YgAvAL8AcwgFxJihA7SPduMhY8AbpyXHxYomJjkuztCINS8D2FYKbs/Iq2KoHHb3CfapiJyoeArQIWB496A3tTDnj0z0enOAg4xT/XS9K9rCQgGCor8r0K+ml8VCf9TYty2soA/oiHfUydr73C48Jwrsm3dTzxTqKdQ+gqSID4txbKWnEJhVVzX5L8xcgGwhbjr3jcmxFkkCVzJ/CAGFN4ApAO2EhPp7VdaZo+19b3pZcE2uD+hNLvCfLDk562B6gzXj9coafosatPonqPryRR1/m1qOXGcV2mf+hYu3NbY2pu033Rivb8z17ZrpWMPj/XFBnMeipYHmq6zDrVA0ZRzmpmFtlCfG86NJ628U7uYGiWan4vKTK4R1As+NkwGfO9zl1DZhCf/xTz+jsNjX9YNid+6dIhZ+rf0KPYXFXV3VQ9sG5hdqdugOyeb+ScrrvlMRga4IbQ9r65iISvliXgQ2S2axZ4XdDAVVyWet8U1D1vRIn3V809CMyIqOQLzC2fgHdm0u5crVrx3ZNjL9gi/cwsWU0leEkB2TRYC1nRIH/6y2/5jqV1X/RJU17ExYbRuLfNZl1k9yAgDAXoqMCHFGGCNfejMULFo55R4v2isTboi0+MOmPGnTXzV10ORDgfwg8TK5HgDRn6PK82O9AqD9OVXmw9dVISx45p4S+S+reNyb0pHUTOGhAsXtKRPmR+QD01VqoIwkga05GGZ05ACukLpFSuF/Ngh0xhNwWqM8Is+MsgJ+GW+oVe1ukhZ4KHxIlefeS1RbCaf4nMMiLW7LXRQ9s/QDe0DeOa3FwS9RxdbMCOUfEY6pJYxuw3qZ2oqnxFtUb1KFtKAtzHUTUg5Szowjz1rGDtCeedap8FsGrwNoETwajIfVimMh+zT/Wws6YgafdYGcIztUySHRqeDpQaGtxsuB7zxzKSvGU2tDTJx9854Di7NDvffPDfZ8rpzPIsvlUu7KZiu5pZBkhKxTmKj2+9I38lMwjyBuISlYb+M1p/2e7SfvOThj9fdkHRFaofRHa7a86BynouQ2JLyi7Ru0vme1vo+r9TXdfUCN7m6Ekfgxx63X6zwGyrl8Sg5aoUgwW6Gi5IeRlEQCiQQSCSQSSCSQSCCRwHkigYSwOE8GKmlmIoFEAo9pCZiQUFit8uLP2gzMZjwkeLk1iSSNZaDxygCkB6w3SSY5FmDSWFPLKLUTnHdeyzMGbFXxnABeAeTAShMSgBdyyB2+IwNAZSy4ORYLTiNLQCcKwjmTL/FG2LSPdgAaGY8ZABwQDkMkQWAAoJHslfElXjbjCngMUAe4Qb/QA87jOgboOJNtbooi+WhKID3T2HBZI0pfrzwVg9Uwv+Aqu2kjSik3RBjcYz/5yGBqcq+IjD2Xdt150km215IupAU6obwZgFBUPIBWFCl83wE3/4RMFM79l/oEOhDc6/V0HXKyAkHtTdkouDpjhVdsVFx/W4hWl5YRR6okIqMYRnbdtUJAMnSecyHEmDNzWhsOy4K3nvK8TCbjpP78o3f6/oOW7+SOVO2Nn77LTs3JQrrJpz7koAVp8MuqAL9YD69KwNzMCVEvfyXzfYXo+Zd9mc23CEz+9fsy27eSb6BTSUV+/crq2Ef2p0e/JxB+cFdtvPHU8v0DAqnRfebA9ao/qgoAChCKNfXq4lsN/3YZ4ZssNUCVhLepWc+Ay9F/JEH4puq7VZljhwRQTp9p0sKAnro+c5V1gX7krE9/O13NpoeVk2PPt6+/8l8Fhr5GYZuqQq0B6SEanlrq9rZ7YfGzio8PhbAziskd3FNkV+2m8LYSQCocPiamICzwPhBqqTBQkBXjW4aqi71d0+ObhzoC8gJX/04Jub8r0uIrut+kAGG/JeQO4DFkKkmXf1H1ZR2kzJoKoYCXDPoEubpugus1QvqYS9NB1kqs4xkj1u0LVX+q9d6QM0qqbXWFVWtn/fjk3dmda6VXx7L/2aoQDKyvyB75PkP151XxcDtReY8OIAwUzxh0nYqun+zaG3sAiGzolrdEKKYJlwpbDhd4zSmrelQXeVHQ/COnBc/+ujgMDazdsAO7EQVhTltthfQp25Zb1SArR42j/MthPP/bG9/0JmEzExYjhw+rMi6/26mjY+nRKQWPO/iM0r1Bf1B82nJOi+YTjLBQLn4LalnIirQUIqpHd8YjBdcVQsYBxrOuHPjmP15a3HPxtpSQdeMhuEPbIQc4dinxyOpC3g3yyhii/kTEF61jHPnNgzcW92B8IS9Xeaa13I7fTXhu8czlGugsv7GC9vw1mreMG30Yffq3f3DB+KbBVC2Tzn/tedfUa5mUIT7iS//gyl1W72LJ6lsoWbmy1t6mN6R2fbR5D+7DXEKC3M8YonQURttGu1Lz47CVMJT6WBDfMG3bTr88LVAMRYaKNmgpgMFEz7h9GHvgKNO2BDooXQvyGc/P92UGXFtJmdJK5Z6URAKJBBIJJBJIJJBIIJHAeSKBhLA4TwYqaWYigUQC578E1iAO4jQK6p0J3WTCVxgvARO2ghflQVVjDQ2gg+WoITtMSCEEZaylH4svpwbsp+/IACACEADgH0tirEkhCgA4IS2QLeADABuyRE6AVxA8AHOG+DkTCmbID9qGFTvtAswxIXT4H8tfABbailcF5q0GzARcpP30CTCG/wFU96uiD7HVuSrje6aJljPR/8fENUpBz+CsP/KkifqWC2WsOpp3SxnlX0h1uUVHpMWRjFO5fSQ1vs+PUrXT9axYQ1DojdGPVSGOGpbzUpEUB6/z5w8/qKggD7hdfUrCvVluH69yotQreoRTRYolUxS43afvg2G92Bc1JqUoXMuAyugQen+c+OdYdqdSjpIdRNvL1YYvK9y61qNSUN5SdRYvHncGvzuuhBidmov+/pzqfQJKx9BzvAdaD9T21PuigBwEw/Km+CGRJvWazVRcXXqCsjUcLKZ31I//2eWVsdeLZT0y6Bc3iyBirjCXsPjHuhtQEvDThJNqv1hd+S3+WPWJgjVfygoZh7R5yJ7ZeAxwHa4JoM26eqeASiObjh0WobFuaRIUrCcmDxHrDQCp8a7i3gDlYyIiNnYXK0/eeHy2W4QFJvYxWWGK8nWMjEzO7958dHq/5zPdNYSx0T0uMyItbHtcJMW8jO1ZyzY00t6XJjYOPiBPiQuObRm+QmFqsrounlydyp2yCC+EjvV13Ze1ppN3CesnSZBNWDuA/vYCCYwHDl40t4qQ+LI+SXR9Kt4qPPdgsCAFCMvEukz+FJI0v7lT4wkNtbEx/8n+oHTjuDc0MO314vHTXmj/i1QhVToTW2sIp7mZUFiAzJBjeApNS78Nyb3+mQ/tjUP6CECe9/2g23LdORnLD2sKHNM8ywheVs4BkRQKDyWT+W7RUdOu5ZSFRXuac4rz5ZSVw+KgjplWsuUZZe6eKpZqjVrNr//ea5+ynozRX9qKHKHtaP/72xut0FkbDqRHNyg82z6RFtag8oMQaqs1rwXnuPL/s0UPyENpydtiQcThEq0ASYAHwY0KmTTWXajcqnmbSTV8W2QY8oc0+i3VTl46nP8+Vbwq+E3DHO9IVuBd0SxGVyBMoVIoPEN/r71vbf8zz8mnQ+4KzsUzJL6fISs0d5m3VO4BcXaJ6otdP9ixYXK+S94Vz9swMWsd3t4avU4XGh2wbn/yxdFVd+2ztxyZtkRsQ4R+UHVMlYnLsxujA0PqnspvskhJsuVUYSMXIuotyHGiV55GW4LQ3hCFoaMGZ7WGj4r8CuJlgqh70inxXmHKtXuUB6WhxN3lRsMvKe2NPzlTOtlwWycQabI7kUAigUQCiQQSCSQSSCRw9iWQEBZnX8bJHRIJJBJIJHAiCcTARvy6uQQe8bLPdxNvGGDevOjGlpiqhrAA6AJU4jxDXizFg3nsFvpnEkjSf8AF40UBSMgLPiQBoA2AJGAYL+qAh/tUAUiMtfmZlJOxpDbACySTsexljAC/aAdRwgHRGEsAJaxgsRgnNBTtNrkBAE44hnTCXBsQjbGPLUObVR9JOZMSkBVzdrqxcaEQ9B3ZmjmQC6Ljvfsql8RjkbIb38o55X1Zpzp5cf77Z1J36AJjDGgOuAVRhUfOctHOq4Ri9n4mvRG9Si3a3qVaJK4ROPUKchgUtFzQIOWxsPzQvnfUqn1LCblHc1HINQFf8bJgTVHu7hg0nRT+nReg2qsY6WURFVnNKpBxme4qVs3c0+ad/js+Ytn+IZkOA8K1F5LoEpoJ0PEbIiiKzZA0Zm5eJK+K5wgYxRp60rdcwgitKnl5hWxvTFm9Ii2yYWOoLyh9SuQGxBzeG1c2T/iKPjl/PfB5UhJ8h92vlAGXWB8I9li3KBzU/14nWBFx+U0BeP+MKl5OzFnmaSvVEQnUbAcbDdFsYulzHkQOoCgEEUD8U1RZdyBPISMJYzOvJL17u4qVLdsPTTxBXhDzC/3dsZuNKTPDfZ68L575Q1+6LTMwuzjjBuGQyArCE+0QYTGt4SZATq6eSX11Zqj33oM7Nw1OD/dtk9fG0xRXf5sIDZM3p13erIeEoaJ9rCdxbpD2g5r/038s5AGdkU8nK3najVcE3hC0b0rEhfHyMyH3+J9ivM/Ybohn5EE4H/QIcopjIRnI09SxCLD9PXnj1BSB586KIwejpeMBsGmHKSZpB2SUKatIwLYboMdUxhGUHC+FOBmz6ukAvUY/hC1HXZETLQhc3q/cAgPiFOVsQdqKcKc8JjwREmXXc44qgXLRD8OtGDco+za5CaK6QOtcLlXxPLeQSXvVTSOr85F0EBRyYb6zJCBvAHtIulXEk3Ja7L4zt/vW7fXJHRv9+ZGBoFCVqX4WbxZTHPmxYFYRQW/RKBO8MLReLF07qtBIdjWXHhicXWwErnvk2JahJ4kU+4POIxi3CZIBj0fIFLy9Gm+a6qyHCgXF/EKWrHvML57xbMODZk09ad4bDx28cBhTrnFAtWJItSbJyDPWzD/uQegwOv891dem6v4WL+VbV9213xqcKcQ5YSr5pVBQlOkN/dVCb/5IqTs7J9LmQXkvMbfQHZ7tsYGJyM5TISqWr8250p1peehAfBBCrFu9kCuHtaCcKGRonyOvRaMRucrFPa5QUN3SnYb0aFrHiu9yj5Yr9clCqT4vT57GEy4Ysu84vGhds633dNvT2rbkeyKBRAKJBBIJJBJIJJBI4KxKICEszqp4k4snEkgkkEjgpCVgABwTygmwqxnMJAYegAgATSmAjybRqQkfxfkmVIQBiB6LL6UmXAOIAWAUMphDEWoAACAASURBVAGIAvgyKAKEAPsgCAAoALM4DiACAAEwgWNim0Q8XM5gjg8jcxNjm0+shrkvoCVAImMHmAE5ASgNIAaQaAgnLDIZQwBO2k07AVVMSCgAHkBok/j1sTjO6t4jXxSWyb698JHS3vLlA/Uofa2Ii7wSa4/Lm+IrxaD3WbYVzoxVLxrflD7sn2HvCtNZdBn9IP454JyZ8+wnTNi2CSczodhAvSIqNgmBex6DTyJrklQEQkJ9WaB7dji2z81PPiEojfVbjQXtIlk2gB1EpwxyLXEU4ZSsd+VXYS+CRaq6Ark0GayaAopUgiAdpiL3mGbI/TqH0DgkW24vb9UGiAX0+FMiLbi+mZdY4D9LbQPAJ5zTqrKtPmUNBoU4J8GW+rTVF5aFrsY8ENd4XcsJa4WUab3mq9TDCV1gQHDmXlmCf1crA8TPa1SxBl+vkKcDwPwfVFkvmJ8maj7zzcSdNyC0WXNYp5nHWHqzD3KGyn0ZQ44D9GfderoqhAt9e7q8LDaNHpvp37l/PDqwa1NNpMVDKKgOkIdE5r7LLnjmjgPjhdHx2dtkuT6mzaxdjgbpsADivd955hWHZc1+qXJilBXeqaKQNc89QT/JOUHuDtp6otwrqBa6eKvqr6oy1gYgBrpmnaJ/hOn6r6qQxugKMgGIxluI5xOyYw2jf6xjyIK1C+IVkhY9wWPmaSdoO7v/jnaLtNgjPdlHsnnVd0nHmCu04RXrXEPTpsmZmPBm/L+06W7ILv1zQMbpkGSAzlRCvp0oTNF6zaav9J1rzWcybt5vhFfk0+luRe/pq1UF1ttWScDysBJsu5p+pDwnDJCSKNsN17WLOVteXZ53vDefKuXSLiGhTna9ZyLxnEBnCLsE+dLJU8Z6MLP1KQfTG+95fuGO73aFlQsVKuoSPC3wZmE+xqGORkSijChjguj1cK9aPy9z/sDVw8v7OQH2eP0UNh2buXls5+isyIpOa4WRE21hbvDMQ4/M7xWz3xBbfPL8NGQC3knoCIQFYb3WIy+5FuQTfaZCzi2IqIiJp2bYJ3STyhhxTUKfMfb8NsBIIO4Dfc9V6lb/XMGa7+9eQVawX2RNbt/uLXek6/7ddjTzYL5UvVsEI/17OEQFl2acY+JU6/GiyC478OUX5ToTahIyy9d9v6bfLhDMm3S01MhRmD+rK/ADeWQ4NV2glsumRWzY6Z6uTHqoL2/yjXD9pCQSSCSQSCCRQCKBRAKJBM5pCSSExTk9PEnjEgkkEng8SKAZKgqsgpdQXp4NIGFepo2lviElEIuxsAeU4KXWWHsv4ZePzQKAQd+MlwFgB6DXUmz4pQJAA1AGgAVIAdEDYAFZgBwBPbBWRF7GEvxMWsq3yt4AfhASjO12VUA9QlTsUMU7BDIDEKkZ9yVuJ1bZY6qAhVh5AgbTbvQBwgMwBDKGaxK7ms/HYq4SdesRL+5/zr68q8stdKXt2kTB6k+Xgy55WXi7gsgt1sPMEeW0KL33mb/zcEDM9TrFWAIQAwITIqe1ECLs/1GdVopldP4SKdgyaEf4e0rZdkRYeDenrOh2HTclxA/dMrHT8d5Bj9DNhTje+VISX1PjayjkTNw/ERB8jqn+q+orm+e2t/+/aAM6jMcFYVfMHAC4B0TuWK6p7J3f1Jjth7DoDipxQuUmWbHWKWtt/3ftgJCBZNini2SUi7muFZK1gfnD/Aco/6ETXPgF2k+lALzjjQUBADAPyMp6gbyRFdcE/MO7i7UHDynmKxWCg7EiFA6EE94HgLPMf6y9IXA2kTA3U2vMjR6fLYl0KIqwALhfUe65apclb4s7n3zLfe/tWSwfzJdrQwr7Fe7fvfnYvZfvyOqcdMNzt4Sue4mwd0iT9sLYM95KPx6D/d9RZXxOJZwZ/YTkIEQT93hts7+sS62eHL+u/5ET93uh6jtV8ZSh/8iEgj6h14SrYmwgbwjndzJkxcd1HB4wX1cdV/ii8s9e88VAOvo1/c+6iYcH90O+kNOblwgKe0YkhDxUlskJtqlKDLbGObK/JVRac06J3hWlSZ/fteyAZ0fp4ZAVhG162wduRXZxXiIxDX2LhajkeQrnVW2kBS4TvU18qLVLHERG4X9qjutOyPNJcZnsXkV3m5PrxTGRHNOa0nNyySjksqnGi6/d0vF5ZUInteSyQN4cSxuQDc9L9A+PmVVF4dquuLHn2p5Lq4e+qZwWTxBpEXvIyONJ4aIWY1JUjiFWaoNvpYd9K7zPtma7+qxaI2UVlG5DBFuPwpH9sJLJd7q82QZhxrz6qiqehRC/8T55Uhgy0HhUsJmx5NkHeQ+JQE4Vxnq9gg7c1Owzz0r6Xa5/2AqboZ9oIHrHdSDXMACBOIOwIIxVq1dOfB8SapOjQqQhn6E8LGjjcjm6beS/Kgn39KZj09+5cM+R47v+YLqdhDlBk1fvlv5E0h/zO6UgHTkoosIOoqBHOrJR/xOsT1GfrKqI5wVHypLyHKU+CR3lt6jirZNyvQl55uBNN1UuN2o9+SBKvCtOeSiSExIJJBJIJJBIIJFAIoFHSQIJYfEoCT65bSKBRAKJBDpIACDJgBExCM27cvMToAfgge0m70JrCCgSsT5WiQojKvpnrC4BGgjrBICGBSbgP/t4rgGkcSzABJ+QAgCHACQmHBPfsfxdlTD4DGgm7TBAEfE7sN403hKAIYCbxgqdPtA2zjEhewBSaB99Yhv7AFQAHwGc6RNEDN+NR06cybW5b0UXHoNJ18/AEK15iZwwoZystsdsO5wq+H3XaloN9ngLpUqQ/1o56r7bD1LrJhd+mI1DbyCjiIUOuNhuMQ9hcaA57r/Rfi9ICynL+5XD4v3dkV/yFD9IoV2MxbIh+zitNaRYCDjGRgN2toCebEcHAfD/j+qqezbbADnxUlXAfeYYHg2rAHjTXsm3WLdTH1VuEMLPCHz2f1HtZI6cbIGMYH4gC9oGCTknC+pAIYkqzmuWrJMFUGJdDmAp6/k4pj8A+xtO4iYQEZ9rOY7zkANhdZiveFC8v7mfOU7FCwRSFMIJEJ41aoeqCaDDHAZ8BVBl3s4r5v34hom5TQt9XQ1Zp+9ReCi8aFYUbbvhSy+6bkxhpEjCPaVVfloeFS8QLIm3A/0jqfFa1uaMPevE7zeP5TtlFeEm2a1X6pIrpAdEDbIgP0SnAilj8otASoypIkf6C6kEkQyRsSJ58bp3Xrrne1QZv5tUkWcrSc93rs1a/rdaLn9EKq/xsRXmTLblVghJvHmJlIi+rO9Y0RNG6kP6/5aw0TdjO/WcFaXyQWXjlPiCehSm/V971tvPBCnJfGYMIMw2CExW2mNXFvKhtrmbskpM0XDCvChDeVxYzNXFVMqtKWdyLZ9NHZJV/YT8aWZTIrTkgFPt782dMDRVS86HVrEuak6zbv2TKvlBDDG3QvTKNXPBXbldsS4puXl92F9MQygWnFzcidHGrFVyslZDTMvRK4esw/kRy1PGBPbPd/GY7Vw0x+d6F8tvrGZSffK+mJU3RuOJd+wJnu7d54iooJhnJr9tmF+sHax/tBPyiWc5v33WIyvQD3T0Y9LuRlS2xv1bpDt1qyxvK85nPjIezEH0EB1EVyGnMBIwBDFzm/WM45cap0crpIVIw1BzltwurAMrigibX1zo79r7wKUX7H33y53F9pw+7cef5P+sY7HXnR7vRa3k09LtPeoEP/aUe8hyREiMiNCaVfMc5TcRYRrNp5SbRoqymE45ReWvwMDDGujNBYUSThdJSSSQSCCRQCKBRAKJBBIJnB8SSAiL82OcklYmEkgk8PiRgCEteDmPQxY1X1gNQMMLtzkmJjceh4A0QAPoCNUk0gaIAyQETMPLApALmRnwwwBHAIucjwU0Vs9ng7Aw48P9+Q64iuU1QDRWolh9UmgD7aSNjDfACW0CWKKN9AcQBQtQ9tNXQq0AwHJt+m8sqI0Xx5kA2ZrNe1x+yJvCHVn0+wfTTs3Lu0UlynXGq2HuYwoJBVAKwXS2ZQzAdJ8q9+tUfmedkdknr4rcQTc3tCF0Z360PokuxWbmqoCBtH2ZGDVExQlGGh1DdwXwxqAxlshreU78wkloDf16177Mpi+JuHA2N6aH1DjCSr1EFbCQ+QKAuFYeBizqAeB3qGIRDbmDVxVEgGUS6fJdseMhLbDu/4rq3aqAn3hivFF1Rd6IE7Sb+7UXwE7aS6gn2ox8sQjvBOYDEpuQTwZ03SPU8R4Fcvqywsg80FWqQPS8v1M7atn0T9FfWXajF1Tu+eJmXa/p/6mdeHSxJtI+ZEGYo9MBLlmDOB9CBk8KCCoK+moICORrCoQFtRUcNyT8em02+0ziaLx7WBeNbhgy3xKJotGM++L/xcjLadt8WO/dH/ldWQXKUU6WerfllRq27TM+ANDI/jZVgG3CNC046flCWB2u+AuXLTbmro5srxSGlVHrbR94uX2S8+NEfaHPyJ91WwmTldQ+sg/6oiUUUmkul3EXRLMPiijdIVZnWJ2Z8Vz3oPJV3C+CYyKbSRVFXMzKI8PM3RPdr+N+jXldpAXPGDxteF6+er0LiVBMH0sNWdStyjGjXBfWRn/OKoqcgLRYLisCmXW+4mX3jk1o1blky5GpKO37Ts9CaXSwvzgkWkLUgp5hAt5F2sCDZCQLQrhB7qGvrSG+IAzXKu8UFfGAVrnhqGrtCw9Zi+ED1qhICwg01i4IBnSRuQOBBT0HiXG9KjrR6rVCzqt2Qq0uwvA3FRZq47ZDk7nxzcPe/EA3c3BFERnDPcilMglBdJrzbPmaTS8LQ1oU5BGXdhyRMVEkz0pL3+VLZkdOIIXSvtB1HDlbOXURXH7Osyddxz2cSdskeolDk/34DbvOpDfpeuqT7EskkEggkUAigUQCiQQSCTxsCRiru4d9oeQCiQQSCSQSSCTw8CSwZCC/orSu0SZUVOtB8ffHC2HRlI/xosD6EmAAcAHAAYtIAC68FwB2APn5nxA1WHsDTuK1AAgK8EV8a6xyIRKUhPjhe6e0jZ8BiQE+AMqMZSwkA/ekzYSMIVwKIB+AGta/ALAYE3AOVqAASyQDpl/EygceAvgCtAUEA+Q04XxMIvEVivR40Q/J4WEV5a9gjqEfgOU9iuF+XKRFvRGlLxOJgQU/YVXI0RCPZfUVp4J3n7hpur85iHag129RJXfAyRZ0BTKDsDkx4aE2xrqg0CLxWvJwAFgBcKCUdBq9fb8q+hmLQrUFwVy3uX+mvcDMyHJBIaGcFxVudZVwGyIRgo5wMRBzWMAzDwAcd6ii+9zjs6qArt9QxUuJeQIRge5TVup+i9dAM2491+Y+AJjIGbAdrwZIhlXeDc1rno0PE67qr3Xxojwsgq/+0JOOzwz3Xl9Pp9h2JgrXgcxhzWG9Y93D8vt0yIolcmCJ+ALoZc1CR1+vSvinM2EABRGBJwJz7e2q6DP6RugoQGdkBjHbsf14iDT13PP67rdTA3fZTnbCtVMsk/HzgTbSfkO8xESHKjoQFe/+Hf434dJiz0YTGi3u+WkW2tQEnhkH+sM9u2QFH3qunc9kvC7Xtruqfni1LPkHtF7v7+3Kzgh/PiZC72h3d1ZpC+zirq2DJm9Vx/4r1M8JW6g5TL+YR8bLD+LxOao8h854uWzyoNVTKlt9R4rW4LEFq7tYudezwv3Oxuh2d2eUF9yuzmnuBta9mo2X2Wl5CqXiuXiyiytrz+2S6IfCCeveaMJKhUesnEiLLj0Vf0z7WB8+popXBddl7MlVsxYZ2kkGP4EuqB6XV5O37wlbD95z5a7U8U2DeA5hgNBe/kIbPqiK99NJzzfpyXryN/OOuTcgooLfPhv0qehP9lZ5XfS4rrUgwqIo4qKRTrtF6cxMEFrHpWPzyntSGBnoqiWExRlX8eSCiQQSCSQSSCSQSCCRwFmUwJl4wTiLzUsunUggkUAigcePBDoAy63AxNm26j5fBM2LO3IBZDLhkQA3DcABKIQFNygVIAVW0IBcbMPSGKIAcBTw52yS9mbsaCdgB4Ar1td8MpYmVNQBfafNbAdM2akKsRLHUFfdoQq4xP8AqoAtWBtDxADSmnjffFJ5rhvPDn1NyilKgLFCX7oUYWNRnhXIkvFgG+PxSMxD2sA9Fd4mJqQIZ3Sigp69TxVPAsIyoRuRIUHepu9ngGBBBsw59O9XVH9SFbD6ZMgKCEQsuyHc8CwCgJ4dTw2W+56ryD03xuGWuDaANaAcYZ4gJMZUP6DK3ABUNawOeg4Az/a4rycIaYS3BXItiLiA0IEwgXBhPLkmoCahovBkeCQKxAlyY52Y6SlUGoMzi/smNw6wTjGOEAEPpwDyQ+pgpf51I6vTJStaGkJ7WTtZSyFO/6/qF1Xx9jhRYvMT9Yf5hfcLeTZYy1gT8egB+GUf5URkS0wU+wuXhKoBRIFAeraxflKMp118nVZ5vO0DseMS+oDM2O+SQ+DhkHymw00ixcwf2tCjnBa1MLTn/CBq5POpybQSJldqjYvTKVfh6KyJej0g+XapS3lmfFUREg/bOr4ZpqgsmaD/gN54yiAbcogwl89YuaF4t3WVc8Aq9mWtUL4vuS1Kzz0XXGY70WUiKl6ip9Rd+mQeHNWoPFE+Dadyf1/nf0mj1B/OWncG9+g6ZSsvomKzrnWNtrM+8Kw0Bg2s4089hc59UseyHn1eFR2MQzIGrnv/nou2lkRWELKKZzA5NdrLm7SB53rszSRZN05m3knP1mse+SzMb4lQpISiatkV9dMPg6iqVOhbtCUKnbAkcmJeujWmkGIN13MWS+V6MZ3ygj0HZ040d05BPMmhiQQSCSQSSCSQSCCRQCKBsy+BhLA4+zJO7pBIIJFAIoFEAmdOAoBJgBxYzFIJAwO4C8AFgAnAy3fASIiA/5+98wCToui6MJizvzkLKJJzEhRMKCqCYMIsophFVAQDGDBgVowYAEEkCCqiJEWRJErOGSSJCogRUQThv+8wxdfb9MSd2Z3ZPc1T7Ex3dXXVqerqnnPq3ssKS/JDfiISIGyQIEYhAGL6BM9F1R1BANHEdSAjqQOrQqkTSypx8QT5d60lVi3zXCaxQp5V4LQR1xMQuJAvELSONHdCB20EF4gnsIDAdS7EclH9QnkqYwcsWYVfOYwnfTE33G95RfrQz8ss9bDE2L0/Qm9ApkE+Mra+suRElXQIK7SdsYsVBPcZIgNjm2vizilIuEAcGGCJsYrQwfiEzIPsDq1sJ16GLUne0nrtQNoA9hDiiC60G4HDBbPmfoH0dSkH+RwBnx12m3ARIt1NuOAazAP0OUQ51gjcS7SRe+iG8MnUE9Kbv9y3qdggirn3saj6xfzjryw7d9nGORVLgAtCFfPaPVEuhDsjZ+FCNqyzsEyYacmJnbQNzMB8S4TYBsm0BfzAZ5klcKNve1nCHRir2BGWEolHQh1Yrc5YZsU6cx3YICTRprgEqbAo4CwRQ64TWbVuvHnIpY6HEI52D3OMBHbMwwTODgkfyQDFOe5cyrGvzp1VyKWfuYda9d+W/3bdYFEWLBbBr+baZ+ctO29dY25/1v276b/dTbAIPaPSsDKee4jnJaQ6xDzYE1idMY+wntRGgG4L2F3kcHMdddQmi3VOI7f8U6ToMebzKRS2OweMzK9s8Vt3bLF7f4uFa/qtyA9bbFQX3b3I6i3Li/yy9ZciZ9j+f614RAriWmGZxfOSLVrcC287cUtXzBIxKpiz+MyGleQES79Z0O2Ny4uHisWVIzZH3K/MfbW8BYXPxeSFOQxLzqTHj6dcxo97l/jHxsbvJnZhYWHzZtEfthbZsuvm//ha5BeztFhrY2vTzluLbLK4J5t+XPtnSoQ3Xxv1VQgIASEgBISAEBACaUVAgkVa4VXhQkAICAEhkEIEXGBOCCxIOAg7CCpWb0MusGIUIgGCE5IBwgvChx/6rOqGTGM/5DNkqxMrnNVGrqoawfUSsbC5PmQsxC7XRbRwcTaoP6IExAbtcSIKJBLfWWXMMfKwj3MheM6zBIkCMQO55lam0xYIEq7lyLdctasQncw7Eav7GTcuIDvEHqTU3869Uh7hESJZw33e1f5CxJ3vuzYk732WGFvEOoGAhMh2rmPSUVXqBenKNVnBDzbgda8lYhrA5jE2P7KE+yYshhABEDkgovnrRDc/icd37kkS9zjj3fueGmQ5lDQRGLa42GjCBfcMMQ1oi4sp4+YaSFXGAnOLIzCj4UodsXIpbgnS3i9wIOCwerunJfzdc38j5Kw+ZM1vm01U2GQCDjhxHOGkQ4SLUVcnWNDvr1tC+CRYOPgyDiD76ZukMYrSUDe3MA6Ys5jHIHmJmREKMG0J8YkV6FjAIaqRmMuoO4IEghHjhbHNHA5u71tCBEGwceMhkfq7euXGGoH7zrmPcq79EqlDJNjcvQMu9AtiHNf6Z9PmLcaFbwHHn+15sWH1uvXEed5sosXWdKyMD6/4/8/GGvcYzxHERlyrYc2CyzfqSr/FbZVQbcOiItX+Xmxs+b4hkWIP01pszb8NglRAZ0z9yiK/W9q/qN1RJlgct/Vvs6DcUmSW/T3LUEQ0S8RCw99HiBQIhPQHz1fGH/ch9zMYbe7S6gJvQ5gTEAc5xuYXLLBAY07BkmwUfey/YKLfw8IXIhz1cJaAu5i1BYG2fyq6swUX2dZxm/75d/MGuytDMU9yI7YlWkflFwJCQAgIASEgBIRAKhGQYJFKNFWWEBACQkAIpBsBR0Txox2SDKKCH+aQfrhMwi0JRBjCBG4bIL9wDeV8mJMPUobjkIUQo87/fbrq7shnykeoQEyAVGQ/pObpliA22U/92HDRAYnEPuoJcQ7Zi3so/G8TjBTCE1KE9tNOiGpIC2fF4cUqXW0rSOU6AQv8XB9B4rkg53ndVkfYYs3Q0VJnS/TpBeExAElN/0N84vYn3WKFt/3Ug9XZuB6CgIXYhYjHdQp1WWYJ4Qxij3bwF3Ib4i6QwQxw6eQI3rzAnWtBPk6z5OYF2gGZXj9cAY4hlDq3bRDMuJzjL0IEK6rfssR8AjFPe9lHfsQFgv0SS4L7FBzoOycuQIgW6dwqdCXGHscINk2fki4K58X1EgJQD0uMV6J04M4K6xAsxzgXiyDmmXQKV6GKhjfmJvp/qSXGAnMy9aD9d1hihTuiCvM1czT14h5DBMICBLc7YOjmMLeS3HuNeD+nSqQFW+caqqiLQxFvJSLkc0Qzf13/gAn4uY14Axs3/7c9LtF2S5EYLoOSqlpYuCAYN+1lTFKv8eG+Gm1/se5j/HNf06f07XqL77PY7CXK7rFl05xdLcL5Xlv+OWDPrebDqsjO/xy6+TfyFt3VdHqsKnJstIYWx7OFnXNtsdlvy7IQSvuHqHmr4VZqsk2+rOi7BOMMET/axpxVLZwBYQLXTn0tcS6/ixmLCErgEcI/nLxlsh8xgloEWZZR+9MsfcBJuCWLxy1UPLA44YK8Ni6dxc7W//4zlWjbfYg1BZZB6XR5GU9VlUcICAEhIASEgBAQArlCQIJFruDTyUJACAgBIZCHCDiRAoIWgh/RAdLUEYOQD1AZ3h/qJ9l3ftSvtAS5wCpfyAZWAfMDn+fgTphBpCLwdhAWYcsLLuHcNLn6uXgTkJOQjJCjzhUJxBDECXVn9TGrpyFU2QcBCO0DQUgCBzBhcwQK11A8i6AOibyPcYHYBSlNf4ApZHFEkj2x4pPKzZiH4J1tCWKMvqY+kJyMaeoMQU4eR67tcKEUxK8IqrwTFCDnGG9YJ7iVxNSPscrY5TPWA6lZap0UjJFPCruI2mqWFmzUlzHgxD5EF1ZSIzjwGUEQQhaxEMISSxLmHMZM8fBnxg0CDfcocxKWDmwc94owlAd2fvddLg/CKvMbc8AoS6eFy2McMD7BF4GTceAIcNxBRQ3OHK5Lwn9ixAgJkboWi8QJP6FI1+G20X7GB+IN8xhj2FmSMTZcfVMhsKZKsKAublwnjFWUE7z1c5+d4MNp/vrnyT1DbAsj1Z1ohFDD2KUPeb4g3DHeub95Li2z7vzF3DsdYh6IDihaZKdjtxTdaeXaXfbfbfddNi0u9+/yhjsX2RIKCLLDFqdYYbEoimy1O5En5labgbdyN9ldsNVJO8EzHXsR89i4t7Dy8W/cH90scd9Wt0QMFiwpWATAfcu9jEAdsk4IbMP/dvKsdRZZiLVNPfkRurlHETlTIhxECMrtRG13jVCdw3m9n3FNFqM5OiwEhIAQEAJCQAgIgcxCQIJFZvWHaiMEhIAQEAKREXDuOZybBrdSF9KO1boVLUHmQfqzShohgx/tEHqQi6zuxb81RCDnQqSFXCelS6wIaAqkCoQQdaSuJFZ2FrcEGUR92ceqeshTXKZQV8gXVm0TkPZUS5TDebSbjTJxe8UqZchTMOIZv7MJJUWsfblxkRK+RKH4A06Q7hBebssT7GKICv9aAG2Iayg/SF/uBSeAhYipNIkS20GIEgPB4UMwX8YqG/UL1StThYoIo5m2ePvbiUEuNg73LfsQPp2Yxb3HhjjhBAj+ungKTpCAdiUvxHA81g+cB3nKfcyY/NTSKEuIJtSBstiPqOEI1lQR9hHgib7bRA13fS+GG03IYDwwL7lxwfHtY4RSYwVNj1WhFLu+8QsLsS6f6HH/OPOT2rHI8kSvF29+b73cswRBHWsLjoUsT7YUKWpjr+iif4vutOtuWzftfuB/f+5WcuMPu++/Zf3vJlbgFmydjUjuleZ21u5bN4TujYOL7m/Puc1F/t36a5Gfix5S5EjbX8RiUBQpanIBJW6xWRcrCratJgUgXGyX82KPbOdekdOdWIFbOu5VLBkR/Hm2cq9gZcF+hGDuS9rKu0BE0TcCgNSQ94lO4XKxhGJD6OG+5PnMcx1RhPs+6S1WUO6kC9aJQkAICAEhIASEgBDIUARSsuojQ9umagkBISAEhEABQgDi3TZICRd0G1ICP9usu4TEwwUUBAJ/ISFYTcmKS/I5n+iIFxAWuQmqtQAAIABJREFUkAm4voCo+NcIfecOKG2Ihevvyqcd1A1rCdyjFLdEwFlIFepI3fElTlwA2oRwwQpQ6k1QVNpAGzl/WXgfAs0oS6zqJIgq1A8kDPjkpSiTNgwLc8EmWLjm51hN63amW7AozNjT9rAFBh+9+Od4jw5ba+wAVThOhiOhcxD1LjMuoSJsTqjlMGUwd7jrbl8JnsKg2oWyqwNWsIOzE50UtDhgVDhXR998U3an2n/NY0wiovFc29+o/90sHWehLDZuXVtkxdY/ixy40+FFzt76e5H/zK3Tj0X3s7g7u5mVw99F1phwcZi5eTrB0p72xPrLvElttn+UkcyGRQgC4+RwQlhkAQOWPdQRkYLnIs9TrEhCwm+ke9dfAWtzUJ2wHjrLEvF7ECYQQ1ycEp7FCBYurhQibjLt0jlCQAgIASEgBISAEChUCMjColB1txorBISAEMhqBJybI1YsYm2ASIErBwgHiHxct/C5mCVWyH9piaChxK+AmGAlJCuT8fWOgOFECgtwCp9fNC9XtXIthAhcSpAQKCA5IHsQJLAEIYAurjjYR71pL8FqYTsgKi+2VCKccEEBvUOQYIQPVuMT8wLyxLkcycv22WW1pRIBjyChfkwlsHGWZYSm27z4x9UXPjI0+JyuEUlM/9pyvwupOFugbAkiAO6B4lKC5RTY7M56qk6deU5a+M+saXj2/GFSj3mLMmFia5Fdix5pn7cWWWsunpYU3afIoQbqrvZEnmrixWFbfrP43L+YoPBPkQqIHFs32f9mlWH53fMZX0Y824dZ4plY2hJWlddbIi4Mz3UE/XcsEUAcQQKhCfHEWR8hGFBH9juR7694RYo4OpD3i88t8XwmPgbWRHzmWcz1EEsQLLQJASEgBISAEBACQkAIxImABIs4gVI2ISAEhIAQyAgEnHUEVhYQ+aMs4eoJ4YIEcQFBD2HAhrUFFgwQGxAGrLxkxSVkFKsuIRogWPJ64/q0BdEC1xmQKxAq+MpHdKBuHMdtFa6u+Iz4QB7cW9BGhBcIGIgd8iF6QJBgNeKOc46LhZHXbdT1hIAQEALZigBzdHJr/LO1xSmot8ctWBETL/4qem4otknIUmWnhqHPf5hLqJ144pn7p3khO8G/TLTYWGSsfYLYx20Tz3cEep5lJJ7ZWCrgyonjlMcznmcnIkVxS4gaWCc6KyQXhyQk+IUFx1yLfRGsI4gBwvsF18fagrqxYIB6s2BCv7dTMLZUhBAQAkJACAgBIVC4ENALVOHqb7VWCAgBIZDtCLDiFZKCjb+IDRD8CBNYVfCdeBVTLEFssMoR10i4f8AqA8KDv04ogBQJBQXOB2DcSmuuDdnhAp1CzCBYIK7gw5768Z2Vo9SXYKG0h2c4Vhmch6VFWUu4iEKcmRveDyZgsTYcWFwEXD50tC4pBIRAViIQlwVNVrYsDyodFi+IT7L9uWOfgwLNrze3aTynve7PeL7zbHwjvN+56MLVEs/vPpacmydnQeFicLjneZ71XzhwOXX7Nvzs5dq8j/xgSVaOeTDedAkhIASEgBAQAkKgYCEgwaJg9adaIwSEgBAoyAg4MsNZFTgXURACiBP4VIGsr2epgSVnwYAlBm6kIPuxxkDQwBoBN0u5CoSZCNjmciooOzqCC/QMwUG9IG74C8kB4cGqTQJqE98C64q6lrCoIP8yS7i3ahpuO0QOLqUQPQiUyoZbKZ73P9u1NuSx66tEIMqTvNNW/lG06jH75RmRlSeN0kWEgBBIBwKheSLFAb3TUc+CUKbf+sFZPrq/3tgxzl1XKD6Tp/H5Oq+HXWRtNmsL3lHYsOAMiTXOfVZB6Ci1QQgIASEgBISAEBACeYGAgm7nBcq6hhAQAkJACOQagXDQamdhAXGP+OCsJ063z/iQrmPpXEsQ91gnLLXkAqcSlBoSn5gRrMyExOcz1g2b8pvIJ45GuE64esJFFG4xqDuurk6x1DD8eUV4P840jrMESVPOEsIMq07BgHYh4CDKsOqTc7DQgEApkt9tpQ75sZlYQb+D60YTLcBGmxAQAkJACAgBISAEhIAQEAJCQAgIASGQQQjIwiKDOkNVEQJCQAgIgagIQOjjCgm3R8R6gMw/1hIWBggUiBYEvGRFI4S/C5j6vX12QamxqCAmBMdxl4TbpUxyk4QrC4h0BBlnGYIowWcCjXJ8jKWSls60VDtcf7eis3wYFwKTnmUJkWKiJUQNnvneVar2tVBuuATbw8QL+v43Ey4yqf8LZYeo0UIgvxF4/L1JQVUIzZeysMjv3tH1MwEBe2Z6q5EjIL09RzOhiqqDEBACQkAICAEhUIAQkGBRgDpTTRECQkAIFHAEnAUCrp2wrCDIJsQ9FghOgPjSPkPOF7NUxhK/sGGiiPFA7AesLLA4mGeJYJ6UsyVDLA6cmwtEFaxDcHOF8IAYMc4SRPsdlhApEDGIa8HGcdqCkOMsLdhfyxIBSSHmKZPgn2x/mzXHv9bmwkjU414E11pgAbYbjYRZZGQL40KbEBACQsAhICt0jQUhEEbAI1bwvkF8ERejI1/dcKmDhIAQEAJCQAgIgYKLgFuRWXBbqJYJASEgBIRAQUIAgWGdJVwbIbrXtHSepX0tQcoT8BIxYqwlrAt+tXSipSrhH9mIAAToJCg15eA3u2jYHVMm4MSPf+qElQUkOkIEVhW4MSI+B+6iqlpyYgV1xoICEt4FEnftgJynjQQkx/KEc12Q0kxqc57hHo5dASZY3SDwVLJUx8gYYpxoEwJCQAg4BBS/QmNBCPwPAQQ83jtOtoQ166GWWCiiTQgIASEgBISAEBACaUFAFhZpgVWFCgEhIASEQKoQ8MSu4AczP5BxC1XcEgQ+rqGwuIDkxycBJDQWCLhNwg0UYgX7scYgxkVZSwS0Jj+r7LEy+CtDLCwcZN4ViwgzuIJCdGgUbq8XWiwxsKRgQ+BAkKFt4IQlCUFJIRbA6itLiBgOx8JoYVEkLFqsMpECUQgrC/4Wt+8IPgQz346L3Fx4h5o+C4GCi4C5fQpqnFaPF9wuV8tiIOCzquBdq4El3FPyDsXiB3+gdGEqBISAEBACQkAICIGUISBz55RBqYKEgBAQAkIgnQiYcIHIjqUBq+FLWYKMx4KCVfKHW/omvA+LC8hnfkwfYQnBAtIfy4sjLWFduMwSrpKWk9cEC4j8fN3Cwoyrg7OAhBRAbECkoV3EpUCUqRHOCNkOgUA8DixHCM79tSUIBUQOCHiCipMIwg1eWBiELDIKqVuo7f1shAwrRolpgmsxhAqCk0+xlMNFlISLfL01dHEhIASEgBDIQwR8YgWLOy6xxHvIjPA7xKLwewWLAPKwZrqUEBACQkAICAEhUFgQkIVFYelptVMICAEhkP0IILJjQcCvYwQKxAisK7AggHgmfgN5WAkIIc8P6tXhPOyrYwmRAhGAH94uWHcRXEJlmJWFCxyOcIFLKNoz2VLjcLtxjcU+3GDh6okYF8TrQLDAZcNKS0dbIu4FOGBhwmfnOoqVw4V+9bARLb8bMUOME4QcAp0jaEHOgCdjJ4QR5I1IGZDQJgSEgBAQAgUZAY9YwbsS7xSPWDrJEs9KFoJ8aonFEtqEgBAQAkJACAgBIZA2BCRYpA1aFSwEhIAQEAJpQABXR8SrgHjH8gCLC8QHiH1+XLNhbYArJUQNYkDwwxprDKwMIKE5BuHPXwSO/zJMrHCwIVpg+cFqf6xKqDOr/6k3OOBHGsGGeAwQ6xx3G239IdxmrC3AgTwEyyRBOmzEqiND2+5pSno/mhBB4G2sb5ZZqmyJYO1XWhoR3ocQpE0IFDgEbNwzbzrhkr9ey2u3P7Qv7EqtwGGgBgkBIfA/BHxiBdaHd1tiEcQSS7jVHGAJV5Sh+UFCvkaPEBACQkAICAEhkC4EJFikC1mVKwSEgBAQAilBwBPDApId8hhBAgECQn+ZJVbGH2sJl0hYXSBQ4AqJ+AQEpIagJ+g0hD4ufyDvETkg/XkOYsGQiRuEAG2krViWYEkBsU7bcA9FW9hPuxBvFljCkoJ8Iy1xPpYnWA9ATCLgINiw0X7cZuW7K6xMAN5Ily1G1CDygB9YXWypmSWEMQK5Y93iFYQyodqqgxDYjkBYfGDsOndyHGOOw4UcogOCrhMsscxiHixhCcs05gFcxTEn4GKOOQSRFEst5qD/rHzmG8qmDPIzH7t5FFGVxPnMv64OnBuKCSNic3tX6YMQyEgEPGIF9zhWqddaOtfSz5YGWXrVEpaphTL+VUZ2miolBISAEBACQqAAIyDBogB3rpomBISAEChgCEC6QYRhVXG8JawLEDAgyCCbcecDOcePaYg08kOs4QYKN1KQd/zYxkIBso6yIN0y2TWSIwZoB2ID7WTVI+Qg3xFbilnCKuALS2MtXWEJgQYBh7bOtgT5QFkE4uYcsNC2IwLgNT2MKSIYmJUHcyNzwBexKCRwiYDV8Ek1Ah7C0Fu0m/f4y3s7cxtzFvMdAi33Offz2ZYQb0+whODAWGZeqGKJeY45gzIQMdnYF888gFDHXBtpY7X1J5ZuDGdYaH+5h+ZYYr7l87/WNgQRiE/mMK5NXRTgPgqwOiQE8goBz9zD/MK80s7SZeHrI2BgXcG7VqYu8MgrqHQdISAEhIAQEAJCII8QUNDtPAJalxECQkAICIHkEPBYWCAwsOoX8YGA0pBoSy1B3GFhwDF+WBOrgbgWkGGQdIgTkG6cPyr8GfKMLbQCOJPdIln7IRWxpKC9rJKGlMR6BGGCNkNilrXUL9zGpvaXlc6zLL1naZqlhpawwEDQ4NkPTmCzKZPbHu6jPPnjI4sZK4hfjCMIHGKHQNRAxhLAHSw3YJmRJ5XTRQo8AuHxx73J/Y6VA+POCa24wWOOq2AJ64iWlhDS2EZbYrzWy3CQmI8QLxA4lllijuI+Wh7+zHxE2wIFZAmEGd67ql5WIxCef3gvwKLiTUtYZLLxjHvQ0muWsDjcvumezOouV+WFgBAQAkJACGQ8ArKwyPguUgWFgBAQAoUbASPUAcB4ewu4sI00RnwgLsMBliDqIPgg8vGxjMUFRDPHIMRqh/9CjEHus7IXEhqLBfISbTuTLSxou3MLxWcIPdxC4SYKwhLyj9XUtJVjbMRewJUL1hSQ67SZfayOJB+khNsAN9Pb76lu+j5CvnhECzDHgoUxUimMN6IR4+o0SzUsfWP559h54KtNCERFwDO2vBYTjClECeYxhFbuRcTIiyxhGYH1FPc7YgVCZdB2apLQe2NWYI3RPVwPVlUzprmmf2PeQUhJZsMyjBS0cb/1sDTEEqIg956zBtP8FAfaEaxzOJPx5hI4O3dd4Eri+emdw9y4cM8GxSqIA/8CkIVxUNJSE0tOrKBZj1nqbSlHLCeJFQWgx9UEISAEhIAQEAIZjoAsLDK8g1Q9ISAEhIAQ2IaA6RXOPzs/rA+2BIGHOMGGiyiIFUd0sX+SJX6AI3JAyB1taVE4P3EwIMQ2mmCR0S4OwhYmtB1yE2EGlyqIDhCbfD/OEu5gxlsi3kIpS1hjkJ/A27hlwf887lhoK4sVwBDRZnMWCDbhLsu7Pz7yD6yw4qkexhW//4wdBDDGG65vwJkxFXEsFXaCx0fY5yBDA3rWEazukDcAtCNa3Tusl2B1+yBmvUS3EzYpzx3bSiBpq5e7lj/4NOe4enKOX9zLEZQ6fNwtBIIAdvEecGGHKME+7kGsJRDBzrKE67a6lrwiYrIDHbKfccj1GJPMB1heMU/MsMSYRRRBdEDQJDG2sWygroxdkotRQZux9CAPcw7tZV5hH/MO4mdNS4gqzCXfW0LkaGCJ+ZnrEcQegTjRBVK4XnvXEvM1lhmI0dQ7UBwsDPdWgAWYwRHqG/qF/qO/cPdF/7CBF/1CnzSyhLCN0D/FEv3GcwF3ifQNlorkpzzKQpRi7NCnHHPlu3JZNJBjrisMfRDGtcD9sbHF/Xy6pc6WcCPntufsw0uMG+bKAtdwNUgICAEhIASEgBDIaAQkWGR096hyQkAICAEh4BAw4t5LYrLSHXLG+WFHvICcgYRhHwIG+SGaIekgYiBYJljCRRTEDaRLxltY+FxiQSy4gLeIMgTMRYiBRIfYI9g22EA+sB/iEmIRchJrDEhECCqw+dfEClkHGBDxbGFiGzIQcQiSFj/fxLnApQ1ENGQx7rcIcu7iqmyPkZLthF6U+ApulTb3mBPCnNUT45VxyHfGoXNpxmpd7l9cjDAmIcKd5QH5ibkCjlgIuQ0suZ8h2DkPEYBxj3s3SHbqgas4zuc87nFIXCyPIFyximFjH33Fedwz9S1xT0GSu/pyfa7FNdk/MVw2+yhrTLhcrkd9EAkRR50YiEhQ3BJCKflPtgQJjHDANSCDI21YVHAdF2vC5QOzry1R728s4V4JIZLyuC5jkDmNz9QbAprNkc1bckM6RlnB71bsu5gUXJ9Ef1A38EbAoE1YvOG6ij5nPkK0QQiMtSEG9rf0oaVllhAKaev2rQDeX15LHD47XLlXGD9gyjOAccIxnn3PWEJI5RnnxPxY2HIcfBGWom3cR4w5+pM5D3IbIYk+pi6UwRh1z6ccz5Zs7594QMy2POFnGuPlPEt9ffXvaN97hPsacTfbmqf6CgEhIASEgBAQAlmOgASLLO9AVV8ICAEhUFgQCCDuIcogxSBQWFXsVoa6GBcQJhCGrGCG5INMhujiB3pIsMgm6wKfYEO7aQfCDGQVq2jdymm+49IBUgsBA1KVlbQQWpBKbqWkrCsSuHk8hC3jDFEIUht3PBCnYIyIQYLABmNWJiOQ4Y4Mcpb9iGaBK1XzmxCKQkiDkpeAxnLHWRAw/sAC92Ss2iYANCv7T7QEGc0xXBtF2r6yA8UtITwEbbgHQgzIxA1BhfZ5N8jaRK0lIHkdGzjIPuMrHnyrWuJ+RXzhWk6o4RiJa20fS/k9fmJ1UHh8ce+4scRfxGTwIlD485YiuYzyF8+4gVDFig4i/b/ciDGx6p6O4777zQkSzsIBEYL+Zw5nbCAKIPaclo66pKjMmVYOroOcBdpb9hlhgz6n/vTTdusm/zUzffymCKOMKSYsViDutrbUxlexi+37aEvMOyHhSf2TMV2niggBISAEhIAQKDQISLAoNF2thgoBISAEshsBj2BBQyC5XEwKSGBWu0OUOJclrDxmFTYEUHFLrHifbQkBA/IEch/BImuCJnva71zTQARBmjsXOayQ5TMkAwIOZBeEJ/khzyGMwCHkyiOb2p4JIzeA0AdXiEWsXCATIdbBnNXNrKbHGgP83Yp+VpUTS8S5JaM/HImXq9XvucXH2uZWyTsLAdoGUcp37pkLwm1DlOC+w10PRNadliCbvdtn9gWLAvLF2ig7nnyxysmU4wih3lgT9P0oS1hcePePC2P7nv3FjRvjCFGR5AQv2uTu7awnDGMIYow35m4EDMRX3NxdZwmxOdr4wKrkNktYniBGB7pkywSyNcL8wbOI9mENwfi4wpIT2XEXlooN0RrrHzZcPCGyTbWEdQRB3BGyscC7xhIENkIY3z8Pfz/T/jI/MC7nWjrJknM7Fat+3SwD1kxYYHBN5gae3bgYQ+jF6oo+Y/6LVZaOpwiBsFjB8+pRS818xT5i33EDhZC6/f1I/ZMi8FWMEBACQkAICAEhEDcCEizihkoZhYAQEAJCID8RCBP2rgrOmoLV3nxGsIB8gQBxvuIhDyF/3Gp4CGNILUj7kGVGNpH2nva7Zzd/nY95SCaILwhwxAosLMAGQg9CCrKJDQKCvAgW8kmd4ID2ko6OwAmT/RD7kHKQe/QJwgXjkXgFbMssQUpC3mF1wRhF1IDEY8wiNiGwsSIZawz60QXDDYqVQD86//XOyojruFgB7HPjhH1cC2KQfaHYJZZcGRCl1BfCGIKYxLjBIgmBAgEGAaI4FwhvrL5lXDX1XMcdm2wfnPslzymhj9yDkPOuHhDNWKeAAWQqGJK4NvctFixgAWbct4hD4MO9DbYIj5Csgy0RFwJrDgha5gTag7shsMbdiRM48dFO+8EPzMEB4pj7BosRyFrqwHeujRsn+hTXUAhTkOmIgvQdcQFgWhEd6Fv2Q7qDG/mpJ+IEdYCARpBAOA3dg7Y5AdH1ccR7sqAThgGEPmMWbMHb4X6rffbHw8DaAsseyHAIdcYR4ymjrE/C7XOWFIybOpYYr4zR88PjIZ4/jDHIZERoxiVu//iMKzGEeoQA7gvnJoqxxxjnL7i4ew/hwLlSc7GNOMdZ7oAfzxDmB84hL/c8z9r7LCFULrNUyxJjPpGNOQXBBFdrwy1xX3AvkGibEzIKjGCXCDjpzGvjkHmR+amLJeZT79bdvmC5xByYUfdPOjFR2UJACAgBISAEhEBmIiDBIjP7RbUSAkJACAgBHwI+wYLnl/OZD9lIghCGqIRshGiB2GQlJ5/JC9EDEQuZE/oxnk2kva/9oeqH20vb2CBwaRfkE3jwmfZ73RCFCKBsardvGGTsV4/LG+cyCvc2kOP47EeQYHy6cYmlRUNLWMhghcFfCHUIQQh33EhB1vKdeAkcR3SCJCQWAGOb8Ux5iAAuuC7kPfsg/XBPBckIMcgKf8hI3LYg4nGPEH8DQQBxgWN9wtc51/6yQSSy2h3inrHG9REXnG98yEYIeVwWUXdW7ELGu/NcYGbGIC7Z3P3Id0gz6oxgQB2dmynGKp+d6xjEDepLe8gHtiQn1nAvUzfIWDcfQHayQXizj+PefM5lE/sdgYwwQX3Awc0tzvWSs4LhumBBu5yVEwQrdXViEHlcuU4Ucm2hToVWkAj3ScQ/MSwwwJV+A39I1nMsMb4ZcwgajGe3IR4hAHBfOLI+zy1UAlw+cd9QZ8YnLniax8LEjmPlwD3G/UJ7mBdoH5+5/9kYg+6Z5oSJHYrOreAVXpXvynWWWPQJAgZ9wHxC/9AnrNpHxEA8oe7xbM41GgIhgcGZIxFhEDd4bnPv0J/bRQxvobltXzwVzOY84f7jmXK5JcQK78b4IZYP4hdjK8cmbLO551V3ISAEhIAQEALZi4AEi+ztO9VcCAgBIVCoEIhA2DvSHuIEYoS/kKwQXI5MhDRxqzbdavSsI+0D2k//O3KUz44shbRyhKqfIM26dmfLII9AuDpynRXVLuYFIgZjE5IPUQOinHyMW4hABIZPw2OZWBCIFpCTkO/EhYAgxFc8hPgZllgB7VZGR3KfA+mPMAL5iYDiNgQDykfoYHUtxCBkKsF12bAa4DN1JF4AljuQrtQRYpF6QcBC6jtXa856wOtuTUFbPaDrY+II+O4vxjvzPRZNT1jyBzHHQudZS7hfY5xuyivS1VdPJ3IRj6J9uJ6Q8LhV8t6rEMZYiowN30+IlNx73LfM5TzDHFkf6MYwr9oXqefClmbud6UTIREfmfsQOhFGW1li/kpkAy9i2WBNgkjazxLWS1hgIX4ylxLDJEeQ70QuUJDyBjyHnPtMnj/EpnjS195v7PvVlrByYZzleGfI73FVkPpGbRECQkAICAEhIAQSQ0CCRWJ4KbcQEAJCQAjkEwIxCHvIXAhTSAu3+tMRwdTYG/ATV1AFzh1SOCi3t3fcMz7rrEnyaYil9bIelzCMU1b/Q1iyMhwRgNXJkJiQSqwuhoxlP4QsbqJYGYugwTkQd7iAgazD7ZTbsGLgfDYIPVYmMwZw2cLGd0gpXCexQVQNtIQbGYQP554FAQRhg/vHxeFw1gaOFKTcHMSpiK3/dYQ+pR6BCIIg8z6WZSUs4XKLeBaIA2y4hkKIw43Uh5Z+tTHqxLTUV9BK9NSR+wOyHhdjWHsgqgRtCOmdLWFJgVjIfe0s4goUcWzY0FeOPGfewxVWS0unxegM5jksN7wb1lpfWEIMQdxl7sO6i/3OlRsWYfR3aJ4q6PNTgFDGMwYscKd2qSWs/Br4cMQlH0IaLve2W54WBrxijDkdFgJCQAgIASEgBDIAAQkWGdAJqoIQEAJCQAgkj4AvGLUriJWtkKvOAoP9IdcsBVGsSB49nZlXCEQgXJ2FjHNdhJjBBtHkdSHjgsdDzkJoQi5BiEJqsmIZYg5LCI7jioW4CazO5jPkoBPyEDIQNRAusKxAyPP6tXdBi3cQ9Ao64ZdX40DXSQ8Cdn9BhiNQfGAJ8cIb0B0ym5X6rPBfY2M5LYK1xy0c9cC1WpPwX3+jX7QdiIWIiIiDkPKBro7cidl+/0UIOs7iAuYx5kFc3eHuC8GUODoubgbxc5wbOi+OCKxOjPXuZw5bZgmhl7GACy0+M6ciYjAuQlaIhmmgtYq/szLhexSXabzrsPHsYNxh9cbf1pY4xr2AJR/zPFi77WH70N/SYsMhMFh9JrRbdRACQkAICAEhIAQKLwISLApv36vlQkAICIEChYBHuAhsl4SKAtXdBa4xUVxK0VbITPfO5tx9OTHO7Xfkm9f6wUuCZhVBV+A6WA1KKwKe+4eV5bgfYvX+tb6LQlg3sjTDSFrcoaVs84gVWHu8YQnrKP/2qu14yRIEuje2UIG3AIgFtMcCzcWQcW4eXbwdvp9nCTEDkRbBlZg+jrCPdQkXm4H4DcTd4byplrDEQbhFBKZPAuNkpFswikOQcDF6nPUd7aXeWKpwDFd/t4T3OeE7CJPRthOrni+sTYg32oSAEBACQkAICAEhkJEISLDIyG5RpYSAEBACQkAICAEhIASEgBCIB4EAwhd3ZgSVf8EScWO8G4LBFZYmG2kL6Zvrza6PtQCr2W+21MJX4Cf2/WlLBDXGDZQsmHwARSHsnRWaC7y+v52KlRjfiaeDZQbxPnC9hVUL1gWJbAhXuJIaaQnRF8sNXCWxMTY4xrWc1aZX0IhlqZPDLWO4TNceznVxpziEBYiLA4SrK8YJQgTiG20uaYlYILgPRLTBTWAi28uWeZQlrI2WyqoiEeiUVwgIASEgBISAEMgPBCRY5AfquqYQEAJCQAgIASEgBISAEBACKUMggtshhAtitCAaeDc3sPlnAAAgAElEQVRc5FxgaZSRt3xOePNcD2L5REsPWjrHUxBBjNtZ6m2JFf4SKhJGedsJcbjUg+Qnzg9EPv1Jf+Bqi7gNCFfEB8EKIdENt10zLSEgIGAgdhHMHSEDKw+uS78ifKy0hNUC+RAfOIbAQX1wz4e7JupX3hIuyjiP2EXUm4DY/C4fYumhcCW9bs0SrTdt72OpW7huuAPcnE1usBJtsPILASEgBISAEBACBQsBCRYFqz/VGiEgBISAEBACQkAICAEhUGgRCCC3WclObITLLCFeeEUFgs43tzTG0vaYBrFcAPnEClbAP2aJAN9uozwsLVj9vzFdcTMKbSf7Gu7rcxf/AqsXBCvcKOHuCSsFLDGwZsCVUlAMjHggRbDgGpQXtBFAnesdHj4YFDg8nuvEyvOOZcDChDgoSxhnlrg2QbQRRxBZEEu2xhrPsS6k40JACAgBISAEhIAQyGsEJFjkNeK6nhAQAkJACAgBISAEhIAQEAJ5ikDYbVNpuyjBhgnw7N2usi8DLOVwERWJ6PXEXCCgcVNLHT2FtbfPX1nCvRAr7At9jIo87egIF7M+Q7jCGgbrB2JiIDjwWxgLB0QsXExh8YA1RKZsiB1YbiCAbLD0liUECoSJdZY2WUKYYJwxdvMlBkemgKV6CAEhIASEgBAQAgUHAQkWBacv1RIhIASEgBAQAkJACAgBISAEIiBgpDW/fXDL84Al3DV5t0H2pZUlAjFvd9/kFy08YgXBn5+wdK2nkGnh73PtLyRzaNMK98wdkuExgYCBoEHQ9n0tYbmAJQZjhUDtiAO4aMKKhnwEr65qicDfQRtupGZYwoqDMov7Mg0Ln4vg8KUlhLTplggKjmXGGkuID4wh3FIxHrEYcaIE45h9oXGq8RWhF7RbCAgBISAEhIAQyFoEJFhkbdep4kJACAgBISAEhIAQEAJCQAgkioCR1KyyJ0Bzd0vEOHAbq9jrWCI48Q4uojyuhyCPW1qCYHbbCPtwuyVcBkUUPBKtq/KnH4EoQb+5uBMzGA/OxZSzaiAINrEqsIRATMD9FIIGrsb4nc0xNoQHxAnKYkMA2Sc8TjiXvJxPHrYc8U4kSIRR0R8hIASEgBAQAkKg0CAgwaLQdLUaKgSEgBAQAkJACAgBISAEhIBDwIhq4k+8b+lsDypT7TMr6SdbCrl08m0Q0pUsYU3htgX24SJLWFaIbNYQEwJCQAgIASEgBISAEBACuUCAF25tQkAICAEhIASEgBAQAkJACAiBQoWArVz/3Rp8gSUCb7utmn341lIzS1hSeDcWe5WwhCso73aHfclhWcFBrYwvVMNJjRUCQkAICAEhIASEgBBIEQISLFIEpIoRAkJACAgBISAEhIAQEAJCILsQMFHhb6txb0s1fDXvY9/rWvL+XiK+wYWWGnry4gZqvKW4AnZnFzqqrRAQAkJACAgBISAEhIAQyHsE5BIq7zHXFYWAEBACQkAICAEhIASEgBDIEAQ8gbSrWJVwCeXdatuXSZb43YQ1xgDPQT63NtHjxwxpiqohBISAEBACQkAICAEhIASyHgFZWGR9F6oBQkAICAEhIASEgBAQAkJACOQSAWJPTLdU0dKvnrJwD4WbqAMtXefZTwyL5yytyeV1dboQEAJCQAgIASEgBISAEBACHgQkWGg4CAEhIASEgBAQAkJACAgBISAEtgXMnmepuqVVHkCwsBhi6VzPvk72eY6loMDcwlIICAEhIASEgBAQAkJACAiBJBGQYJEkcDpNCAgBISAEhIAQEAJCQAgIgexHwBccGwFimaVTfS2r6fk+zj5jYbEh+1uvFggBISAEhIAQEAJCQAgIgcxCQIJFZvWHaiMEhIAQEAJCQAgIASEgBIRAHiPgEy2wtFhi6VBLr/uq8pJ9v8XSckvk0yYEhIAQEAJCQAgIASEgBIRAChFQ0O0UgqmihIAQEAJCQAgIASEgBISAEMheBMIBuL0N2Mu+XG/pKksjLD1v6Q9L211B+cSO7G28ai4EhIAQEAJCQAgIASEgBDIAAQkWGdAJqoIQEAJCQAgIASEgBISAEBACmYmAiRg7W82wTCdtsrTF1VRiRWb2mWolBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAJCQAgIASEgBISAEBACQkAICAEhIASEgBAQAkJACAgBISAEhIAQEAKFB4Fdd91tt8OPPPqYVLd4v/3/7wBSqsuNVN7+Bxx4UF5dqzBcJ5Px3GWXXXfd1wZXYegHtVEIpAoB5voSJUuXLV2+UpW99t57n1SVq3IyFwHNlZnbN6pZ4URg51122WUfe4EpnK1Xq4WAEBACQkAICAEhIASEgBAQAnEi0OLWu+4dM2flr9Gy9/r0qwm3tu3wWJxFhrK91uujYS907TMwkXOSzVu+crWa01b+sfXUsxqen2wZmXBe1Zp16vb8+IvxRW3Lz/pkOp7Nb27dljELAZufOOnahQeB8y667Or3Bo+amI0tZj654Y52HcbO/f435knS5KW/bHrqte59DzrksMOzsU2ZVmdIyH7Dx02r37DJRZlUt0ydK08585xGo2ev+MXWNByYSXipLtmFQDbOy9yTExav+fvAgw85NLvQVm2FgBAQAkIgmxHYKZsrr7oLASEgBIRA4USgeu26p67/44/fI7UeK4kKVarXSoRE38m2Kka+Rys3lWhXrFrjRMrb9O/GjaksN6/LuuSalrfwI3arbXl9be/1Mh3PyjVOPMkWiO+b3zjlZx/p2nmLwOkNzmty+FFHH5u3V03N1W5ofe+DCM6fDujT86pGp9Vq1uCkyi883v6e2qfUb9Bj4Ofj8tISLjUtyrxSShxfqgyWKwccdPAhmVS7TJ0ra9c746x9bJn53xs2/JVJeKku2YVANs7LvF9h+bThr/Xrswtt1VYICAEhIASyGQEJFtnce6q7EBACQqCQIoAYMWvapAmRmg8Jw7ElC+bNiRei40uVLY/LkVnTJkcsN96y4sl3QtkKlcg3Z8bUSfHkz9Q8WDbMmDxhfH7XL9PxZEx+t3jBvM2bN23Kb6x0/cKBQJVadeouXbRgXra19uBDDz/i+lZtHhjQq2uXZx5u15o5ctG82TP7dOvy0g2XNDzNDh91Z/vHnsm2dmVafRkf1CnTxkimzpWly1essnL50iX/Zvkig0wbh4WtPtk4L/N+tWThvDn//P33hsLWX2qvEBACQkAI5B8CEizyD3tdWQgIASEgBJJA4OhiJY4nVsHsKMICxAJFL1k4P27BoryJIJwze3pkISSJ6kY8pVS5ipVXGfvx+2+//pLKcvOyLHwaH1P8uJIzp076Ni+vG3StTMYTnI48+tjic2dOm5zfOOn6hQOBo44pVuKggw89bP7smdOyrcVnNWp6yW677b77O6+/+LS/7ovmz5nV882Xn2t08eXXZHLMmmzAvHK1WnWw+FowZ+b0TKlvJs+VPGMgbTMFK9Uj+xDIxnl5z7322pv37rmzpk/JPsRVYyEgBISAEMhmBCRYZHPvqe5CQAgIgUKIANYVNHvW9MiWEKXLVary3+bNm5ctXjg/Xogod6MtHzM+Yma85ySbb6edd975hDLlKs6ZPiWrrSvKVa5WA7db0axdksUokfMyHc+SZcpVoD1zpme3NU0ifaK8+YtAhao1Qy7n5s6cmnUiWfnK1Wuu//OP33/8fuXyIBRHDP54ALFgylSoXDV/Uc7uq1cwNy8rl323GKwzpSWZOldCNCOmLDbBLFOwUj2yD4FsnJcR6nCZqveX7BtvqrEQEAJCINsRkGCR7T2o+gsBISAEChkClarVqo0YMW/WjKmRml62UpXqy75btGDTpn//jReeStVq1qZMyo73nGTzHVeydNnd99hzz2xfcV++UtUaYLx4/tx8JXEyHU8EtJBgMSO7Bapkx7vOy3sEyleuWmPbmMs+kcwM6A7eYlsk1HAPdU2T+nUmjP3qi7xHtmBc0cLp7FfsuJKlMm18ZOpcWbZS1er0/KJ8ftYVjNFXeFuRjfNy2QqVq9Fj2Sh+F96RppYLASEgBAoGAhIsCkY/qhVCQAgIgUKDAKtCsYLAGiKo0aYD7EUw0YVzZ8+IFxRiVxDDIprVRrxlxZOvTEX3AzC7XQThRmuR9UUiwlA8+CSaJ9PxLFWuQmUwAqtE26b8QiAZBMqZmPiH+ZtjBX0y5+fnOdTbFrP/H6JupHrMygA3dPmJUW6vXbZilWpYx82ePnlibstK5fmZOleWq1glJFgsnDsr7veKVOKisgoGAtk4L5exuULvLwVj/KkVQkAICIFsQ0CCRbb1mOorBISAECjECODXvEyFSlWjxZkgYCcugubPnhG373ZckHBOtLgYqYS9XMWq1fEdbhYWWe0TmIDbc2fkv8uZTMezrPU3YoWCtabyLlJZkRCAiGYeZPU880y2IbVkwbw5tME05ErZVvdsqa9bNT17+pSMEiwyda7EwuKv9ev/zEYBMFvGZEGvZ7bOy4h1i+fPm633l4I+QtU+ISAEhEDmISDBIvP6RDUSAkJACAiBCAiwkh7f5bOiBNyGROd0EywiuozyF1/R3EGxL69iMdjq1urLv1u88C9zHp6tnX3QIYcdfviRRx+TCYEYMxlPxmvJMmUryB1Uto707Kv3UccWPw5/+7OnTZqQfbUvUmTi+NEjqXftU+o3yMb6Z0OdS1v8j82bN23KpKDsmTxXsjJ+wdyZ07NRAMyG8VgY6piN8/Juu++xx3EWcE3vL4VhhKqNQkAICIHMQ0CCReb1iWokBISAEBACERAgzgSHZk+LvCo0mdX2lLvu5zWrIwV55ZrVa9c9FdIit52DJQfBYjPNd3ii7XLBz+fPnh63MOS9RmHBExcnEHHRxmyi2Ct/4ggcU/y4khdc3rxl2bA7tsRLyJ4zXDDqTFs9Hy+C1PuXn9euqX9u4wvjPUf5EkMAS8WQ1dfGf/7xn1n8+BNK16t/9nmJlZj73Jk6Vx5tAqB5KDtg7ozEXDim6hmXe2RVQiYgkI3zMvPEzrvssku2v69mQv+rDkJACAgBIZA4AhIsEsdMZwgBISAEhEA+IUD8CqwSli1ZOD9SFQi4vWLpkkWW7fd4q0m50Qjlppddc33XAUNHvdbro2HxlhkpHwGiibORab7DE21X+SrVam4LuD1vdqLnZhKeBx96+BEHHnzIoYm2Id78FW1skTeaVVC8ZRXkfCeUrZBW9z9Xtrz1zgeffvmtPkPHTun16VcTjjqmWImCimfl6ieeRNvmJEiwZgoeW/7777/PBw/sj1urgtxP+YU38UFK2HPISMjJ/jqwmvr9z8fPeLnHgMHEdcrLOuZmrixeslQZXEamo74u4HYiq8xT+YxLR5tUZt4jkI3zsovdMifDXMflfe/pikJACAgBIZAfCEiwyA/UdU0hIASEgBBICoEKVWrUsh9OEf2yIwQUt4DbiawGO/yoo4896OBDD4v2g8wR2kujCCXxNsi5rEqkjvGWnZf5KlateSK+5pMJuJ0peOJTuvuHw8dcdu2Nt6cLu4rVatWOJbKl69rZUu55F156Vb/h46btssuuu6arzk91uOf20ysVP/jpB+9pVbJ0uQpv9P1kBPNFuq6Xn+VWqVn75DU//bBq3drVP+VnPXJz7aED3+/N+Y0vuaJ5bsrRuTsiUKl6rTo72WYxlHYQLPbdf///wyIMwf/nNT/9mJf4JTtXYgExYMQ3Mxn36aivi/eRyDM7lc+4dLRJZeY9Atk4LxPf7Z+//96wZNH8uXmPmK4oBISAEBACQkAICAEhIASEgBDIAgT2P+DAg6at/GNrq3sf7hSpusSiIM9lLW5qFW+T6jdschHn1DnljIj+0iG2WW0KkRNvuZHyPdDphdcnL/1lE76Bc1tWfp0PHqNnr/jl4Wdf7ZpMHTIFT4g7+r7+ueenzfXMJ2OnL3qjz6ARyeBUWM55vffHn/U3wjGv2otrKPr94quvvzmvrplX10GEmbR03b8vvdP/07y6Zrqu099W+n8+ecEqXJKk6xqFsdzb2z30BOOf2D9B7T+6WInjscLIa2ySnSuvu73N/VNX/L6Fd4R01Pm19wYOHzVz2c+JlJ3KZ1wi11XezEQgW+flj0ZOmtv9o8/GZiaqqpUQEAJCQAgUdARkYVHQe1jtEwJCQAgUEAScZUI0v+xlyleuSnNnRwnK7YeDcgmkGW31JMeXLEzOmmDH61WvaUUF+g7Plq4iHgA+vZMN2JopeNaud8ZZYD514vi0/CA/4KCDDwGrWdMnZ2Xw47wYj1hVVK998qnT0tQHQW0Y8mG/Xn+tX/9nNJEyL9qejmtg+QSmC+fNmpGO8vOyzP69unU55LAjjjz97EZN8/K6Bf1aVWvVqYvbLbOQC3Tn9/3ypUvMwOK3vMQhN3Nl7Xqnn7V08YJ5v//6y7p01LlM+UpVE40Hk8pnXDrapDLzFoFsnJf33meffYtZPJtEx37eIqurCQEhIASEQEFGQIJFQe5dtU0ICAEhkGUIRHMJU75StVDA62ixAAgQ+O+/GzcumDNrerxNNy6iBjEvjJ/5NegcrCqw3Ii3vGiWE/jYJrDonOmTJ8ZbXqR8rDpmFWek47vbkj4CY6fDD7kTj+bOmjYl0XZkEp7mxr3CD9+vWPbrup/XJtqOePL/L0h83ggWhx1x1NHx1CuZPOkq+9gSx5/AfZFqUoRyI7WTOYI4OAUxPkKVmnXq0u54YsvEcsG19z777pfMWEnVOUM/6vcewtIlV19/S6rKzLRymMPz0oKE+Zf5e8Wy7xZzH/jx4FkXbVwkOyZitTM3cyUu3lI9fzhcEMxw75RIDKJYzzjccRGzp5y9e6Qr7kamjfNMqQ9zPmOcBRd5WadE5uVE6sXcwbteIue4vNyT0cYf7qAYq3OmTcn1+2oy9dM5QkAICAEhIAQkWGgMCAEhIASEQMoRgNwkwO1nk+Z/P3bu97+93X/IVzfeed9De+61195BFzvjnMYX4BIGVyYfjpw4h7gS/nwEeV7946rvo/nVLlOhctWFc2fPIK7CQYccdjjulzBnxwVGkDsnfrCVq1ytRjSyg/gG7w768hsCwEYCih+NLVu1bf/F1EU/Tli85u++w8ZO/b8DDzrYn790+YpVIIO85AfxM26++/5HcK9Ur/7Z58XqDMgZXOhMWLTm76/MTUXQKnH2gT3BhT/4csJssI1G4Ma6pv94OROPWKEL1omem5940t9tH3m6M8HTX+zW9+NaJ596xh577LnXc2/2+oD01Ovv9Gtx6133JtqmSPldkE1IV9yKjJu36vd3Pvp8XLzkPwFwuY8YT+9+MvLb8y+58tpI1ypVrmLlod/OWe4V1yAX736o0/PDJ85bydj0xuqAiLjwimtvYHyMmrV8XV6WTXDdV9/9cChui2gfbeL69MGzb7w7oOMLXd7JjdBGvw4aM20h80EkvBAojbsNdPFmXNaBt7bt8Bj3PW6J7rjvkScjuYPjWh2eeulNL/HDvX/vo8++/NiLb/ZM5X3nb8tJp9Y/G8ze/+zr6V36DPqc9jo//ovnz5kVqe3xzLfUe+SM79acfPpZ51LOTjvvvPM1N91xD5gwp556VsPzU3WfRCpnw19/rR8+aEDfmiedcnq8OOZV313a/Mbb/HMFJPSTr3bv0+ahJ1+I9KxzbaWeDz3zytvj5v3wx/gFP67n+ZFqPBmHt97T/tFuFqeHZwBjmucoBGfQ+ChbsXI1+rdZ85a3BtUlmTERbzsTmStp1zNdevZ/pecHQ5jHsc5AhHHzR6dXuvU+rcF5TVKBJ4sgKGd2eJFBg8YXNuNeY+7CpWDQNaI943i3oS+YV3oPGT2J53Q8z/142tL6gUefpv/een/wSN4ReM6BEXXt3L3foOff7v0R8+vFV113k7c87q/2T3Z+I9o19tp7732iLZCIp34uT26ul+x8y/z93FvvfTh4/KzvwOiLaYt/4p00kXrHmzfRefmqG267K5Z7Qqwdgq7P85P3a3eM5yb3Bs8E3imDBEbun0eef737+AU/rf/W3lefeLnre0F96xamzJo2abuFKHNcu47PvHTvY8+9kptndLxYKp8QEAJCQAgUbgQkWBTu/lfrhYAQEAIpR4Af8fwgx43HJwN693j9uccfgqC9pc0DHffae98dfnRde8ud7fgh/beRU/3eefMV/GffdNf9D/srxo+naMIChBor5slTvGSpMv2Gj53a9LJrrof0vb7VPQ/cfu9DT/jLhIAxTnd/R0YEgbFm9U8/sJ/AnkHHISohBSCDzPPP+I/69Hgb4vCaG1u12aENZvHAPidYQC5CGNPeJpdefV3n7u9/UqNOvdMidQrHECGKH3dC6T7du7z0z98bNjzwZOcu3vz4Sn6s85s9/9u8efObLz7Z8avPBn98QpnyFe97/PlXU9XZ5SpXrUEQxo0WjTHRMvMTT7ApW6lKddx18AMdn+cbNvy1/oijjy3GWChhAdsRuhJtU6T83AubN2/ahBDyy9o1q0cMHjiAPr+t7YOPx7oGcRbe//zr6Y0uvvwagnYfdMihh0Hkn3LmOY2CzsWaBhHCtLrQqmlWBfcc9MX4q2+4/W6LvfzDHnvuvXdbIxoQvCAR3+z36Zf3PvrMyxCXfxszjLgXaWV1qstG/INIQVg0ve5wMIJE5d7HBQXj23S9pANwb7ENDI6KcM9yzPi3fX/7Zd0OfumZZz76avK8G+5o14E5ZfPm/za3uO3u+4LmD8rh2EVXtrixxAmly/IdbN/58LOxxNGh7yBUY/V1oscRSCG7EcFYAW7ecGZTbyMlP6lsY86mhb+WmgVJULnxzrfMGcxt3CvcN116f/z5XR0ef/YAG1dYpZnVQ57E//iw9ztvca+CcSyc8qrvuE/ubP/YM8ROcHXiHukxcMTX5zS5+HIISI5Hqu+hhx95FPP4OU0uuXzwh33eXTB75rRbTFg44uhjisVqY7zHES4JRH1Zi5tb/bTq+xU8XxnTiGuUMXfW9B2s49b8tO1Zd0yx444Puk6iYyKRdiYyV/IsPvyoY479zx5yB9rESF153h15TPESofnD5nF71UiJdVDpctsWKvBecc/DT7349Os93i9lUbjrntGg4evvffwZCw78WEV7xt332POvFjuuZCnedfp2f+NlYoU89VqPfqmIj8U8arfsHvtY5HTu2z///P13MOL+5bnG+8OZ5zW9+AB7OHjrzJxwhOEZaWzxPvP55IWraHO84y9avtxcL9n5FhGJWFUjh3868K3OTz1q0PzGO2kk0SmZdiYzLzOX3Hx3+46mR0Qcr7wLjJ276ndEI3+9sNJx+xCR+wwbM4V3hL333W8/3intURp6LrmNOabPkDGTGzS6sNngD/v2+nbsVyMaXtDsyqCFL+VtTvvl57VrsELlfETavkPHTOHZBp7dPhg2Oq8tVZLpF50jBISAEBACQkAICAEhIASEgBAogrk9FhWs7vISv10HDB318eipC/wQsQqS4J+sRIZs5Tir4Fh96M0L8UG+aKvfS5haQR6IrYGjpsznehAbrHQdOf27Nd8uWr0BAtJbLj/UOIcV35G6jx+55EEECcoDiUzAT4gqd5z2Ymnhdw/F6lvwgYCD/Pl6/o9/9hs+bhqiCivkuQ6ESNB1jrTGEOgabCBFycMPR87x/mhk9TT7zm16yRWuHFbZ3tD63gdTMUTpJ+qdbMDtTMGzqrnOAadIAkBusYKIYMyRIDNdeQSWZXxGK586UTesKpy1EeOYVaEv9xgwOOhcVj1yDvcKfcQq2ynLft3sxuUd93d8iuOMA0Qy7lEEAsqCiOaYG1f+8tNZ9pt9P/miz9Axk3OLt/d8MKM9V7a89c5I5bLSlhXZOc478uhjsDYB52onnnyKO8YKZe5bv+se7mP2j5mz8ld3DIGC++O8Cy+9CkGBehDHJJXtYwU5cw6CrCvXBZDnesw/QdeLd77lXCyRJn7380ZW9rI6m7EEnrSZsZisG5JkcGCsModHc510eB72HQQuOLvA5ohvwybMXTHQhK5Tzzq3MRZNrJwPaivzAmIFlhXOAohnAeUxdyeDj/8cymX1NPcV1gccp99Ycc91SEHCOPd/tGD0iYyJRNqZm7kSEYZ7IVlXVbHw5nn86dczlzRpdlULsMESBiyb39y6Ld+9opUrK9IzzuHrrMrIT17eeWLVI7fHEeSx8GPMelfTgz1j5fLrbr4j6Bo8S1iAMmX5b/9xj+W2Hrm5Xm7mW96beCd0bed9jvmZ96rctsmdn8y8XLnGiScxjrBcCKoHAgPvELw3+I+z4IJ+aXXvw50QKLFQ7jN07BTXJnfvu/MQrnj2fzVj6VoWLrCffZQf9Mz4fPKCVSyiIR8WkNSTd1gsNK64/pbWfL/k6pYF1l1fqsaFyhECQkAICAEhIASEgBAQAkIgnxHghyCm6fwY8ooVkFsQX5Ci3iqysjTTbrsAACAASURBVPDLaUtWQ9h7VxdCqvCjy5vXEW24A4jUTFYO8gMKlwcQ+94forif4djBhx5+hPd8VkzyIy9a3AncSfFDP8hk3hETuIzxlgt5eHWAhQUkKe4k+JGIyxoILq/Y8M3C1X9BUge1ERcPEKFev/sIOLTL6y6AFfXsg5BPx5AobitYnTCUTPmZgqf7wZ1KiwovHhAI4OS3FoLIhDSIhB0r5rmHIIn8biAgmyARgs7FYgKRDFGu2TU33Mq1Went8uIain3cixCZWBa5Y5By7I9Up3SWzb0ayx1JouMMko37mjYHnQu5Ccl5W7v/WbqAG65zIO8cmePO5V4GO79bIgQf9j/+0tu9yFu/YZOL+M5fvje+5IrmfPeKH4m2xZ8fkYIy/XMO+ZhPOMY95j8vkfmWcxmjzOesqvULsrltgzsf1zQQ/LHKgxSmXc49lT9/Xved6wMnGOEehWeEs8JDxEbgCXpmuLac1eiCS1w7EMxpXzxYxMKKZxnPFoQ35hJv/rMbX3Qp15m89JdNPIP8ZRG8muNlK1apHnSdRMZEIu1Mdq6kji907TMwlgAcC7Nox2kzoiqiJK6+XF5EaLByFiveMiI943C5xTmILLmpU6Ln0tcDvvh2Fs8ev6tKJ3R6RXVv+W5RB+9QiV43KH9urpeb+RaBkH5MRRuCykh2XuY+4b3OLdjxl40lHWMGqxT/MffOi+XLkG9mL8XFWCTXUZyLm0LKOum0M8/xloUloN/FnxP9sU7meThhydp/ECvcnIY1W+g5ZAsh0oWpyhUCQkAICAEhIJdQGgNCQAgIASGQEgQgSVm1+dSDbVutMx80rlBEBgSJSePHbPezyzFWKOK25on777wZ1zDsYwVtyTLlKi6aP3umt1L43cbFwdyZkYM8Y2HBOac2aHj+4/e1vsmZsbNv/fo//gj9NT8AOcq1H12L5s2d9e/Gf/6JBAJkyuxpkydyfW8e3KXc88hTnYmr8dZLTz/mPTZzysRver31Sg6ylLYiNuAP+PZ2Dz9hXNLRbW686iJvsG/zgrObef/JUUfKhUjCZP9tu86qlcuXumuVNv/atJMYCW6fueb/hc9BcUBS0dG2erca5dDGZMrLBDypd4UqNWr9+P3K5d6xmkx7Ip2DYEScjw96ddvuG5xVnVhATJ/07deRzmvzcKcXELHat2p5pbdfyW/eq/6MZAUBqWBeumbh6ggifuLXo0f27vp6Z3cd3CyF7oE//vj9zusua+IdZ8eVKlNu1fJl30WqU7rKRgCgrbOmTgoU6ZLtD1xC/fTDqpWHm5+ToDIgiCFepk38Zpw7TjyParVOqvfi4x3aLl4wN4egBO7k82PvVsiPG/nZUOa4Ng92ev6zTz7o9+XQQaEV07GCWifaPrC60/zUE8fHP+dQ1p/huWPqhK/H+MtOZL6F1MQ/+Xc2oFrd93CnHl06PzN80Ad9E61vtPyM0Qc6vdjFK5xFyo8rNY5FskDI675zcQ2+/mrEMKzjml3T8tbOTzzYzqbi0D0U6ncbX/72MH6uu80ISjvPtYk8pcOxVhbNixx3JF7sITa5r7q+/Mzja1f/GHLx5DZcBPHZnqOTzZvfBn+ZFavVqo2bP6tHjucv+RIZE4m2M9m5knpBtKd6/nC4IISBZdUTT6r3w8rly17q9ND2+Eb2yA2/U+z4vI70jPv91/Q+myONkQ5PvfzmcfZ+9IA9U/xu8IgdEopHFdDntN9ZZuKaLd4xGC1fbq6Xm/n2D3svwo1YKtrgLyM38zJ4LJw7a4ZzY+gtm/dFRG9cfeFe1X/d6rXrnsp9fNKpZ57Nc//ulldc4H9ncOfwDGeewiXW+FFfDPeWNfiDvu+OHjE0ZEnhtopVa4asjudMnzLp0Rff6MH7Qce2t7V078Eu/lPQ+2o6MFaZQkAICAEhUDgRkGBROPtdrRYCQkAIpBQByLob7mz34PjRX34GYectnNVc/BibYfEd3H7ciTRrfsOtY7/8bIg3ADVm5xC6/IDylkGQ5xVLlyyK9uPI+eqdNN6c8oYJLlfGPvvst5+59oeL2U7S8GOcH8BzZ06N6I6GPBDbM6fuSM6zog4XCa89+1iHIPLHD7BzO7XBmA78/772zGMdIARdPspCsFmxdPEOpv/X3Nz6HoiGvub32uWH/D7z3CYXDf6gTw6sjKj+kh+V9eqfEzOAdzKDADyMF/3NT+rGU1am4Eldq5140ikzpvxvTMZT/0TyWPn18BO/7uc1qzmPvm1vBC3imF/McuWygvSshk0vHtjv3W6LAoIm77nX3vtstGHsrwdkIoLY/Nkzpl1z8x334Ou60wN33eLIBa7tgjF3an/3rWuMzXdl4DYCcnp6BCzSWbazPEhHP0AwRnJhcsqZ5zbyzkmMSwj9pYsWzPuwz47EnBmJhXyH+7EvXb5iyL89cw5+xsHq+Ufbb49dY6F7QgTZ77/+si6RsRMp76XX3nQ7bkDeeOHJR4LmHDMgOwpf/tMn5xTEEp1v3Wprw6nxOou98sbznXaIKZSb9iAw4FrnyfZtbhvy0fvvxSpr5bLvFiMG1Kp7Wn1/3vzoO+IaLFuyaAGCwM133//IgjmzphO7aPtcbv0OQeoXuS8yixJWQBPXyfssJN4RIpNXZI+FSdBxyr76xtvvppz3e7z9mj8Pz1b2Tf523Oig84l/MsfEDAhS//FExkSi7UxmrqR+zJdYkaRj/qB844uP592G9ITNp15cXMwBt0DA4RXtGUe/fL986RIshVIVwDrWOMGKCfd0zBlTAvqdPl/+3eKFQYs2OA+LSt67eFeLda14jufmermZbyeM++oLxCe/lVw8dY6VJ9l5mXIr2YIY/wIdd70b77rvIcTPCWNHfUEsCX89eKdkEQ5CBEI7i2ci1fXGO+8NzTkvPtb+nljt4TiiG89I4k2VLlexyoN33dTc+8xx8aF4L4+nPOURAkJACAgBIZAMAhIskkFN5wgBISAEhEAOBM5uctFlBJ/saStx/dCcfHqDc5fY8j1Ibnfs9LPPa4qLkn7vvLGdgEfYuO/x5179dECfnn5rDIK8sio0GuwlSpYKWVi88UKnR/z5IBL9K8iPt5WxuEqIVi6r0iB/CabtLxPRASLys0Ef5hBoItWxgv24hMDC9B48elvQbG/eE8qWD/kwXjh39g7xO06se9qZA/v27OqCXLPyDtdZy5cuXsjqZ285P/3w/UoCKZ5xTqML/D6MUzFsXfBzPxkXT9mZgCf1xF0YgeC9K+zjqX+8eSCjqtSoffKcGVMmcU6I8Hr57fdYwf/QXbdcC0EUVNY1N7VqU9R8Q7z75svPBR2HcAwiv50LI8bVZUZqD3i3WxfvNbgu9xuk6BdDPs4RtwHLHeobtCqfOqSzbOoFERMJj3jxDspn98GKw47c0cKCtuJibrJZfBHMnHPPNBdOuPN516yiWG3sL++QI7YRvX7sIa4hIX/7dd3PLW67675333zpOe+q9mKmonKfmFHUkty0hXMRnZhzqPPgD/uFXFB5N+Y4xvS82TOmWgz19d5jic63xNPhfASfV57u+ABib27r787n3iMWwgfvdX9zQK+uXeItd9qE8WPpI79FRl73HeMHfBCxQ6KxuSJ84bEH2nhXSGPNhMjibxuCPNYA7pnD84c4Krile6rDPbfHi0WkfI2tfPBBPHFWi968zjIkiLimXZCU3oUF3nMTGROJtDPZuZK6MX/wN13zuLPaZCGG34rDuVZaFbaqcVhFe8aRBzGa+7Re/bPTsqDA22e4oGrb8emXvhkz8vNurz7XKWjcsBgkSBzfFgz6gUc459sxI0cEiVjJjNfcXC838y24U18EnGTqHemc3MzLzIWMI6x8/eUjFDW68LKr2R8kFuFCyoxmKuDm9LvFC+YFWWC4MnlvwH3pOLPsclZgsTCoWKXGiYxtBND+vbp1mTNjauhdxm0WeD78vjorx/tqrHJ1XAgIASEgBIRAIghIsEgELeUVAkJACAiBQAQub3Fzq0XzZs/EDY03A4QO5LqfBKlzav0GrDz/dtyoLyBS8TX/Ss8Phkz6eszIR9u1usFbBj/qWFUczRIC0sPIwVKskA5yD8GquoU+N1POT3c0wQJ/yxCOfvdHrGwrcULpsvxIjJfM4wcgZRFk8Wlzm+UnRl3QRdwDeNt/Yr3TzuTHKSuR+XFMUPH3Px8/nTy3XnnB2X9v2PCXv1MQMVhVTZyGVA5ZSAysUmZNnZiUC59MwBM8nLXBtInjx6YSH1cWRBdj1niE2ZCs3T4YNrru6Wc3vPuGKy747NMPA4Oq07dnn3/xZRPsnghatYjoAYmxZOH/rHK2kwflKoQIZtx+0EfdXslJTrnA291fe2EHf9PEW4BsHTfy80Af5aXSWDb9MG3S/9wypbIvflq1cgVkjjc+DuUj/hHI1EvwnGfEEK40hg7s3zuoDgRFZpWx1zKFfKz4xWVGg0YXNDPueS+/5czxpcuWR9CI5nIu3jbjOgQrmhEmODnh0nuui1kTREYnMt9SJu3lL1YEzr1VvPWMla/5La3b4vruzRef6hgrr/e4s0bzr5DO675jVT8i9pzpUycRLwhxePI3Y0e5unLf00+QiN76M+aKHVeylLMowVXi+5+Nn17zpHqnt7nhiguDSONE8CEvLrN4xgz5qF+g1YpzvTQ94J4rZnMLrm0iCRbxjolE25nMXOlwYf5ARFzqwzpR3CLlZ77l2KD3e3X356Ev2bfQ3nu8xyI941weXAQiOra49e77UlXPoHIQrp55o9cALDPb39HyqiCXQ4xjXEfynPKX0eTSq1q4OGCpsmDJ7fVyM9/yDjfVnvcXXtHiRm/csNz2QW7mZZ4PXH+JzwUh+4h9hbUOn4PwP6b4cSV5x+N491effzLaAhIsZSjrw97d34ynvbyLIHbx7r6zfXn92cce9J/H+yrvnlgMxVOm8ggBISAEhIAQSAYBCRbJoKZzhIAQEAJCYDsC/HAqZxYQbgWbF5p6Z2xbRej/wYUrmNnTpkwk+OSwCXOXX97iplYQWHe0aNbYv5LPhIVQzIR5s2ZMjQQ7K6lZrTrB3CH580AwIYr4LRcol1Woi+fn9FfvPb9S1Zq1WbXud0V1uhFD5Pv804/6xzMUEFTKV6leE+GBFe78cPafZ155KkEq+F0tgRXiDqtjCaZKkE/zQfzZ5efUrRbJBcDEcaO+ZMU8AXMhCeKpYzx5iCUCzjOSjF+RCXjSTny106fJuLWKB6eqtbYFPMcapf+Ib2dCJlx2zslVR48Y9mmk8ytXq1UHIiUSQQwRRgB7/0pHysOthC3yX1v3jLMbvt/zrdecGyqOQWo0aHxhM8aK33c1Y+Nks2zi/uT8oLqlq2yIXeaOGVHiecSDdaQ85q3ne+43fywXBD/EiS+HffIR5yJo1DZRcNzI4UOChAWCGFvX1CN+jpcUwk8/K1cXmN8vC8p9NyKh1384pE9IKPUJkMm26aRT65/NuSMizDm1Tzn9LI4HrTZPZL6lDCPSKvD3/R5vvpqMJVWkNjIPnnXeBZew0pc4HIlg8XM4LpKXbMyPvnMri7mfGl102dVdPO6dQtjZRM5ff78792d/m/kLwd0JZI/wdOV5p9VE9EgEi6C8zMvMOxZvacJPq75f4c+DBSQkIwR7kJ975mbOiUROxzsmEm1nMnOlaxsWIVg/pnKMenFjwQXfTUTe4b2ibMWq1ek/v7gc6RnnyiVmVe+ur3VGbHEiY277Puh8Ar9bmKxj77u1xWWR5nbir3BPLv9u0QJvGYjeBIN2ZPTMFMUYys31UjHf4toOt2m8F6UK89zMy26uWObDn3Fnz+xLwR83TH5RjLo7y0ee9SZih2L8RNp4X0Uk+9oXuyJSft5FeW9A5OhimHmto9055FlsbiuDhLBUYatyhIAQEAJCQAhIsNAYEAJCQAgIgVwhgD9mChj1+ZBB/oLObdrsCvZ5V23i/oJV56eedW7jG+5o22HU50M/ueDU6mXe6vzUo0HuWFhVByGBf/5IFT22RMkTOIaFhT9PzZNOOZ19EDneY6Ws3MXz582O5uoAa4igAMm2Srs+P+Jiualy1yt+fKkyrHjEvzwuVoLaUcqWtEF++H3T41oIsunxl97uBUnW8pKGp7W7pXkzb7DuoPJYZY9Q0+TSq6/LVQd7Tq5Z55TT6Qs/lvGWnwl4UldIeFZcpovoqhp2VdLUsB/8YZ93W1zYoG6slYgIEtTNb6XksHX32dgvhw/2412p2ol1IHQOOOigQ3q9mTPYe/1zG1/I2PtiyKAP/O0lRgHERLRV9Okqmz6gHf54C/GOpVj5cI1GniOPKVbc5WXeYRX6x+YexN1nzC+IEhPNuiuozBp16p7GcT/uzkWOxTrdj5XICEXe84+15dkQ6qkSLLge82MQoYwwg6VMaK71xSJJdL6FrDT3emUQc4d9PKBPLJwTOc6KXdzUxTtvesvew9Q6vm+yirn9+dF3zuIIwtlChYz2xmCiXv8TLHK69mMe5zhEMkLXw3ff0uKyc+tVQxBPBMNIeSGD6bspAQHXOYfxATltBP/XQWUwN2NR4w/KTN5ExkSi7UxmrqROEM+0eYYvXksqsHRlIDhC9ge54WNeIN6H/50l0jPOW68+3bq8xOr0q8zdTirr68q66obb7mKe410jmgXbUccUL8E5ftGl6WVXX/d/dqN+PWrEcOaB+VEWiyRS/9xcLxXzLa5GscC9tMWNtzOmE6l7pLzJzsuUx3yIkOCPT3HzXfc9zBzJMwzL4qD34pJhK7ihZnnLe2Wk+nGfsHBi8jfjRkfL5z2/QpVtAbdxaxcU04k5nOeKifVyB5WKQaQyhIAQEAJCICICEiw0OISAEBACQiBXCJhJfJ0fv1+5nOQtCOLm+FKly0GAeP15W4zMo8k3xPywN6pb6fgOrW+4Oppf3VLmJ36VOYF3/uaDKutcFwSt2sVXNCshvXEoIG4skGDlBXNnhlwrBW34Foaw8BOq/NCFtJpqPtXjXV1WoWr1WqE2D3z/vSDf5rvttvvuuJgwUWYHKxL8XbOq/urGp594/UXnnBLk8iWo/vjdxo0KpHmuOthzcs2TTzmDeAOxxJJMxhPymf6bPX3yxFTh4i8H3+rEEYBwYLzEM05YVck5QeOD1fqNL778Gu4Tv3AHcYAbFlZDfmyuS7zWFdSrSbOrWvA3SJQ4+/yLLg0dC1sb+NuRzrJZHQ0ZRsDidPTD6h9WhQQLSCFX/s1t2ndEoPTGfXGrqCMJohdcds31CD1+jEqWKRdym1TXBNveYQIyx/wXdvcRzTIskXYjIpjnkBlBq+OJi4OoGYqnYfOtt9xE59vjSm0jvgn06g8onEh9g/IeYK6S2P9LOBB9IuWZ1lSS/F6rsvzoO4hCMMa6otvLzz7hb8PxpcuUDxLYmcc5754br7qoSb0qJ+CSLIiITAQTb17GB9+D3D2x/8IrmodcLUZyrYhgGkk8TGRMJNrOZOZK2lG+So1aCHWzp09J2zzOe0XQOwUkNe3kHvH2QaR3Bn+fcl99+kHvnqeceU6jVMeZoh9bP/Do02O+GD44UiwkVx/zmBeKzfOjuc9z+3g+3tC63YPEFyOGDfNzvG4vY43d3FwvVfNtr7dffYG5MlUxRJKdl8HqEBMuvdizDyuoBo0vuhTLLQJeR7JucQHIP/sk2MWk6wssgbhPpnjc1sXqJ/e++vbLzzweJHI48SjofTVW2TouBISAEBACQiARBCRYJIKW8goBISAEhMAOCPBDMshkvVnzlreuXbP6R/8KVFsIfhCFDBs0oG+Q6wr/BRAWMD2PBr0VeTDH/WQdBELdMxo0xD+/190LRAQro6OV61aA+13WHHnMscUh9H4wESXe4UDMC/LivzroHEguCOd5s6bnECwQMnADxMrAZIiZwR/0fdeRK/HWNVI+6oH7DoLNJlNWJuBJvS0ebijOg2lVU5JpR6xzDjGGGAEBYtCshwaxstn5mo527iHG5qwztzdBVh+nGSFNPIag8VM5bJmBKPLe26+96L0GK7lrmIURsRf8ZCTuoHBnEVrJGeBChnLSWTaudZYsmDcnVWSYH1tnYUFfcAyf3Oc2veSKj/r0fNtLQoI7x41D38FFEcTWaWef1+Rrc2HkF2SdT/+jix13PK6T/Nd3K+1TReowl61asfS7oDF0zU133MP+IGuOROfbMuUrVaWskcM/HRhrrCd63Fm1HHDQNuEika22BYdnJbLXUik/+o5+py9+WLliWZBrP/qdYLV+N4L0A4Ijwlc8AmYi2JDXBYH+fvmyHcbIifVOPxPyc9sYyWn5wT4ssELWChHcsyUyJhJpZ7JzJXXGJQ1//c/MRHGLlp/3CguRkUMAJH/ji69oHrpHfEJvpGdc0DV4NvMcci6FUlFv3Ow9/XqP939evfrHh+66qbn3WQIRXqNOvdO81znwkEMPg5D2WpBgnWHvRvu++9YrzxPkOkhAT7auublequbbUZ8NGcS9iViUbDu85yU7L1OGTYOHrVuz+idveXd1ePxZLJKxesFCNhL+ZcpXrop4G+Qi0luei/nDop9420u8NTD6bNCH/YLOKWUTQrrvvXjrqnxCQAgIASFQsBGQYFGw+1etEwJCQAikHYEjjjq22BpjPL0XYuUrLo4gQvyCxX7GaJDXFldvjFU5F6QRYjNaXlsUGAo++Pfff+UIQH3xldfdhFsWb4Bd8rFilL/RyiWYIqvV/dYfbkXk2gR8sFew1aCQpJFEhxMsQAX1IXC5t53/w2pjTKyC8HHurNzqxFh4RztevXbdU8HSH4A83jIzAc9Q359QOtT3LohvvPWPNx8uQchLQO++3bu8zD1wZctb74x1PmMY//b+fAhZrHjF+mJg355d/cexVGDfJAt473c7dVqD85qwunLksE8/8gshdU6p34DVtNHiaqSzbAhSc909NxYuyR7HIgu3bUeYwohFVbuOz75s+K7vZgFKvWVunzsCsG/Zul0HSEV8zvvr4VxyfDLgvR5BFkfmBa48pE+kODOJtsv0wn2Mr89BblHGWY0uuMQFkZ87Y9pkf7mJzLecW6ZC5ZBg4Y93kmh9g/IjuCBQYZWSSHkEqIaw9AdFz+u+I07EUWbqQd1ZqR3UBgSLoNg49EO6xDnqsdfe++7LXxfrw9UN66w2Dz7xPN8R7YOeeQjqzBPTfe7EXBmJjIlE2pnsXEm9mD8QYv3CUCLjKlpe5gzmR1w3efPhYqfxJVc0N6Fkir+fIz3jgq4D0YyFmZtHcltv6vuEuY1ExLv3tmsv81tHQYS/+u4HQ52wtW3M7L2PNW+9uzai+HW3tbm/q1kOMVaI/5Oq+Su310vVfAvmc2dMnZwq3JOdl4PwwOqjdr3Tz3rh8fb3lLCFFeQJwp84Pgjx8czRib6vspCH9/evv/p8WKT5CvEL67AlC+enxJ1dbse+zhcCQkAICIGCi4AEi4Lbt2qZEBACQiBPEOBH7+ZNmzd5L9b24adenDDuqy/wq+9W5EO8ksd+H//JX0c2RavkoeZ2gePLly5eGC2fIy28K9m59tU3tWqzbPHC+VhYeM8/zFwdxCoXsjaInIcY4Nw9jbzy18nc1pfGjY53P1YSJ9hqUNxHRIqZwA9Azlm8YN5s77kb/vozjNWeIUEm2sZ1KlTZ5nrKbUWNhOKzLaLM0T+xygo6jqUK+4MCkMZTXibgST2PPHpbTAOsGVy9IeSwIImnHbHyuFW2+LdnleQH73V746Y77w25d/Cfywp+RyisM3OkA8Muc7z5EN04FzdGQcR4dQvKTv7hgz7o6y+fODHss6CcH/iP1TVyhH3jzU95pDals2wIF28fQJQ4VxOxMI73uFlBLYN0I44LpP6rT3ds73fxsm7t2tWU58eee7LZ1dffQkwRf1Bk5gBnQdG/Z9fXg+pjQYrLf7dwfsoEmX+NPYIw914LMaztI091dpYL39kE4q9LIvMt5+JqhHGbSqLS1QnR7Suz3MBtzXkXXnpVPP1IGx/o9GIXiONeturbe05e9x0kOcQ+Y+irzwZ/7K8/9zIpqN/pB9MkY87j8WASlMdZENoQyTFGrrz+1jshZ0MBos0nfVDMporVatVmblluMSyCyk5kTCTSzmTnSuqIlaTNmdvncO5JJ9wli6H3PJ7ViJ57hBdDuGNYM/FuYe6WcoxFjkd6xnGMMe/egfi+k33hb7QYWom0o+Ud7ToQ5+jVZx5tH/Te8rm5DuL9yBvoG0GGceGuc9/jz72Ku7beXV/v7OJNpHIeSPZ6uZlvmafpLy+WvBeZZ8BcvxNRZrLzMuduw+OfEP4IYfc9/vyrxKQgzoZzZbjmxx9yLAbaNkdve5fA8jbWGClaxL2v5pwXQuPVhErq4C3D4l3UAO9vx3w1IlLZvM+ykMc7dmLVQ8eFgBAQAkJACCSDgASLZFDTOUJACAgBIbAdAYgO3CS5HS1btW0PyWSczipcX8yeNmlCI/O///W8H/5glawL8Ohf4cYPtHYdn3nJBRemPPsNtx9/CXwZDXLiKnDclQmp9PBzr3VjJVrnTg+287vgiFUulgQVq9Y80W8dwjVWLlu6hL/VwkSxqxff+w0fN63JpdtiBriNeAms0p4cxYcwefjxt3b1jz94z4XggxzzY8WP2xa33X3ftbfc2c7lv+iqFje9+8nIb1mNzD4EjOssD0SfBcnOlZ9vfvA3vODSK8E5VvDooH7KFDypGyuO+bvnXvvsw1+I0z5Dx0zBgiQVtzUBLiGhZk6ZEHKd1fmJB9uZ54YVr/X6cFjJ0uUqeK/x1Ovv9Ov4fJd32IfrIFa4lqtUtYbLw/2CP/JF5hKtpwkW/vohspCflZD+GAuQDpUt0C9u0oJ801cxC6JQQNXZMwOD2aezbO7PnYw12tOsBmgTYsXb/YeMfOiZV95ORR+4MiBVSpQsXfbO9o89g5uN/u/uKC7Mn73NDRtxINx51KfTK117b9y4CtUyNAAAEW1JREFU8Z8n7r/zZn+dEEEQaiEGgyx1uN9xxcEK8FS1h+DMrL7lvnbj+PGX3noXtzouUPtPHl/07rqJzLecw1wzb9a0tLhLo/znOj5wN66dHnn+9e6XNr/xNoZCJIwQf1/r9dEw4vs81/G+u/x45nXfIUJR10/69+4R5NvdiVg8+/xtYu5kTLj+4zhtZ/7hWZXbceKCd59y5jaRkg1y+vZ7H3riG4tnxJiM5PqtWq069bD+iySoJzImEmlnsnOlG/9u/uB7h6deerNr/6GjuHdzi6U7n7bQ526RAgQvz13c6FnsgBzucqI94xA/e378xXiEa1c25XDOpPFjY5LOsdpTq+5p9W+++/5Hvhkz8vOeb7z0bFB+rM3Y/4+9ELjj/3isRy679sbb6597/oXPP/pAG54LuCMiXxBhHqs+kY4ne73czLfdPhw+5vm3e3/k+rCmuUhEiJ/0TWyyP552JjsvU7azqAy9rz77WrcDTDV/6cmH7+PYvvv9Xwj/IMEIwYBjWPnEqqNzKVXtxJNCCxvc1vzm1m15XzTj3pBFndvc+0ek91Xen7BQTuY9MFZddVwICAEhIASEgB+B0I92bUJACAgBISAEkkUAVzSnn92o6XW3t7kfQuaMcxpfcMW59apff0fb9vyYa26kOiIGq2P5jnhAINrmtlIRgo3Vwac2aHh+wwuaXQlBT+BgVxeLTbmOzxdd2eJGhJHa9c44q9k119/S7ubmzbz+w1kNBjF7wx1tO+yy8867nHJWw8Z1zOc5ZQW5vHHlXnNT63umTvh6DNeGsDy3dvlirFQ1L1clWM3Mj/Y+Q8dOeeOFJx4miCV1YVU4Aa3xPc2KxDEjhn1atlLV6lx7va3IhMzK+QOwWoiAnhcQUNvlg5h2q6T9/TDMVs6zShaCY8GcmdOJI8Gqe8SYjm1vb+nyY0XS5sFOz+PDmpV35WylHCLQs4/ce2e0gOXx9PsV19/S2hEYnbu//8mKZUsW/fj9iuUGxQ/0yyZjdlk9Csm9h/2HIIS/avIM+3hAn0zCc/l3i0Li1j0PP/kCVg2Xt7ipFdgRpyAeLGLlYfUj49v1J4LRzZeff+bbA4aOem/wVxPf7/n2a1ipsLoYn+Iu7sSn5tP81rYdHnvqtXf6skoW4q31/R2f+nvD+vV3t7zigiD3DLgag0AYNXTIIEdIufodY0GKEbaGfDRkUFBwXwJ+rjJ/95FW+KazbOYAc6m95PRzGjW1WBMrzjqv6SWQIDdd2rh+LHwTOU4sAUg4LLAeaHX9lUGxAxAlce1yiwXk5t43zfB7yL8S5tOpjQVIdoS/97qIIHzv/+7bgdYVEOwQxP6YOonU3Z938Ad93r33sedeeblH/8FmMTOAeByIbNxf82ZOm4JPdrvkrv7z7FZdEO98CzHIvDLdxJ3c1DXauQiwzZueedILXfsMZP6EKMXV0wyLjbPGlD1WPhN75aTTzjznkmta3sK881bnpx79qE+PHcSsvO47+p176cPe77wV1EYnWAT1+3CL2XROk4svR5QbOvD93sXMGu+Sq66/Gdcv3mdesrjzDOTZhOsf8w613+67774HzzdECETTdwaO+DpofHA9cxlYwXS7SU+83PU9+ufFxzu0dfVIdEwk0s5k50rqhpjA+L+t3YOPY/nCewftzO2zzov/sI/792nz0JMvPPTsq12ZK6+99c52WJN2aH3jNX5xJ9ozjvceiOPrb7/ngeNNtD7iqGOOhRgmTsxEexYk2+ech2D55Cvd+kB61zrplDPeGzxqosVO+mTS+NEj1/704w9777vffggtt7R5oCOCn91mY9317Dm+GJH8ubfe+xD8Ph3Qp+foEUM/4bizzuSdJjf1856b7PVyM9/SnvMvufLaN/t9+iWWpieefGp9e+Qse++tYJduibY12XmZ6zAmEKGpG+8CD999Swu3aAX8Q1Y+YYtkb72wRCTuiFuoE63OY0cOH8J8xOIWM9j9g2ddg8YXNmt62TXXT/l23GisObznMy55Xvpdobo8xSzKOKJrkPvKRLFTfiEgBISAEBACQkAICAEhIASEQFoRwDXDoDHTFk5b+cfWUTOX/ez8UmNtMGXZr5vZh29ebyWwRhi/4Kf1nEMaZ9YXkHF+d0qc0/GFLu+4fPx9s+8nXzjy3FsmBN7kpb9sIs/UFb9vgRhyq+n9ALA6uv+Ib2a6cictXfcv1h0uHxYiE5as/Yfjr703cLj/ehCSn02a/723Xu8O+vIbF+DQe717H332ZeoDsRDUEaz8+2rG0rUDR02ZH3QcVzWfjpux2F0LTF/s1vdjggj782PJ4nDt//n4GWee1/TiVHR+e3PJ8s3C1X9NWf7bf942x/p890OdQm4zMglPiOQeRt65cfLUa937+l3tJIsZ45dyIQ39ZXAMkpax4HBjLCMquLwXX339zfSvO87qUBc0OqhON5gbEPKXrViluv84K0kpByIq6NzB42d91+mVbr0jtTWdZXNNgpG7e2zElIU/eC2rksXffx7jH7yJ8xCtTAi9UbOWr3O4D/1mzjLwi3QOIkj3jz4bG2l+IcgxZV14xbU3pKotkERc09WRdmGlgJsXSCb2Q8wFXS/e+ZZ5mjkUkjpV9Y5UDgInpBkEa9A8QvsY/9H6gbLzsu/aPvJ0ZyyeIrUJ8py2BD0HmOc7d+83yNtW2s59kCqsudcnfvfzRu84Rrin/Jd7DBjMuA66FiutOefj0VMX+N2yJTom4m1nbudKe+047otpi3+i3t8uWr3h+lb3PJAqHF05PBd6Dxk9yeE5fOK8le79xn+tWM843A6CP2UNmzB3xY133veQ10VUsnW/w0TtcfNW/Y7YzTx394P/3979hVhVxHEAJ6UnV3fVqKjA0iwpekio6J/5EhtpYilooQSSSBAGBVHqQ5ahhZHSQ24SopaFRFQWFgUm+SLCShr5YA8RUhAWGokWKO1XuHA43b1/9np3bffzsCDu3JnffM7cOWdn5sy8sv7r3qO/lr9Teb4ob0uYZ5JKv5e3EIpbambCO3ms79n+n+0EBxrrQMtrpb/Ns9s7H+7em7p8+8OxEy+/0bO1vEXUQOuTz7XSL+eel34uz1VZ8FOM4+FHH38iMWdCtxxf2mTeKGo07vP32h9/O128d6zZ8Pa2PAeX88hzcfqB/vLOW6LJZ+XaDZsaLV86AgQIECBAgAABAgQIDJlAtjbIoGllYD9/YGYSIAMhWS1bLbDO8RMmZhXt9Nvvurfe+QE5GyL7U/c36F/JP4O7GWC5ZtJ1U+phZOA6g/4Z8Kq2jUS2cShv4VPMMzHnUONZ8xYurjZ5UEmb+mcFaK148iZErbrFNyvwMvhU7ZyDYt5JG9t69W/m95XtFM7/gd6353H+4L+i73yRTNxkECSDOBlYzLXM4GkGk8rX9GLyTD3iWJwsaMajv7RxyiB5rQGRtIecB5L2XHSt5BnXtOFGznNImmwHUi2eDIZlBXK1MpL+/N7eNdpJO/OuxJu2lIHLWtsCtXpdqg3KVMszbSFvTaUNp29opdyY5+DSfBdbyaf82Til3WRVbrlfzcHulfNQBtrfZvK5PLl8IePvL6+0w7TjvIGQt93y76z8brTsi+XapT3nXlUr7twnY5wB4Ubr10y6uCX/lFPcfirf56ysrpZX7j2Z1Kr2PRxom6hXzwvRV6aPS32L9WzGqpG0mZTMvTc/5f3+y5+vd49LnXNuUSPlNpombT+TJcX0ccl5GvkuZSFHtt7q7z6QQ7grbwaVy8yij/mLlixrNJZG0rWjvEb62/SN/U0wNxJ3rTSt9MvpB3LPL+cfp41bdu6qdi5LrmvehGsm7nzHu+fMX9j90LwFtRZBpC3Ue87OM1+9Z/ZmYpOWAAECBAgQIECAAAECbRfIAF1WoVZWcvU3QNL2QBRAgAABAgQIECBAgAABAgQIECBAgAABAgQIjEyBrNravmvP/mxvlO2VMmnRyJsOI1NLrQkQIECAAAECBAgQIECAAAECBMoCo5AQIECAAIFWBbIFxfu79/X27Z5w6WOzZvQd2nfyZA5jPtZ3sG6refs8AQIECBAgQIAAAQIECBAgQIAAAQIECBAgQKCuQA6PzMGBazZu3l45tDF7727a8clXdT8sAQECBAgQIECAAAECBAgQIECAAAECBAgQIECgVYHKeRVPPrtidSWvHID4zaGfji9//sW1rebv8wQIECBAgAABAgQIECBAgAABAgQIECBAgACBmgLzFy1ZlnMqnl7x0qvFhJOnTrsp/3/f/Q/OQUiAAAECBAgQIECAAAECBAgQIECAAAECBAgQaJvAmI6OsfuO/PLne5/vPTBq9OjRxYIWL33qmUxYdE2YeFnbApAxAQIECBAgQIAAAQIECBAgQIDAsBNw6Pawu6QqRIAAgfYLzOyePTeTFtt63nz93NmzZ4slznxg9twjh7/rPfHH78fbH4kSCBAgQIAAAQIECBAgQIAAAQIEhouACYvhciXVgwABAoMoMGny9TekuKNHvj9ULPbaKVNvvPW2O+/Z8+VnHw9iOIoiQIAAAQIECBAgQIAAAQIECBAYBgImLIbBRVQFAgQIDLbA6VOn/kqZ47q6xhfLXv7C6nV54+LTne9uGeyYlEeAAAECBAgQIECAAAECBAgQIECAAAECBAiMMIGp026+pffnk+dee2vrznGdXeMvv/Kqq1eu3bApZ1esWrexZ4RxqC4BAgQIECBAgAABAgQIECBAgAABAgQIECAwVAJLlz+3KhMUxZ8Pvth3cEzH2HFDFZNyCRAgQIAAAQIECBAgQIAAAQIE/r8Cl/x/Qxc5AQIECAy1wPQ77p7RPeeRBR1jOzsPHzyw/6MdWzf/8/eZM0Mdl/IJECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAgQIECBAgAABAk0L/AuIgWkCPYjfhgAAAABJRU5ErkJggg=="},{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"U3RyZXV1bmc=","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOydd3gc1bn/PzOzva9678WWu+SOjQuY0ME2JXQSQrjchHQIuQkp5Ia0m5DGj4QUQkmA0GJMDdjY4N67bFm9r1arXW2vM78/1hZ2sEEGBxs8n+eZR/aUM2eONN855z3v+x5Bo9HsVBSlGhUVFZXjIAhCsyBJUjiVShlPdWVUVFROXyRJioinuhIqKiofD1SxUFFRGRWqWKioqIwKVSxUVFRGhSoWKioqo0IVCxUVlVGhioWKisqoUMVCRUVlVKhioaKiMipUsVBRURkVqlioqKiMClUsVFRURoUqFioqKqNCFQsVFZVRoYqFiorKqFDFQkVFZVSoYqGiojIqVLFQUVEZFapYqKiojApVLFRUVEaF5lRXQOXEMJktaLVaFBRikQixWOxUV0nlDEEVi9MYncHM9LkLmXHW2YwZPxG73UYiHiMUDCJqNFgsVkRRoLN5P2tXvsZrL/6TcEQVD5X/DOpSAKchFmc2N9z2VRacM58ta1awfvWb7N29A9+QF1lRjjpXo9VTNXYC51y8lPnz53LfnbexfefeU1RzlU8qkiRFkCQpDCjqdnps42csVJ56fb3y6euuU/Q6zQldW1w9UXl6xQYlJ9N2yp9D3T5ZmyRJYUkUxW8riqJF5ZRTVjeV//3pfdx1y1WsXbOOVEo+oev9Qy70GcVU5FnwxrT89tGn0af87N3b+B+qscqZgiiKSdVmcRrxhW/9L/d/5w46unpP6DpBlLDZ7QhAMhEnMyOL2+68luV/+xNX33grr/3rzXddE49FCYfDJ6nmKmcCqlicLmjt1BZbWb951wlfmlNczd3f+wGCkP6/qNExadJErNokueV1fP+XD77rmoPb1/DAb377YWutciah2ixOj03QOZTlq9cpwkkoK7NsvPLQww8roFWWrVp3yp9N3T7+myRJYdUp6zRBifvY3TzI5Zdd+KHLyskpwOXqxZiRT2jIdRJqp6ICqoHzNGLrhrf573t+zoS6Kvq6O/F6vR+onNJxkynNMOIKKhRlm1j5xsqTXFOVMw3VwHma4Rvo5vYrz+ecS6/iju/+grzcLDrbDtLV1sqAqw+PexCP24VvyI17YICA33/McnRaiWRCZlLDdHZs2gCARm/mS9/6Ho//9kcMeIY/ysdS+YSgisVpRioZ51/PPc6/nnscnd5ISWU1JWUV5OYXUFU3gekZC8jMycWZkYnZbKa7rYmXn/0bb/zr9ZEykkkZSRKZffbZ/OQLvwbgwmtvY/rsOXTtnsvTz754jDsLVI+byGBvO17vO2JitlgJBQPHrqwgYjIZCYdCxzxsMDu4ePFiXnr6cSKxxHs+t95gwmI143G737uBVE4dqoHz47uJkkapntCg/PLR5crnP//Zkf21085V/vSP5cofH31sZN+Vn79TeW3LQeXldTuVF97epkwYW3VUWbd9+5fKg4/+Q/nHa6sVm0mnAIolq0h55vW3FI2AYsuvVO79yX1HXbPo6tuUb37rmwqgXHzTl5RFC2cfdfw7v31C+duLbykXX3SugiAqX/z+r5SX1u1U6ifVHXXe0s99TXl2xQbloX+8ojzwpz+dFCOvup3cTTVwfsyRU0kO7t7KD+7+KudeumRkf29HC3X1M3nusT+N7Hv6oZ+zdVcj3//CNTz7wqtUVleMHNNbc7jgnGl88aar6PbGyMuyA3De4mtZ/cLfSSqQm1+MxWg+4u4CV1xzPc/9/REAyitqEJBGjhaNnUZNjoYXX3wdvdHABdfcTpE1ya9/8wAzZ541ct7sC6/l3LMmcf2Fc7n9usv5yQ9/iHLo2IJPXXQSW0vlw6KKxSeAzOw8/EOekf8HBjo42NzKzh07RvbVTl1AsS3Ftl2NFBQU0dfTM3JsyU3/RXCgj/GzzydLE6al242kM3H1DTexdcNaALJy8wmEfSPX1EydT1mmRHNHf/p43tHHF197M8v/8RjWLAeCaOHmm67mJ9+/B6PBQiASBA7ZUe76Fn/61Y+IxBJccuMdnL/obADGTDuH666/+j/QWiofFFUsTkdEDZdfezOZGY73PbWgfAzf+eGPePjBIx2sZF547jmu/+ytAOjNDr75vR/yqx9+m2RKwWw2Ew1FACgfP53LLlyAtWwSd9xxK9/64q2kZLjpy98lP9OGkpIBgXMvvJTi4sp0eSYbd93zA5LxtB3CkpnPjBnTKDl0vG7aQqaNK2bZshfJzMzl4ms/y/N/vh9fIIJGq0dRUgB89us/oDgvg3AwgEZv4tIlVyInU4gaPV/79nd58P9+fJIaVOVkoEadno4IIld89kssvepqPH3t7Ny6mY62VgbdAyiKgtFso6i0nCkz51KQ6+TBn3yPDRs3H1WERm/mF399huHuAxTXTmH183/mrw8/CsAF136BSxfNZO2GbVx6xZXc++WbKZmyiCWXLOSlZcsYN20euRaZp5e9wa233kxXvxd5uAtb6RTcrTupGD+Nlx/9NbXzrsSYGKK4diKvPfcEV1z/GdasepOG6dP49u3X09bZy08eXs64UhtXnLeAWFKmpmEe9957D83t/Zjw88rKTdzyuZuIpyQUJcmKv/+BRGYt1dlw7/fuPQWNr3IsJEmKqGJxGiMIIqXVYxk/aQol5ZVYLBYEARKxKN3tLezeton9jY0o/xa2fhhJq6d+xlkEBnvYv//AkSUz57xLKczLZNWrL+AaGASgruEsJk+eRH9nM6tXvE5KVqiqm4zdomfb5o3ojTYaZs6ip3U/7e0dSFo9DbPm4OpooqOji8KyGsrLS9ixaS3BQz2X4soxCIkgnZ3dI3evmdCAzaRl26aNyIpCTkExcjzCuVfcSm15IXUTx/C5pRcRCKu5OU4X1BB1dTuttmtv/46yZk+rMqGu+pTXRd2O3tTZEJXTBlGjZ+a8eTz+u5+we9/BU10dlWOgioXKacEVt36d8bXleD2e9z9Z5ZSgioXKKceSWchVSy/iiccfRxTUP8nTFfU3o3LKufyGz/PKE3/AH4oiIJzq6qgcB1UsVE4tgoaLLr6IZc88g0bSkZDfO4ZE5dShioXKKaV4TAOBrt0MDocx2GyEj/ACVTm9UMVC5ZQydlI9u7ZtAiA3Nw93n5qs53RFFQuVU0p2XjYDPV2AQHVNJS3Nrae6SirHQRULlVOKb8hHbmExk8++mLirEU8geqqrpHIcVHdvlVOK2ZHDfb/7EyYpyX3fvIO2zp73v0jlI0eNDVFRURkVkiRF1GGIiorKqFDFQkVFZVSoYqGiojIqVLFQUVEZFapYqKiojApVLFRUVEaFKhYqKiqjQlQURRUMFRWV90RRFElUFEVNIKCiovKeKIqipiVSOTZ2hxNBUL8jKu+gioXKu9AbjGTn5lM/46z3P1nljOGMEwuL1YbJbAEgr6DohK7Nys075v78opIPVJfcgsL3PedEvu6SJJGRlfOB6nKY7Nw8YtEIkXCI7o62kToKokhOXsFx2+xE23I0GAxGMrPf+3nU3s9HxxknFgXFpSQScRzODERJev8LjiAjM+td+yw2GwbDB4vDe78XzOZwMnXWXEwWy6jKKywpR06lPlBdDnNYbEorq3G7+rDZnen9mdkIgkBmdu5xrsv+UPc9FiUVlQT9/uMenzBlGmWV1Sf9virH5owTC51eTyqVoqC4FFdvOhxaFEU4IlGsVqtFEAR0ev3IPrPFSiQUBqCwuDR9nk5HXn4R/b3dCIJA1Zi6d91Po9UyedpMcguKkCQJ6ZBAWW12IuHwUeem63EYgZLySrZtXEskFEKj0SKKYvr6I76mh7+sgiiSnZvHsG9o5Jj+kIhptTqycnIxGE0j50uShCiK75R5CEWWcWZmoSgKFquNUDCAVqslJ6+AQbcLQUjfU9JoQBAQBAG7M4Nhn5eS8koKikvRHGq/w/XTaLUI/3afI59XFEU0Wm26zCPbTqMlHo8DUFkzlqLS8pHfk95gQFFk+nq6yMjKRqNJ31NvMKLXGyitqBpp/3Q9j/5TFwRhpE1FSUJvMCJpNJRWVB/VJlqtbuQaSaM5o8VJ8/6nfLIoLqvA7nDi9QySSiWZNvtsnBmZtDTtR28wEPAPM2HKVLo62ggG/LQdTC/7l1tQSE9HOwAWm50x4yehyDI2h5PSiioad++gtKKK9uYmkskkeQVFiJJEZc0YPO4BsrJzKCotA0UhFotRUVXLyleXj9SrpLyKsxacy/rVK3C7+qmbOAVnZha9XR2UlFei0eqwO5x0tjYjyylsjgyikTAZmdn093WTkZVDbl7ByFKGFquNqbPm0tZ8gLLKGvp7u7HaHeQXFuP1DGKx2QkF/NTUTWD96hW4+g7lkRAEcvMLGRp0U1pRRTQSoWLuQrweNyaTGZ93iIn10w+JhBO9wUhHazMtTY1U1dZRWzeBpsa9ZGRl4+rtxmy1otXqSKVSpJLJkRR6WTl5nHPBpbz47BPMW3QhNruDQbeLN17650ib5OQVUF5Vw2vLnyOvsBhFUdDp9djsDgRBQFEUSsur6O/roWHWHIa9QxQUl9DX3UUqlWLshMlYrDZ0ej0OZwYvPffUSNmTGmYcEieFRDxBflEx+3ZtJysnB2dmJjqdnmGfl+ycPPoPPUc4FMJssUDLmbkI0hnXs+jv6cbv86EoChU1Y0glk0QiEXR6PTV1E8jNL2Tvzu20Nu2HI9YQNRpNxGJRBEFAlmV0ej0H9u3G4cygr6eLZDLJ3h3bSCaTAPi8Q0xqmE44FEIQReLxOEajma0b1iJJEt6hQYKBdBdb0mjIzS9AkRVMZgvjJzfQ3dlOZ1sLgiDgHfIQi4RJxGN0d7ajN5jIzs0nOzcv/WXNzKa1qRGPe2CkvsGAn0G3i9KKag7s240sp8gvLKa7ow2jyYTFasXV10vrwf3vCAWHeg2SdKhnZaCorIKmxt3IskxOXgEe9wCFJWW0NDViNFno7epAkiRMJjNmqxVZUcjKyaW3uwONVot/2IcgCGTl5NLUuHvkPmWVVSPDQFlO0d56kMGBfo6oCDq9nq6ONmrHTSSZiBMOBbBYrBSXVRAKBNi5ZSMIAgVFJcSiUZoP7MPd34ecSnGwcQ8FxaUc3L8XhzOTzrZ30vVlZufi8w4hSRJ2Zyb79+6it7sTg8HIzi2bsFhtbF73FnkFRTQ17sFoMlNcVoEgCOzauunk/kF+jDjjxMJqszHkcWOzO8nIzCYQGGZwoJ/c/EJaDuw79AIrFJWWkzpi/F9QXErN2PGUVlSTSiawO5xk5+bT3tpMIpFAFEWcR9g0otEIPu8QeoOB5v17kSSJ/t4uIP3VNxrNI+daLDasNjvbN68fGWIEA37kVAqNRkt1bXp4095yEEEQyMjKorOtGVdvD6lUkr6eLsZPnop/2HdUfRVZwT/sQzz04ns9gyQSCXq7OgkFg1hsNvbv2XlU+zicGXS2tZCZlUPjnh34fUOgpKdSRUnC4czAP+xDbzSye/smYrEoGo2W0opqFFmhtWk/A309pJJJAsM+yqtqUBSFoH94pNcjCAK5+UXs27WNnPwCdmzegKuvh2gkMlIPo9HE3h1bicdiOJwZeAYH8Pt85BYUcbBxL6IkoSgKGo0GjUZLUUkZFVW1CIKIVqcjOy8f/7APjUbDgX27iIRDI2VrdTqqx9SRSMQJBQNkZGah0+mRNBI5efn0dnWiKAoB/zCCIJCdl09z415EUSQ3//2N0p9YBEGIcRosvKpuR28l5ZVKRla2kpNXoJx70eWKIAinvE4numVm5yrnXbLkP1L3KdNnjfy7qrZOmXn2wlFfm52bryz6mLbpqdoEQYifcT2L053C4lLKq2opKatkaNBNWWU1viHPyFf540RFdS1DgwMnre4ajYbacROZPG0WgwPpJQMEIW0I9gyMfgmB8qoaPIPuj2WbnkoEQRBiiqLo3v9UlY8CQRCw2h0EhtN2Fa1Wh6zIpA7ZQj5OaDRaAJLJk7fKmNFkRpFlotF3hiwGo4loJPweVx2NVqtFVpSPZZueKgRBSKhi8THn/MuuYPLUmTz7979ysHHPqa6OyicUVSxOQyzWtLFTFEWCgQDBoP+YX0BBELh46TV4hzxsfPtNrrnldpKJBK+98MxRsyIAoiRRUVXLpKkzyMkvGNmv0+rYvnkD61a/QTKhrjGqcnxUsTiNEASRhedfjMliYXDAhdFoIievAKPJhMFkIpVMEotG0zMGQtqpa/Pat9i5deNIGbn5hZx3yWLszkw0Gg3RaAQBgXg8htczyIa3VuLq6xmZ5dHp9Mw8ewFzzzmfZU89xp4dWz/0c4iSBjmVRDjkcKXI8ocuU+XUo4rFe2C327Hb7Xi9XgKBwH/8fuOnTMXV243b1X/M44IootPpMVsshEOh9x2jC6KY9glJpRABUYDkcex5kiRRVlVDe3PTUdPFHwStTk8iHhupgyoWnwwEQUiosyHHITMzk/nz53PZZZdhMBhGdY1GoyEvL4+JEydSWVmJTjd6DRYF8bhCAekvdCwaYWjQPSpjniLLI3EiGhEWFoD2OL/tVCpFy4HGDy0UwIhQHK7DJ5nK2roR35qS8iryCt8/mK6yZux/ulr/Mc44d+/REgwGyczMxOFwMG7cOLZufe8uut1uZ/r06cyePRuz2cymTZtIJpN0dHS87720Wi19PV0nodYC6Wnxo4nLEEjAtGxYpy5SftLIzMpGr9fj9QzSMPMs3l7x6vteox/lh+d0RBWL4zA0NITX6yU3N5eqqiq2b9+OfIwvpSAIVFdXM2/ePCZOnIhOp6O/vx9ZlvH5fMco+d0kEol3XJ3tOYizLkHZvxGlfQ9Gi4aSsXa0ssyw10D/hKUkVj8NvqPfeqFiMpJWS/LAZgAKamxMXlSIaLbwRvBqdgz0cF3jbxgkhd0BdjOs2QPR+AdrH50G5k+C+ZPTQxz3MPxzLbT0jr4MQRDQ6gwkk/H3jJYVBDgVLhFVY+rIyS1AUWRSskx3eyt9vd0jPSZZTqHRaikqLae3q4NoJEJ2bh5ejwedXo8syzicGfi8Q5hMZsLhIKIoYrM7jvK2/bigisVxSCaTvPLKK4RCIWKxGAaDgfAxokRramqYPXs2Go2GUChENBqlra2NLVu24H+P8Op/R1EU0OrR3Py/SJKA/rJbObfn+0ybm6AoQyaSsPKLge9QKSkI02cw67GbeK5VxhcHoXwi2rseAUFCuOciyouC3PSzaax/tp1O+6coOXsuhMOIbpn1eb+m35cWiWQKbrsfdrSMvl00EkyrhTuvghljYfVOONgDY4ph1S/g6dXw4yfS4vF+OLNyGT9tPt3tB2lr3HaUk9SYYrjuHKivBr0ONuyDP70C7ccfqZ00DEYT88+7EFdfL5vXv0UiHkcQRex2BwVFJQSGfYTDIeKxGIlEgryCIgZcfZjMFsZMmITXM4jDmYnf50Wr0xGJhCkoKaWrrYWxEyZjNJnZvO6t//yDnGQkQRDuAU4sscPHFEEQyMzMxGazkUgk3neMHg6HSSaThEIhAoEAsVjsqOMmk4nx48djtVqxWq1s3bqV5cuXs2HDBoaGho5T6vERZ11GQf14vhm4g2mzBNZn34rjb/+PFY/s52XlM2SIw9xd+FNetd/Kkr6X+cEYH0G9g/3/9SSpV/8MQ304xpRz0+cFVv+thTef6Mb/qe/ydeNPqS/bzSPJb/D2z57i7ofCPPQSyDI88CXY1Tq6l9BqhPtvh7uvSfcibrsfHn8D3twJy9fDU6tgai1870Z4ezcMvodgiJLE3POvYua5S3Fm53Fw92YS8SgAU6pgxf9BOAYvrIPXtsDECvjZ52HzfugcOH65H4aMzGwsdjsLz7+Y1a+/Qkdr8zs9HkUhGo0QGPYRj8coLC7F4x7AZLbg6u3BarOTlZMO7HM4M2g7eACNVksiHicnr4D9u3dgtdvxeYdAURjoP4Eu2GmAIAjyGSUWkiRRWVnJ4sWLsdvtBINBgsHge17j8/nw+/2EQqF3uQeLoohGo8Hv97N792527NjB0NDQBzMU6gyYb7ibL0u/w9yQw2DnAK/5LmTd4y/T6jEQvPx7dP7oq/Ss2IFz0iReHHLw2subKF9yMyarlcTjP8AfiVP1hc9h3PMiq/+0jyuuqUVuuIjp6+5h68EEydqZNDUJRFv2kUwm2dYMe9rhL99I/2ztO1yZd3JRHKY4Gx69G0pz4YofwLL16Zf5SAIReGMbpGR48CvwyiYYOs5EkiCKVNY1kJVXzPCQm33b1pBMxMm2w1P3wEMvwtd/D9sOQnMvvLwJtjTBrRem7xE/Sc6XRU4T08qzcQcilFbXkZGZzZqVrx8VeHYsLFYbblcfgwMuQsEAGq2OcDCIwWhiaNBNwO8jHouSX1iMq6+HorJyopEI7S1N6A0G/D7vyXmAj4gzTiwURcFoNNLQ0EB1dTWTJ0+mo6PjPW0LiqKQSCSOGUeQSqUYGhqit7cXt9s9Ep4+GjQaDVarlVQqhSzLSNVTKK8poFpeT2tUzyPf3UasbCYEhhCcuQgZeaRefohuN/SHrFTdsATdrn/ySv33adj1KL8v2Yu32MjuqltRnvgtD94SIDbtCpa9FWf5b1/hwDYfZy3MoajqGsZlO+hubyYaCdHWl34hH/pa+mXsdr87VV2GFf56FwTCcP1PoMv93s+2vRkiMfjF7bBuH7iO8V4oioJnoAefZ4A9m1fjdfdi1KWvGQ7Bt/8CiX/T3A4XvLQRknK6V3QyuGVuDaIgEEvJJHVW9AYDxWWVxKJRwqHjf0gC/qO7TcGAn4Dfx9DgQLr3EYsRCYfo6erAP+xjoK935JqPm1DAGSgWAH6/n1gsRlFREUajEZPJhMvlOm4PQxDS4+fL5khcPj+LBRMTNFTLGHXQNwSJpHJCAUl6vZ7KykqWLFnC7bffjtfrpbe3l2RmEWPKgsh6P8/8fDeh4QRCfgWCyYo4ZgZK226U/elcCqngMJFFX2XpQh8bk+ew+9f34C+2s/BLY/D785g/SSRyYBf3Ju4hvOIZ5O4myowyn8n1Uzn/CmpKqxno76OtaS8AHQPQ3AN/+BpsPQjdR3Tz85zw52+kbRy3/kpHXHRgMFqJxyPvaXXcecgO8rPPp20axzJ8RsNB+jqbCfgGybLD7+5I20Nu+9XxbR6pkyQUFr0Gi0GLNxRDFAWaXX76envp6Wqnq6ONUPA/71vzcUIQBPmMM3DKsszGjRvp7Oxkzpw5JBIJioqK8Pv9RxkwrUb41FSYWQcTxo+jcPLtZBbPJBH109W8gWs0UVytb/HSq2/xxjaZpu7j31MQBOx2O/n5+SxevJglS5YwefJkBEEgHA6zf/8BorkWlKEWnvvDHmLh9CdVbtmB5qq7EK1Oyvv3YJ27iP27txBwdxHcuIZ/nPMV6sTNFNyYz4RrKzE17+Pnzv9haexxjAMppJpsJrvWcM4kuKEaXtnShDh9A/mZkxA5uhf0ymZQfgeP3Q1v7YJl68BsgK9dAV0DcOv9GgqqZzPlrPMIhfysf+0ZXN3Nx33mlAz/7wXY254Wm5Xb4f+ehoPdR0/uaiSFuRPgp5+D7kE4585j90RONtFEijH5DsYVOLAatAyFYjQPBPCGYijHmH5WOcOjTjUaDQUFBQiCwMDAAJFIBAE4eyLctiSLqrEzUWyzyB97JSlFi0ajISsr65DhMwGpCEnfVva9+V1efGMff34VgpGj72GxWJgwYQIzZ85kwYIFzJ8/H7PZjCAIDA4O8sMf/pCHH/4rqaoJ6Dq3Mjx0hCFAlNBc912MBiM3FhjIyS9jy9qV/OuZPxKzZaO7+i4+Pf5Vzq4dYkakCW/jAPc/A68nF5G65vvc1Px7but7jD1D8NhBWNkDY+fWU1A8li2vvY5n8N2WwhwH3LgIFs8BvTZttPz1c4Bk5OxLbmT2oqVEQn5efer37N74xqjauTAL7roazp8Gbf3QP5TuqUgiVBak7SEPvQS/W5YevnxUmHQSi+oKCcSSrDrQf8ypcZU0qrv3IQ7ncxQFuGIeXH9RCUWzfoIxcyL5+elEu319fWi1WrKzswkGg9hsNoaHhxkaGsKiT9D81rfYtuFVfvqkwuChGVNJkqivr6ehoYEFCxag0Wior6+nv7+f559/nhUrVrB//35CoRDHc6iCdLzF+YuvpeHsC9i9fRsrnn+YgG9w5LjVlPZ78AXTX3SdTk9SURCScUQBEke8A1llVhLZYxjevPk920Q8ZLaQlXfaqHbKXGafdyWpZIIXH78fT/97O5IJoogjMxcU8A72ketMz3SU5IDDkh7iNXbApv3Q/xEO4yWNDostm3ljiuhKZlGcZWMwpOBy9zPs6WbY20siPvqQ9zMBVSz+jRsWwY2X1WAZ8z9Y86aiKAplZWVIkkRPTw+xWIxwOExrayuLFi3CaDQSDAaJxWIE/UP0bv4ujVuXcc9fwRtIv2B1dXWUlpZSVVVFOBwmEomwc+dO2traCIfDo7J36LWQlWFk5vQxKIkgbS1t9HmSBMJpXwlZgcShUYXRbGHy9LPBns2ON54nEjza1yOzyIRcOgXvxs2QPDGPLK3OQEH5GCJBPwM9bRxP3A5jsWVwxefvxmA08+yff4q7t/OE7neykTQ6svMrqf9UNUZLJgF3GYImndVbRCYaDuPrayXoG6CnfRsB30fg1PExQRCExBln4Dwe8ybC/3z5MuTCL1E5fiGZmZlotVq0Wi0tLS3o9XoKCwtJpVJYLBaSySQOhwOdTofBYEBvMOEsXoAU3ku+qZU1u9Mv8dDQEB6Ph+3bt7N161Z27dqFy+Ui8T4h4YKQ9rIszk7/dHmS7NnvorN7iJQsIwImAzitaQNsdWFaONDaueCqz1M3dS7heIyepqNzXNhzDIh5pYQ6eyF1YmHpcirJsKefUGB03QBRkpg67xKyCioIDg/R2Ty6fBs6g5GxU2bjyMwh4POclJgVo9nJ2KmXUjNtLuPO9eEsdjHs1pCM2Ukm44iSFhDgqzcAACAASURBVFkYJKPEg8Fkw6AtYtjbQzIR/dD3/iRwRs6GHAunBe77YiWOcXfS6UoyYcIE9Ho9RqMRWZbxer04nU4sFgupVIrMzEwMBgM6nQ5JkgiFQnR0dFBUXIqjaD6aoWdxuQO09KanCCORCLFYjFQqNaqeRI4jPStgM6V9H1y+9HQhpHsQgXDap8EfTvdgej1pB6gsO+TYFRxZBWRk5dA+HKFz+zqO7AHkVzkx1cxDcA8Q9fuOUR+BI9dQ+TAkkwki4TA6g5HWxm0M9o2uZ1FSMYYln/kqVeOnEva76ev5cD0SkyWTCbOuwJlfjqxo6W3S0NskopFqQNYgIKAz95NV3osiG6g9u4dIUIZYEd7BLhT5w4vVxx1VLA5x3Tlw4eJbsRafz7Rp04nFYuh0unQafq+XvLw8YrEYQ0NDBAIBLBYLkiTR3d2N1WpFp9NhsVjSixNJBtxuL+Wmdby6+d2+Au+H05Ie03e74UDX6K6XFYgl0tONvYNJmvbtRfJupC2cxOsagvg7Vte6GeOZOfkSasprcHW1HB2jkJGPeNZihOKxKOFhCB8xhNGbEPLKIJWExNFGWKFoTLorFPu3cb5Wj0cy0Lp5JQOdB98dhSodnow7WrD0eh01dZOx2Gy0H9hFb2crHxRBEBk34xIKxlaRW9uMLPeTihUjkAOyZqTnkIhCwBNHUVrIKFKw5UUIDSlIShG+wc531fFMQxUL0tODd9+YQeHUb1NUNo7Ozk7WrVvHmDFjgEP5GmWZYDCITqcjmUxiMpkwGo3EYjH0ev2IgTQej2MymUiIWfjbnmbQG6X5SP8CSfO+UVHxpED/kIA/DHYd1Dmh2Jz+qdMIBAwZpGKHE7IfQqMDexYk4qDIWHN01C2wUTHNiZiTT7irl1g4iaQVyRtbTKZtLBaTlYGedlyHv9qCiDh+DhpPC0Lnbhg7B/pa0MhJTDoR49zLMUgCSsk4Uq7OkSGMUFSLNP4stKXVKHozysA7Rk+hdhrYMkmYnchDvWmhOYR2TAM5l16Ko6GeRE87ydA7ghYOBulpP8DBPVs4sGf7h8riZXXkMWtxCaUN7Vizh7FlWzDZIOB2IooSklaHzqgQib1Mdrkboz1G0GMh7JNIKR5S4WwiwTDRyOjjfD6JqGJBuldx8UUXYi67GqPRhM/no6SkBJPJNLLgTnNzMyUlJSQSCcxmMx6PB4Ds7GwkSSIej9PW1obZbEYURXQGC/5AiDLjev615R3jI4r83uGTJhvSDfcizbqUy0vauPtLWcy7vpJr5uq5sFhg7yUPEr70a2hyihF3vUlcJj29+tmfoLnm24jV9UzJ2cuN99UjKAodG7ux1Jaz5LY8mrd6EIuqCSfgwKpVeAddtHd1EPWn7Q9S+VjmXFnGkitk5i/NIyfPxIzMQv634CDnzp3ExHFl/ErzEtNr8yirKGW20opOI8KCC1n86RTnz/cizrgY74EuYi43GMyYZ1+KtXUbUU8/VDeAuxMUGSmviFnfvJLrLulhzASRoosWUlUSpG27m2RcBnsWgbwaBtubSIbecY7SizArB4bjEBvlLGdJxVTqzkmhMYbwu0z07JqOnDKQiBrTSxoqCuFQF4l4lJC7nv7WBGZrJcmoGYvTRDzmJua34/OcjBQCH1/OSLH4d1fmr10BtVOvRuucDoDH48FisWAymUbWuzycMctms40MOYxGI+KhbFRarZaMjAz0ej1arRaXy8WgL8G0nFU8/q8ogcjR99fpdBiNRnQ6HVqt9pCbuIB0xZ3k51q4rGY/rbNvxbV7FetX9rENJ+vnf4G4qKX4qS9ycO63+JHxLdY2eYiXTkKz5Csk7r0c84XXMX2enrd/9QaNLzRj0xbRsldDT3M30766mIFhMwMr3sY/6Kavs4WoIkJWIZIzi7O+cj5XT+xn0aatTGjqJJEt0NZwIa++3MyTpnnsWPYcf9sdZHtTD91FM6n07WPWpdPh8oXc1PQczX/bjdftJu/mT+Ne9TaJjEpmTJ/HnPoZhAd78EhGMFrAP0jhp6/mgvNjbPzLel788UYOtpopbChh0WIr21Z6YPwC8PYjVk5BGehETCUY54QH5sA5RfBMG8RGMTzTaA0UV03AXuQjIz+L7u0ziEcNxMMaFOXQlLmcRBAT5FUnMFgUjMYKRO0+HIVdDA+6CQ1HIFaCu//gqYmTP004Yzw4TSYTxcXF5Obm4nQ6cbvdtLS0MDAwgM2sYLRX4w0E0Gg02Gw2srOzEUWRSCRCIpHAZDIxMDCAyWTCbDaPGAVTqRSiKBIKhUgmk9jtdgB0Oh3xlA6TowyjfgeQFpyCggLKy8sZO3YstbW12Gw2enp6eO6559jVP4w4bT5ftt2DG4lnWpaw6bfdabuB1oc9dwp3THqcz3wpiNT9Oq21F/K3hU1cbz6L0K5VTJiQYuyYjSx7eyLmzb/gwvnFlMy5jfGY+ee2XZjaYtSY99EefMe6LwY9NGTEmX9ZBQXj29A/uJL7d4ZZ2QPe1DaW/q6C9oVX4VqzB7k33ZvCH0fY1kjbrFsYN2Mi3b/+C02bm/lcLVzt28AfA/OJLJnEusYSov3taMdMpKxmIgdeeBzhrKVorFZmXJxP20v/ZO2T3cyYvwRFo2PVyzL2Sx1M+9KlrH9sF0rHHgQUCsdP4EfWDczNh+XtcO+2dM9iNBiMNowOiPkn0HcgRjwaxejwEwvJyMlckEUEjYvisfvJr4mTSsi4WhvZ+UoBOeVxkqFxxPwpRCmEgHCGWy3OkHwWZrOZ+vp6Zs6cSTKZxO/343Q6Wbt2LZLoI5UIMRgYxGAwUFRUhCzLuN1uotEoubm5DA8PE4lEUBSFZDKJRqNBlmU0Gs2I4fNwYBikhSEjMwshlnb00mq1nH322cyZM4eamhqys7NxOp3k5uaOCE1Pc4SJhtV09nr56/2txG7uRMjIRwn7wZFLJKHniW/+i4z7JnGWYSP/o1xNrg8uuGACb+7YwSVfGccL/+9JDBc/zCu/srDbVU6nKZsciwOp4+/seXsd//2H2Wx4Sk/EE6M+Gz43BuaPifPG0lwe+9kWNr4cJiXpEJ25GCI+Wl/awuIrB/n1/W8e1Z4G914uu2QsGx7/Awdf3gXAFjfkGxXO0m8lf+liFsrNbHjqESJtUxkeGkCOBNGIAlNunkelsJUHHtiHKFgoqZmAxeak5/VlLF+Rx6euz8XywDJmFsIt1ftwTb6cvrW7uOSVMPt9cCI+lslkjIhfxFHQRTKWi0anJzIMGq2VVAoEEZDtKAQJeGSsWQZyK3WU1g+y+41CBAxkFRbjat6huoBzhuSzEASBvLy8Q+tiamhpaWFwcJCuri4un53AkVdHRum5hEIhMjIy0gsf63RkZmamoyM9HnJzc7Farfj9frRaLaIoIssy4XCYaDSK0+lEr9fT2NhIXl4eQf8QFt8jPPRCAG8gbd+orKwkEomMDD2Gh4fZu3cvq1avpkOGXP9qnn9oP0FfHKFiEmj1KO17EOvPRcgoYPAfjxKVJQzTqumyfIronqdZP/kb3DB7J9YDjeS7GrFNm8umtd388S9NmHNKcfV2sO21Zwh4QjhyjMw8O5uvSy5urIFV/QIrpoylL6iw/IH96QCt/EqK513GVVfdgCFpJ7cuQOuOAQKe9AyIpBVZ+s0JCCEvbzyw/aieeTAJjQf7KJxbw+fDK7je2EdrezvbO9wIksC5F8DCRTJP37OG/uYAiXiMVCKKLMu0bF2N+cAaLrpQ4ItZPq5zhFnTk+KXTWaWexwM9PWf8OuaTMTJyKpESc0kFrJSOXsd/e0HiAeL0GiNKIqMIOjxdDhIxHQkky4cuXqcBQrtO1I4s6eQiIUZ7m/D3dt00v4eP46cMcOQUCjEypUrWbduHeKhFc0jkQipVApvAILu3Zir32mKjo4O9u7dywUXXEA0Gh3pRRwuS1EUMjMzcblcOBwOnE4nJpMJRVGwWCwIgkAi0MKwt59o/J3gta6urpHZFUVRkGWZWCyGx+vFfvUtbHy9nZAv3ceWNyxHc9WdyGufQ6yYRGr9MgDefrKV8vocsup8RG7/MxaDhvL4Hm6070FzpcIfG5fxP8XfYULBHawsm0P9ugdYnB+kzglzBltovnQOXfud3PGijynX11ExfyHL7n4JOaUAAmJhNfqufeQsOpeCnFz2bWpl0a21PHLXJrR6iUu+PI7isQ7+9OUNh645GiUaZvjV53ljYQHu5wTuqldYeraNNfVjKG/I5snvreHgBjeiADpRxtf4NjW+DdxXE+ecQljT2sOK4hKuf8CNLw4Y9yHOuBiGPTB4okZGBXdfE9kldcQTQ2j1Ccomy/j6duHtKkWrLU2v1m7IJjRox2jvZ6g3RCopYLHNShs/vQP4vX2c6VOncIb0LCCdJi8ajRKJRIjH4yN2B1GAuvxe4rYLKKuoRqPRYDabMZlMI56DeXl5aLXppfiGhobQarWYzWZ6e3vJyclBr9eP3MfhcOD3+9n2yp3sbuxg2bpDLtmyPBJL4vV68fl8DA8PEwwGEQQFQ3UdQxs2o6QOdbR9AwglY9Fc8Q3EkrEk//FTiIVRZNi7uo+G0jb8+kw+5f0980PreGyNzFd/B7H9TUQzimm/+v8o613PVzt+Q6FJQVbg4Z1JNrREKfjcZGoXFmKZWM8zT8BgIg8l6E3Hflvs+HavJzzswaN38OZjz9JwQTZ1C0spXHwxZaVJ/vatDbg7Q+lp4OwShMLq9FTqIT+LiD/B/Bur6DcY2ZyVS+Y148gOhznvja0sjHi4thJuHQtfmwg31MB4e4qdHvjOFnhybYBp11bT2hLD55EhGkLx9CHWTgONFoYHORGSiRiZOeWY7KUk4t3UzbNSNlHA6/IQGy4llUwgShokTZK82n40+hj+ARlfTxZKSiIw0E1X6+Yz3pNTEAT5jI8N0WvTmaLMlbew4Mpfkkql0Gg0+Hw+vF4vZWVl6HQ6EokEw8PDOJ3OkWGKLMu4XC5SqRTFxcUoikI4HGbdWy8T3X4jv31eZvWu0dVDWzuFRNPO9PTqYSQtQvmE9Ivc3zayWxTFQ06WCsgKWk3aKesdBLA4IOxHkFPvfBNFCRSZ/CoreRVWWsI1+JtawTeIMG522kbS14Kyd226lOxiMFrRDx2kdvEshg0V9DcPE139AsgphIpJCJmFKN5+xLxyaFxHytOHqBE473O1zFxajm9I4bWHDtC8uh2nRqHaDvkmGEho8FTOoV+bzXBbE8mWnSO1H3vpFKidyYFdMRR3F8r2FelnNdkhEoAT9Kgsr51L8dhZ5FQHmXxRO/7BBDuWj0MjlRCPhdJrq0gStpwgBeM3EPU7cLdL9O3JoLt5C70dO07ofp9E1NgQ0lGaGgnG53eQWXMd4cg7jlZ6vR6TyYTb7Uav14/YLA7HhoiiOOLtaTAY6O/vZ/v27Xj2PUjA08pDL6XLHw2yp593dXUVGYb6IJj2shRsWWSX1jB9wUUYS2rwyyKJkJ/U4RxzJhtCfiVCRj54+4+O/cguQZx5MUJuOYHWbvr3DRDPqAR3F4SHoa8NpbcF+tvSYoSAEg4gFI8h6fMx4DXh27KdVDictqdEQoiVk9EdWE9Nlp14537iY85CGexGicVo3uFn3d5CdrQV0B/JQbZkEertoCsE+4ZFOotn4Y5CeO8mKJ8EWl06Y7nehLf6ctwrVqHseBMhpxhBp4dhd9rN8gNMX4ZDQ1gt2egsfrJKI6x5zI7RNA5BENFodYiiBkEUSUQM2HIGad3owNct0tG4hf5udf1YOEP9LI5FuwvmjYtQUDqO4ZgTh8NBX18fJpMJi8VCNBolkUhgMBhwuVwYDAYikbTzhMFgwGq1MjAwkE6x1/wWZt8jPPiCTPtJXqNDVzaOhkVXMmfaHHJtFloatxPOqUwLg6IgTDgbJAkUEMfPTXtM+gfBbEecdiHK5lcocTqoWfRpQgEfcUcuSn8bHEqUm45CTWf+EgQhLVYBD+L4uQhmG0r7HvC5EDQ6xAnzkPe8xYTqKm7+769TVl7JzrdfR66sR/G6EKqmIIfDxDe/gdK1H7FkLOhNMOxGKB2HkFOKsu11iIVQ+loQx84CSYM4fi5KfxvKgU3p+3t6EcrGI+gMacH4AKSScUJ+N1qliPZtoNPXIEoaUskYsdAwoqQBBYb72unZE2eoe4imXWvwuttP0m/u488ZY+B8P0LRdFancdNfI7d+GslkEkmSRgTBbDYzODhIRkYGpaWlxONpI6TRaATSWcBDoRAhXyeGgd+wZleSdftOfj1TFifulj14c7JIpWQiri6UZCdCdQOKqx3BaEHe9i8AlK5GxEkLwWhBsGejNG1GDHmZOrGeqrFjyMr7Ais2riX+7/Ech1AOD4ciQeQtr6btE4fctZWu/Shd+wHwZdiIJ5Lk5BdjS0UYCAcQp56H0r4HpevAyLBK3voaQu0MxLlXgiCm63l4OJFKIG9+BWH83PSw48A767eSiKHsXYt0/i3IgoDSsfcDtV3QP8C+ba/iyCjC6vBjNDsQJW1aZEWJRDxCcNiFd7CDcMirBo8dgzPeZnEkF8028cv/+wnGnDkkBDuyLJORkYFWqx2ZFbFarbS2tmIymSgoSK9I7vF4aG5cz9DWu9i7v437/g6RD7h4z3shNHwKoX0P+TYbipKityPtVSiUTUAoqERu2wV9RwRdSRqEgmrQGVBa0/aQmQsvZsaCS2g5uIfX33iJWO8HD9KCdLaxaWctwGZ3sObNVwkFgqAzHBW8dhQmW7onc4K5NLBmIM66HPntp9N2i5PBIW9eAeEdcVQ5Jmd88htBEHA4HEQiEaLRdFf8gtl2/veeL+Isnodr2EB2bgEOhwODwcDg4CBWqxVJkkZmRwbdLja98VtS3Y+wu2mIXz2X7qlA2jkrNzcXo9FIKpVCEASCwSBDQ0MjszInVN/6RSiNG979sogacGSDb+B9jX+SpCErr4BIKIjfd+JrmxyvTFESSZzg84yqbDE9SaMAZOQj5JQgNG1CltWpzI+SM1osDjtqFRQUEAqFOHjw4MhU6cRKiW/cMo0pUyYR047BUXgWtoxSzBYLQ0NDmM1mgv4huls2ET74Cwa7tvLCenj6rSOCxoCSkhIWLFhAdXU1tbW1VFRUjGTX6uvr44knnmDNmjX09PQcmsoVEGdegjR3KdKqv1HV8wYNkw3UFCuYhSRbDOcSWLWSgx0xOgNpJ6hjIWlFSsY7ya+yEg0mad3mQQlGmDsBqgrTSXM3H4CBf1sBoXSCk4YLixFEaNropvGtfqyiwvgMmJAB2UZw6kFrAgogvxySJgOrPLmsXB3iwKbBE7I/WjP16E0avH1hUkcs8Z7jgHPr0zk7M2xw5x+gsRPsWjin2kaTK8QejzpM+Cg5o8XC6XRSWlo6kmG7ubn5qIxMWgmmj4GzxkPDGCPZJTPJKJiCPasSBJEh1wG2rv0nL69uZ+1ecB9j6RGr1Up9fT2LFi2irq6Ompoa8vLycDgcI72KV199ldtuuw23241YPhHLN//KdW0/ZeXUb3CZ7VEyNfuJJ8BmlUjGcrg+/iwZ7SH6N8BzTfBsG6zrh8PvWn61jcu+Pp7ccistWwfJytJSXOegtPcApYNt7GqF4hyRqgKFVTsVvvfX9DogJeOd3PSzaWx7pZt4OMmciwrR7ndxxa59xFNpd+6+GCyYAZPngGSEQdHO64564oMJtBk6Xn/Tx5M/2E4y8f6KMWNxKZd8eRxDvWGScZlHv7mJgDvKNQvhnuvSCX+efBNe3wptfXB2HnxrChwchq+th6iqFR8pZ6xYlJSUUFtbO2J/aG5ufs+VyfIzRaZUKuQ6FSQpnalqTzvs63j/mbzDEamZmZlUVlZSX1/PggULKC4uJjMzk3/+85/87Gc/o6NpH/abv8eiqXEWVq7i+dZxvMktRO9cgByTyasuouTCehbNcuNcs475pQn+8QRclJNeIf3H26E7P5PrfjyVjc93sP6ZNuZUxvj+TdAWsbCteCprn25j4wv9TJ4xj4IcE2cXrOKiKT6+/oiOyd+Yx5qnWmld1sp/j1FY2mDkxaVzePu3u3lpeT86fXqhoclV8MeXIJgQGfvfZ7HsSRcb/9bM9Q0CU77ZwJ4DKZbft50Wz/FtABMW5rP07kk8+f1ttGwd5JzP1DBhYT65G9bzqbFRvvEHWLkj3UsrNsP3p8K5hXD/bvjDPoioQvGRc0aKhc1mY+7cueTl5ZFMJlmzZg2tra3HTXd3eMnDZDJJe3v7h04XL0nSiHG0sLAQnU7Htm3bGBwcJPt/HuCa6uVsf62Rtc91I9yznNTff0i238Xsi66n1R9gfN3bDLsCjHc3cvlZsOQ7MD8b/uuSDLYuncm/Hmlm9eMHuftqhRvOhZ//Ax79F5jyLPzXg7NZ9tMO5iz4OkaTiTf/+RdsoTe5874qdnqc+H+1mc9VKzT64N6tEBqTy5X3TOHhr6zjy/P8NFTD9T+GrkE479ZaxszO5aEvrkNOaLFn5ZHv8LH4u3XMl9y88KsmHtoAoX8bKjnzjdz621mse7qNNU+lHc0cVvjOL2rJrMrgZ5/ZQGOHgk0LS8vhrsnQ6Nfww116dvaFkc/gMPFTyRnnlCUIArW1teTk5FBYWMjGjRtpamp6z4SwBoOBhoYGKioq6O7uHjGEQvrFP+zJOVoOZ9TyeDy0tbXR2tqazsKVmUnO+ecztGIZ655uRU7ICFmF6PLKKBMSzLrkZgoy81j15HLOu72U3/ysi2JnipsvgIeb7ZhumYZuVTNLulqYv0jh3Glw80/h+TXpdUFDvjjhQIJzPlND1y4jBoMZuXcXeYIbadFErtPuojQZ5Ysvw893QlcI3J0hBtv93PHLKUzX97L02yn6vTB+Xh7n3lLLP+7dzlBPlIazL2LqvEtwDURZ+cwW8q4Yz40LYtycEeBAJ3Qcssdq9SJX3TMFd2eQV39/AJT0MgaP3AWFspcdxiqaGsPUy/+/vXuPbeu6Dzj+PbyX5OX7/RBFiXrbcqw4fsV1nLrJ2i5L1i4BNhgI5mIFhgDJP/mjWIY9uqFYu6HrMGzpgKLJijULkG4B1m51k9VJ2mRpkzpxHn7GsmxLtqwnRVIUSfH92h+UKMt2LNp14i06H+D+Yd7Lc48I8ud7zz3n98vy/Xvh023wlUOCl42fJrTtPoqFPAuJj6gqsnRNQoia7lZ34uMkhCCVShGNRnnppZcYHh5eM8u2Xq/H7/ejaVpzMdkyu93O0NAQe/bsIRgMXpFYpxXLgUbbsInCyPu8++OxlRnf2QVqriDT5RoxnUYxPU86VmbkVzH27u/jL56BhMHBHz+1g9FXRjn401E2fKHOF3vg378Hx86szAlVBEy8NoFFl2fIcICHp/6Bb/W+zxefGOLcOzG+/Kcp3DvB0b1SZ8Rlgy9tnGNT7jz/Zd5FeHeYh/9qGw9+ZYgffvMY4yeS6A1GQl0DBMM9hHs2kJwt8OxXj/ATbQjtAT///VX467vBbxHc+wf9+LttvPTd04h6nft2wBv/2Bgz2feXNU48fZLH/mwTT/6GwnNn4e4fwyvTAleon8jG7Qxu34uiyKlBt8q6uw1Zzk5VLBZbKmTsdDp59NFHyWQyHDx4kNHR0eY+i8XCzp07ueeee4hGoxw+fJgjR47c0K2K+d7foTR6isrFlZKAoncr+if+FQpZtP95Dt0bPySbTmJyCB777l1Ez2eIbHZReO8cv+sew6TWeeZlOPgq/M0O6LQ2Bj/nCtBvh4AJzrV5Kf3+NiYPnEO3q4PUQpnv/9FhitkK2/rgX55oJAqemYff3N54YvLot8E8GKZri5t0vMA7ByZIxRrzKIROIdI/xNCdezlz7C1GjjfqsQ7s8vGlr29liylOWy7NiYyXgtPMC994l8JCmi/fB3uH4LmfwNuH4cEO2BWEFz+7g6MnM/zbP400P4fOgdvZdvf9TI2d4t3XX5RzIm6BdTlmcb2cTif79+8nGAzy/PPPc+LEiVX7XS4X+/btY/v27VSrVZ5++mmOHDly3ecRnZuoTwxfMWKq27sPgNqb/7lqrYfda2Tw7gCxi1kuHJvHoDQS7eSWEm8LGkl+H+pqBI25fKOcwLNnwb4rxNC9bYy8NceJ12YoXPIM1mWF++9sPL6ciMHL77IqLSCsVHBbpqh69AYjxXxu1Q/Z4de488FO2vrsBEWGxyJjeNUyRgFiAqY/gHIakkX4jzH4wTlIm4384ZO7+d7jh0jHl/8Ygclso1TMU63cePJe6cbJYNECn8/HI488gqIovPDCC1cNBIFAgP3797Nnzx6EEDz++ONMTKzvBK+XE4DJCG4zdJjABJhUOJaAWH51Al6r20i5WKV4+eiodMsIIcrrasziRmiaRqFQuOYtSzQa5cCBA/T397N7924eeOCBZrLfteh0OoKhMIZLcmJ8EtVpXPVMJuHQNLw6DS9ehMnslZm6F+eLawYKf1sIj8//0XVYuoIcLWpBOp2mVCoxPT39ocdcuHCBp556ir1795JMJlEUpaWye7VajdnpSXr6N6KoKhfOnaFcvv5p08u3BlcbZK3X6+h0OlRVT3tnhI6uHsKRbuwOF5qpkcW8VCygU5SlICdIxKJMjJ/n6DuHmI+3vtpTCIGqqpgsVqqVCtVqlXK5RLWF8aFWdfX284Xfe5jv/N03blqb0trkbcgaFEWhu7sbt9vN8ePHVz06vZzBYCAcDlMsFpmamrruc5nMFgaH7qAt3EE6tUA+m2U+EUNVVcwWG1DH4XLjdHlwuj0YDAZsdgeFpdWxy+n6hBDUalWE0CF0glq1Rr1eo1qtkojNMToyTHxulkQ8RrVSXlpn0RiDEEKgUxRsNgddff1s2b4Lm8PJ6ZPHeP3lF694eqRTFLbu3M32T+3BanNQLhXJ53OUikWKhTxGzYTBaMRktlAqFijk80xcGGPkg+NEZ6evq4CQEII993yevZ/7G31KLgAAB/5JREFULf7+639OsfAhi9Wkm06OWbRICLH0A/z4RuGNRg2Hy43b68OoaZRLJWq1GnMz02QXM5TLpY+vP0IwMHgb9z+0j8Nvvs6h138OgMPl5vE/+RqH3/wFb7x6kOw1ZsE2mhE43V46u3voiPTg9vqwO5xUKhUWM2mmJ8eJRWfJ57LUajWMRg1fsA1/IITb68Pt9TF2Zpgf/eCZlp5kSTePDBbSdRFC8LnffohITx/PPvVtnvja3/LPT36LudkPvz1rhaIoON1ewp1deHx+bA4npWKBarXK3Mw08ViUeHSWYrHQUmFp6eYTQpQRQiwXzpSb3FraNt2+tf7N7zxT37LjU7e8L3L7eDYhREleWUg3RFFUqlV5K7BeyEen0g2TgWL9kcFiDZGePgA6u3tX/XuZXm+go6v3mm20d3Rd9fXeDYNXfd25NLD5cejuG7jm/s137GDj5i031HZXb/9VX4/09KEuZRpr9T03y1pzWvo23vaRnv//Mxks1mCx2tBMJjTNhBACu9O16ssWCLWTXUxfuw2bFWgEluW8j0ajhqK7+sQtbyBIJp36tfptMltaOs5qd1xzv95g4OzwjaXDd7o8GAxX/jBtDudVH5maTGYMRg3gqu+7GfzBEKVi8UP3a5r2kZz3k0AGi8toJhMujxezxYrVZkdRFDq7e1nMpLHa7CzMJ/D4AiiqijcQxGZ3NL/4vkAQvcFAqCPSbE9R1eZyD/dSdfZAqJ1AqJ10agGDUeOuz3y2mdMTwOX2YtRMzTYBrDY7Hq8ft9ePoqjY7A5cbi8ut5eBwc2EI93N95vMFgY2bcZgMOL1N/pqtlhXnUMIQWd3H/lcFq8/gE6nw+XxopnMqz6P5YlVRk3D7nBiMBix2uxLn5V5qV0DLo+XSxon3NlFoZDHF2xDM5lxeXxYbXYsVitmiwVNM7F56w78wbbm2wKhMPlcFlWvx+FyN6/moDHTtS3cgdPtadaavZSqNl4zGI1Y7Q6EEHR09aw6xulyY7JYUPV6hBCNpzAuN5rJTCAUxqg1cqUuByxpNTmD81JCsPG2LdSpozcYyC4uUi6X8fgCdHT1Mj0xzuiZYbp6BwiG2hkfO0dbewfhSDcnj77HwOBm0qkkM5Mr60I6u3qZungBAIfTjdcXIBGPEWzvQCcENoeTfC5H9ZJqRIqq0tu/kWKxgMPlRqdT2LnnMyiKQnRmitmpSTq7e3F7fUyMj1EqFJgYX8nS3d2/gWI+z+DtWzEajWTSKWx2B5l0iuETjepaW3bswu31M/LBMTbfsYOZyYuEI9384mc/BcDucFKv15kYH6Ortx+3148QoNcbCYTa+eXPD7Lzrr2kkvNLdWMrJBON0oJbtt2JzeHk1PEjeP0Btu7czVu/fI2BO7azkIhjNlsJR7rR6XSkFpLNfgfbw5jMFoTQkc9lCYTauXi+scq3Vq+jqno8vgD+YIhgKNzsq8fnR6dTGNi0GergcLl47+03sTtczbZ9gSBOtxer1Ubfhk243B6mJsbp33gb58+dAQFOpwun28Om27dy9J1DN/Ob9YkgrywuEWxrJ5lMNP73tNpJzEWJRWfJpBaIR2cROh21apVqtUKlUmE+HqNarRCdnqKtPczY2dMcffftVeMNmslELtuYrKTTCRRFZXZqArPZQiw6y8J8gnhsjtpSVm5VVenbsInj7x9GpyiUCgWC7WHGzgwzOnKKQi5HpKePudlpTrx/mEIuR6VSIZ9bqf9Rr9XQG42US41l+L5AkJmpCdKphUuOacz0dHl8jJ09jcVm543XXmnO0OzqGyCTTjV+tG3tJOJzVCpV3D4fo2eGCXVEOH3yGLlslkAwxMgHK3Uaa7UqJpMZTdOYnrzI3Ow01WoFIQTJ+QRWu51zI6eWZnmuzIgt5HMkYlFMZjPxuVny2ZW/Sa/X43J7ic/NYnc4V10leXx+vP4AyUQcm8PBxfOjzM1M03jq19DW3kGpWODC2FlMZjMujxe3x8evXv8ZFpuNsTOn8fgDnDp+hMVf8xbwk2pdZcpai6rXs33XHqIzU9RqNTKZFCazmVqt2qgbUq1isdrIZRfxBdrILS6SSiWpViqkkkk0kwm7w0U2u9gcc+juG8Bqs2Ewao3LZIMRqLMwnwAByfk4oY7I0pcbbHYHsblZOiI91KpVFpLzVMoVMukUsegMxUKBYqFAoZAnk04xH4/h8vjI5Rab9+I2u4PJ8fO4PV6is9MsJOcpl0rEY1FqS+tVQh2dlEolZqcmMJktJBPxRp+WFAt5ejYM4gu0cer4EXoHBjl94mhjGnouRz67yNzsNOVyGUVVyKQWmucPhsJAvRlsctkMi5kMLreXer3G1MQ4beFODEYji+l0cy2MxWpbaqOOXm9AVdXmupTuvoHmGheL1crkxQukko1SBnqDEVVVSSYSxOYak7dsdgfVaoWFpWMMRo1ITz9nTp0kGApz/uwImXSKZCKOw+HCZneSTMSpVMqkFpKUSx8+rrEeycLIl4n09NPR1cMbr750q7siSf+nyHkWl3F7vGRSV8npL0mSXHUqSdLa5JWFJEktk8FCkqSWyGAhSVJLdEKI+tqHSZK0ngkhajohhCzCIEnSNa27imSSJN04GSwkSWqJDBaSJLVEBgtJkloig4UkSS2RwUKSpJbIYCFJUktksJAkqSUyWEiS1BIZLCRJaokMFpIktUQGC0mSWiKDhSRJLVGFEOcURelb+1BJktYrIcTo/wLzExJ6O0R/xwAAAABJRU5ErkJggg=="},{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)", "background-pattern":"" , "items": [{"x": -626,"y": 96,"w": 2749,"h": 510,"type":"text","text": "","text-data": "WnVzYW1tZW5mYXNzdW5n","font": "sacramento","color": "rgb(202, 222, 236)","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -656,"y": 602,"w": 2803,"h": 770, "type": "color", "background_color": "linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)", "border-radius": 0 }
,{"x": -611,"y": 599,"w": 2740,"h": 776,"type":"image", "image":"png", "image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydB5heVbX+9/SWPiG9TBrpndB7R0Cqgg28ci1XsWNDERULdq+KvcFV0WvFcpGuAgISQghJCAkJIZCQEALpyfT/+k2+N//DxwRmQtpk3v08+znfd84+u/zOnmRmvWetVZBcTMAETMAETMAETMAETKCTEWhubi6MJRfklt2cOza1hqGgQM1ahxR95V+g77KoHEujNkaty9Xm6O9FN3Qy/Lt1uZnnAX8qvHXkWVD43uRn8fKPIm9/64che2xhmeOcgmmrP0cvP5JbmIAJmIAJmIAJmIAJmEBKxYZgAiZgAiZgAiZgAiZgAp2QAEZsqgyvRTkGu8LYSh9bo9Inv2/3iLohKsbyhjAAM+Z20eLlBJFO+Gx21ZKzRvTGHHf1bbGifZTZs6pwlRjEHqfW5/Z0YN6+vy3OtY+xW5uACZiACZiACZiACWT+QDMMEzABEzABEzABEzABE+h0BHKeFiU5oyteEA35EF5OUGjFw0JdYODF04KKWEGVYVdv+vNGeqfj7gXvuwQy+1kCBZNFlMBbiHOIcQhxVISL7rm9vTn384Ogwc9Siyhoj4t991l7ZiZgAiZgAiZgAiawLxKwh8W++FQ8JxMwARMwARMwARMwgT1CAGNqGGgRKRAQFCaqXSGbXkJwoJ+t0T8iBcZehBGFJ6qN+7aLFntksR7EBFoh0ErIp6yCpp8J/m58gSdF5udlU65bhAr2tLyU5MVk7iZgAiZgAiZgAiZgAibQZgJ+navNqNzQBEzABEzABEzABExgfySQC2EjTwjeEpfhtWW5r9QDImMQRrTAAIzhF2NuXfT9Io+O/ZGx17TvEsjtT/1dyP6kKJwW3xErFMZMPxvZ/C/yxGBPvyik2iv9+dl3yXlmJmACJmACJmACJmACu4OABYvdQdV9moAJmIAJmIAJmIAJdBgCOcECo2xVzuDKW+JbZHx9pQbXvDfYESv4Hbw8KuPgabEr8mbsk7ybb20RZ0YVnJgWMMH43jcO6+I7YYX4DgdCCq3KLWBMHBfFdXuf7KEnmhcCSqM6x8oe4u9hTMAETMAETMAETMAEXkjAgoV3hAmYgAmYgAmYgAmYQKcmkHnDXEmyMaJjUG8xqu9iwaKly6h6c70lhE5HFy1CeCDcFd4iPaMiSkyIOizq6qis8amox0ftH5Uk5Hi0UGqjro36dNTbow6KynM4IOrjUedGRcx4PmpxCBmE13IxARMwARMwARMwARMwARPYTwlYsNhPH6yXZQImYAImYAImYAIm0DYCrSQZRrBoCdkUtXE3CBaaGIZ5heBhnA7jaRECBX9HDI6K+IBYkRUpnozveEogXjwTdUDUWblzA3Nrvj8HYXruuDyOeGFMi7oiap+oiBScY5yseIFogcjxZAgY7co30rYd4VYmYAImYAImYAImYAImYAJ7i4AFi71F3uOagAmYgAmYgAmYgAnsEwRaSTqsRMPM7xV7P+T1n7/mbKLv5hAtOoQBPgSLyljIxKjvjMrfFHzfGBWxB/GCI4JFfSoq3ZIa6/CyQNhABFoXtVsOxPo4EhKK/B4IEYg4Fbm2CBZ4ueBhwbFLVHKMwOg7UR8OwYLvLiZgAiZgAiZgAiZgAiZgAvsJAQsW+8mD9DJMwARMwARMwARMwAR2DYFcTousaIGxfYdCwi7ywNj+e/m+LFqEUNE1WJwY9dSoQ6LiQYEQgUAxMireEYSC2pCqxvZOhZXFqedRFamoqi6V9gu5Ym19Kulamdbe+UxaN3Nzqn2CvCF4SyBYUOlfiZ0RNviOdwVeGo9FRbhA2MADY1nUv0W9NYSLDbvm6bsXEzABEzABEzABEzABEzCBvUnAgsXepO+xTcAETMAETMAETMAE9jkCmZwWzA3hArFih+GadpFgwVj7nGiRS4o9NOZGHR91XI4JPJ6LSggnEpaTg2JgqhrTM/U8vjSV9OmaSnsXp8JIVbHlscZUObYyFVY0pNLqolS/uiltmP1MKigtSOtnlqQ1N65JxVVFqWETHhTktIA33JtSca9NqWlrWWrajPcGYaPIgUGuDEJM9crMZX58nhf1CaqSeu9zm8sTMgETMAETMAETMAETMAETeEkCFiy8QUzABEzABEzABEzABEwgQ6CVEFG62qqXxS4ULBin5ffzve1lEUIFggHixKFRyUcxIipeDIR7qo66JOqcqCdH3ZzKh1em6hPKUtXELqm4Z68QK5rS5kdLQ3AoTiU9GlNJ39LU8OzGECnqUvmw6tTwXH0IEU0hbJSmxvUb09ZFDen5exrienTXUJkKKppS+ZANqWFNSapb9WyqHF4V1ypS4+a6tPbvW1NT8z/S+nsHp4a1eHmsiUrYKLwxFkcl78W9UeeHcNFh8oL4h9AETMAETMAETMAETMAETCDzFpdhmIAJmIAJmIAJmIAJmIAJvJhALkSULrxItNjFggXjIFqQz2KPPY4QKPBWqIlKiCZyT5Bj4oSoeD0Q7onJIFJMjbolKom1ETDGpuozu6eynmWp68EV4UHRIzVsXpi6jOmbmkN4KBsU4aAqg1lxYyroHp4YzY2pua4wFZRFv40R2qkw+m18NjVvWp7q1/VKzbVlaf0DG1JZ/x6pqW5daq6vi34GtwggDRsKUuPzERKqoDDaLk31awrSuntoH9fWzEzNTYSi4vkQNgqPjNuikiODXBiboi4NAQOvEBcTMAETMAETMAETMAETMIF9lMCe+ytoHwXgaZmACZiACZiACZiACZjASxHICxG1JwQLprNHPC1CqCCc0/FRJ0QlTwTiBDk7EDDIEYEIgOcC5/BWwPBPeKjyVNx1URrwtgPDE6IqVY4sTrUrVqaq8YNSUdctkbOiORX3DneJkqJUUo64URMVrw36wo1iYVTGJuE2YyEq4LGxOG1Z3C3CRw1NW59sTIXF1ZEHo1+IFuFVURfeGJuLUlF5QQgWG+Nzt1S7YGOq37QyPX/3prRp9tYQMXg+CCnkvcD7AoGCRN6IGOTXmBv19hAuCCvlYgImYAImYAImYAImYAImsI8RsGCxjz0QT8cETMAETMAETMAETKBzEcgLQaXF73bBIsSKC2IwEma/Leqfo+JRwXdyRWDsr4iK8X9lVESFutz3A0KsWJGGf/6EtPGhpan36X1T16ld09bH7k+VU6pSUbclqajkkGiL+IHHBv3gqYHYQf8IH4gVeGogXtC/wkzRDoGDdjNTU+Oo1PhcWdqytCTVP98jFRZVRxipqlS3PISLLuvSpkUFqWJkUap7oi5tXtaQVl47P21eiAiCMEL/iC4Do5KoG4+LM6P+gO8hWvw6ji4mYAImYAImYAImYAImYAL7EAELFvvQw/BUTMAETMAETMAETMAETGB3EwihYkqMgZfEjKgY9ydFRZioiYpYgHG/R1S8FBAWRkclqTafn0vVpwxOPU/tnXoc1SdCOK1NXSZH26InUmFJvxAU8MQgnBTJs5dGJUk2Xg+IFwgeiBeIFE9FRUigT4QMxqQdbRAwyEWBdwReGbURPapXalj1dKp95uAYZ0xEhQphA00jQkoVVxSkzY9tTRUjKtPau7emDQ8sTKt+9WSqfRKPkbVRaTg4Nx+EDDw51kW9PyoJumfH0cUETMAETMAETMAETMAETGAfIGDBYh94CJ6CCZiACZiACZiACZiACexOAiFSlEX/50bFk4HaOyqiwZFREQ0QDDDwc0R06BeVEEp4KCA60LZrqhj2aBr30wtS5aiKVFAeibC7bk3FJQgQCAuEXUIcYCwEEPJI4E1Bn3hOcA3hY2RuDO5BoEAcIdcEosazUVe3jLWtPaIF4aK4xvnKVL8+vDYaJkU6jPpUu7w2lfUrSgXFXSNRd3Fa9esVqdvk0vDIKEwrrm1Kz9/yRCT35m8e+mI9HAkHdVfUQbnxSNpN/X2IFwgtLiZgAiZgAiZgAiZgAiZgAnuJgAWLvQTew5qACZiACZiACZiACZjAniAQYgWCwClRz4hKmCQEBHJT4MkwIioeEZxHuJDBHsEBbwiM/HgjdEl9zluehl35qlQ+dHCIA4si7BPCBwIAeSEmRkV8QFQgnBTiBcKH+kF0QMDAm4MwUQgQlJYE47nPHPnOvQgdmzP90B4hhLHGtLRvaihJjZHXov7xZam4f59UUBTraGpIzZubYn5lqXZZ5LdYX5CWfWV5ev72utS4SR4eiCN4cCDK4EXCGljrX6LeFKIFXhkuJmACJmACJmACJmACJmACe4GABYu9AN1DmoAJmIAJmIAJmIAJmMDuJhBCBUIEoZDIVYGIgMDw76jHRUWYQARAGOgbtTQSZa9LFaOKU1nfptT9qIZUPrA2NWxYG14V4dcwtmsqG1IZIgV/P/SJSiJrvCC2hWzaduQcwsfSqLTjs9qRA4PP8rRAHEGgoHKekk1ojhcEwgEiBR4ctKEitnAvogNeEYgOIUY0VMTdZalp4/pUUBqeH4XRprYxbX40xI/mgrT2zk3pyW9sTVuXI4asys2Xz/R/R9SDc/3hUUJuiydDuGAMFxMwARMwARMwARMwARMwgT1IwILFHoTtoUzABEzABEzABEzABExgTxAIsQIR4qicIR6jPmIAoZ0w8iMebEilAw5MZX2WpwPOqUgN63qn0gOKIj9EQYgTvVJh2XOpqeSR1OXAfhFyibBMeGQgGDwR9aCoeEsQVgrBA++JyqiEc8JTgZwUCBgcESgQNvi7gzacR4BgPtxLxcOBIgEDoYNz+k6ftEPEkLjBdwkOfKZfvCX6pvqt4dnRVJIaVjel4m7dIyRUQ9o0f12qe7o2koQ/llb8NDwv1iDgLMnNjfUh5hCuinnieYKwc2eIFogbLiZgAiZgAiZgAiZgAiZgAnuIgAWLPQTaw5iACZiACZiACZiACZjAniAQYsUBMc77oyJaUBAoEA/GRp2dintMS9WvqktdJxel2lVVqWJo7xAo1qSeR4cksKYolQzdksoG9E8FBavDU4G+5D2hnBMIDogKhHxCkKBvxINtQsg2cYFz27wftnkxIHAgXBAyij4lQmQ9LJgr3xkHYUV5LCRc5JbTMhZt8LagMh5zwSMD74/NqbmpOjU11qam5vJYR3lq3rIpQkZVpC0LG9L6e59Ny7//UNrwEOIHjB6KSiLyR6ISrgoBg4JY8fUQLZiziwmYgAmYgAmYgAmYgAmYwB4gYMFiD0D2ECZgAiZgAiZgAiZgAiawuwnkEmsfHuMQ3ghBAA8IxIKBUbu3jN//TY+msqHHpLJBG1Lz1uLwsng+VY7snwort0Ti6vg8YmG0OiQqIgFJuBEC6IvwUXg4IEQgWPCd8EkkriZ0EvkmlIOCUFTkvegZFe8L2svLQqGdmA2iA2IDf5Nkc1nwWV4T9Mv4lOzfLmrDeYQKwlIhcsgThHH5zto3pYb6PpHbIoSO2rivsCCtn7k+PXH1nPT8P2OOzbdHmxNyYzDv5bn+8BhBmMHb4l9OyJ0j5IMJmIAJmIAJmIAJmIAJ7EYCFix2I1x3bQImYAImYAImYAImYAJ7gkCIFYRbwuh+clQ+Y+THaI+HA14Io1L/t4xK3SY2pJIBfVJZ5KeoX7M2NT63OnU7cnMqjdBQxd1Oj3aIDRj/ESf4jAiBOCFRgeUgYigpNm0IE4WnBcIFbRElsl4WiCb0xzX6wwtDfSNaSOgQqqxHRdYDQ6IGfZHHQmIH60O0eDAqAgXXR+fmwfrxyKhMjfVbwuMiQk1tjVpfkOrWbEnLvvBseuYP81tCYm3rY1FUwlEhsiC4IFggmtwc9bYQLfjsYgImYAImYAImYAImYAImsJsI8Iu+iwmYgAmYgAmYgAmYgAmYQAclEGIFRn+ECkI+4clAyCW8BDDoj0+l/XqnbgeXRjLtotTj6C6p/vnC1LRlYyrp9VjqfUb3CPs0PNodERUjPaIA4ZuUJJvPCBBK0I3XAQKExAcEAQz8eCZwjb4YF48ODP6EVWI+hFpCOKAtnxE9+Fsk+wKVhAvWw3Vdk4Ah0URiBfNifMZeHJX1cw0Guh+PEObSEAnDn4uVVKbm4n6pYeuWVPvkM6lqSnnqV1qelv+sKTXXEcIKwQPh4tGorJ3vhISaELUoWP8pRAvW52ICJmACJmACJmACJmACJrAbCFiw2A1Q3aUJmIAJmIAJmIAJmIAJtJVAc3Nzi2G+oKAAw/zOlAvjJgzq5G8gsTZiAob6yN9QUpkOOHNLiBabUvfDhqbG2pWpdOCQSLD9XCqpxpD/VFQ8FHpERVBAtCCUEsKCQkqR0wHRgb8dGIP2iAp4SeBVgbiBJwKeDRjz6eOZ3FwQLbgPAYH7WCvJsRE2JFBo3dnviBAID0qyLU+MOLU9XBR9yhNkTK5f+paXBYm1ERuYY01UvECeDIGmJJVUdkvdjxmWKgasS/WHDUgFlc3pqW8/nJobGJO8FsxZScP5zDhcw3vll0xiV5bcHmj1+ce+2JVDuS8TMAETMAETMAETMAET2KcJWLDYpx+PJ2cCJmACJmACJmACJrC/E3gFQkWKN/5PCT4ToyI+YJBXOKNp8fmBCPW0OZX165uK+5anihHdUt3qFali1NpUWITxHWHhnNwR7wi8FegHg311VAzohEDCI4IiQUEhnxAMMODLuI/ggZEfkQCxgJBUCBhU7qXditw1+uB+JePmM/cSLoo5MC798Zm2rEtz4KjwUIxP36xlfFRyapBzAjFFHh2IMQgqCBdKRL4lFRV3SaWjmlLRmoFpwFvLU2nv8rRh9rr03G0bUsPztJ+e61fJxeEzEebhZXFTbj678pDN47Er+3VfJmACJmACJmACJmACJtBhCPh1nQ7zqDxREzABEzABEzABEzABE9hGIIzm5Ki4PCqG/FFRH4tK7gmSblPwZliWJl5/WKocU5SamzamipEVkadCxnf+DlgZFYM/5/CEQJjAMwIPBfriO+0I64QAoZIfzgnvA0QDhAnuR2xYkuvz6TiSCBsBgDnTN/1SaUf/iA30gScHYgftmL/CStEvHhckAadkc17IyK8wTfTBOeYxLzcuoZ7IabHNw2IbL/pn3PuiTkwNm7akuhWb05bHN6Qti0vSql8uTmvvQvSQUPKv+EworJFRyXPB/Z8P4YJ1veKS87DIJhLf3qc9LF4xXndgAiZgAiZgAiZgAibQgQjgWu1iAiZgAiZgAiZgAiZgAibQQQiEWIHHwGVRCf+EER0DPiGbOI9hHyP76lTz8UGpfmNF5KwoS5UTHwyx4oE4T24GJc0mjBKhmQZHXZCrGPHJ4aBk3fSHcID3A6ICRnU8HpRPgiN/U+hFKIQDBA6EB4WJWhqf8XpgXng5IJQsy/XDeMyHglDB2IgND0VFXECI4T4EFfrEawKvjKznBvcyB+aFVwdtECcOiopYQl+Mh3iCYKKE4azxwJb7iqs2p/LhMZemXqmguFs64JxeqcskBBXl54AtjGENc9hflnsWjP+KSs7LRixfUV++2QRMwARMwARMwARMwAQ6MgGHhOrIT89zNwETMAETMAETMAET6FQEcgby18WiMdDjHYHRHQM6xnqEBwzw81Jh5ZDUZUJFqhr/ZOoyEcP71Kgk4sbQzn0IEIgRHPGmUIgmjOYICIgHtENQ4H7Gk1dCNucEnyUWcEQMQKj4ddRxufkgYByXGw9vB3JsKHE24gRiAH0vjYrQoPwXiBuIKsxT7Zkf4awQJVg3JZv7ghwbtGXerIn8GnhzIHIwL9bCee5hLPpmPl0jTNYzqfrUulS/pl/a9MjgtP7+ramp9qm0+VHmwNqYD2NSYcO518UzuT48LRBaXmmBnT3gXylF328CJmACJmACJmACJtChCdjDokM/Pk/eBEzABEzABEzABEygkxE4LNaLsf3IqHg+IFJg8MdzgOMTIVbUpn4X16Uex/cMsYLf98kLgSBAEu2hUTHcK/zS4vi8NCqGe+WDIBQSY3AfRwz6XFP4KP0NIeFCHhsY2xmD439EPSIqYggiAiGZ8HZAJCCpt4QS1sD9eEFQ8ABBGJgTFY8IKvNgTlRybVAQDRRCKSug0IbzjMsYXCOUFDk5ZkV9JCpeEwgn8sigP8QC7l0QyciXpNL+a9PgS7ulXqdUpYrheIRkGcOcefMM6J9nsquKvSx2FUn3YwImYAImYAImYAIm0CEJ2MOiQz42T9oETMAETMAETMAETKCzEYg3+clPQZJtkktjdMdbAuM/HgQ9U+XYxtT9sHtT5fDxqdfpq1JxL37XR5zA04GCQR7PCUQARAJEDISOhVHxIiDsEoZ4eSzgySAPCu7PhoPiu9plX4JCKEAg4BzjI1BQmC9zwTNCwgjeIbRDWEA8+FlUPCHwyCA5NkKAvCmYKyGhWCtjcB99cl6eFhIw6J/wVayRdtxDP4g0M6PCQeslJwWCDJ4YzG1S1LWpbEhTKihYkvqcV5NKut2bVl0/IW1ezHqYM+IGAgjiyXlR58WzWRdeFuS52OlCWKhMLgv6UV6One7TN5qACZiACZiACZiACZhARyNgl+OO9sQ8XxMwARMwARMwARMwgU5HIAziZ8WiCaukBNb3xOcTo9al4h7PhhfAqFTWf0uqPmVlhIHqkroe3isVl9MWAQKjPiGLMNTjKYBggeEeAzyiB14RFIzweDdg3MfQj9iA0VyGeoQBRACEB64hWKgSaon7uJ+xaEsIKkSFmqh3R0VwQZjA6E9SboQF2kho4N6noiIwIC4wN0SEGVERVhBUmA9iBHOib+aDgKGwWJoPfTKOEnrTz+NRlYuC+5kL90rgYA2MTz6PSMS9eWGqfbx7aq4vTxtmVqTHP78qknKTUwPvDPq9NSqiCiIQfd8RosUNcdzpEoKF8oHIa6TJSbd3GqdvNAETMAETMAETMAET6IAELFh0wIfmKZuACZiACZiACZiACXQeAiFWnBarxbMCwWFiVAztiBBdU9Wkran6hLLUZXxjKhu5IXUdU5AKuj2ViisIwUQ7jPwY5QljxBHDPYZ8/g7As4Ik1ZOjYoCXBwUeBxQM8fKi4BqflXhbOSU4J1GDvrmHI8Z/hJGa3DxoT24KxA7EBe4hHBWeDZyfn2vH96VR8QphHggSCCokvGYt9IMwIu8D/T3DPJQgXHOOUy1rkicHYyNyMDfWgXiBN8eQqGLD3Omb0FQ9U2Pt+rR1yaq0eUHPtGVJr7T06s2p/lnmwDwJVSXR5OH4jOByU4gWNzLwzpacaKG5I1hIvNjZLn2fCZiACZiACZiACZiACXQYAg4J1WEelSdqAiZgAiZgAiZgAibQ2QiEWHFwrPnNUckDgaEd0WJLKh/8eOpz9kHpgAu6pC2L6lLFqMJU3HNWKulLqCMM/Hg5jIqK9wCeExi9Cb1ExYMBwzzhkBA+lkXFm0FJsyUSYOwn5BSGfXkr8PcDoZkQQ+gHwz+fOSIwcJRXAyJJNr+FPCcQFhSeaml8JgwUXgt4NzB3xADG4TzCBWIGuTcQBOTZIcEiG46KeSIiUBASNBfmQ2ENnM96jjAu3hyIKMrbgbCBiPNAKiorS1Vjy1Jpr4rUsL44dZ1YkJ6744m4Rp94YtCOdRHCCo+W/vHM1oRo8e/cmDt7kBBTHAKGGLbalz0wdhax7zMBEzABEzABEzABE9gXCdjDYl98Kp6TCZiACZiACZiACZhApycQhm+M6V+ISjgk8iVgJI8k0CNqUvWZhanHwRjtI/RT97Wp+6EbImcFYgRGc9pyxOCvZNkY9hE8EAIIX4RHwYio9LGipd9twgPGcYz3eDRQMOJzjrGVE4L2iAec4348FBhbeSC4n+8UPC7oFxGASn93REXMILwS99Av7RFQJCogqJALAxFDokRNri88LeiTtXCvPDsknDAn5sfY9EdYLIo8L7gOG9YME/4mQkSBCcID6xse9b6oE6Iujfp0atgwOtUu654Wvu/Z9NytJAUfFBWRhLBWzJ+xEFz4/rEQLUjWvVMl52XBulkThTm3KlxYsNgpxL7JBEzABEzABEzABExgHyWQfSNpH52ip2UCJmACJmACJmACJmACnZLAqbFqDPYIDHgFDEi9TuiZDjijV6o+viDVripLlePWp/IRW1NBFZ4FCAUY3RErMMLjWUH4JIzefKcPDPkIAzVRETNojyEcbwQZ/jG668UmRAYZzTlHCCWEBoz5eHHgbcERgzp9yYNbOSI4rzBQGPcZZ0pUPDsQEhAuyFExLSrjMjfaIYaQ5wLRhvUgPjBPKuPRP30wN67xd40ECa4prBWeHMxbIa2UDJzzChWlxOLMn88IEbQ7KCr8mFNJKiiek+pWz0+D37s5DXobnhVPRoU5bRFX4Muz4pnx7Ha6hAhBKChYsUbWzPxhwtqU52Kn+/eNJmACJmACJmACJmACJrCvEnBIqH31yXheJmACJmACJmACJmACnZZAeFe8NxZ/TFS8CTBab0j9LtiU+r6hR2rcXJKKutSHV0WfMGPflcprBkToIsSJB6MSOklGbe7DkI4QgTEdgzwhkTB4IxYgcugtfsbB64DziAAIDdyP4V9CBMIDxnO8L+gTDwU8EeTJgZcBBn+JCxj7KYxJfxjdlYuCeziPaEIh5BV9Mh79Mg6CgMJMMS/EEc4jciBacL/Wqv4lWrAGiQn0L1FCoaSUqJv1MxclIIcJYgZrp38K/RyTiirWpm6HPpPqnnw+nkFN2rKsKa35G+3wtkBYYS2IKwdGHR/PsHt4Wfx3ro+dOiBchLcF90pAYk583u5tEddZUzYB+gvGsgfGTqH3TSZgAiZgAiZgAiZgAnuJgAWLvQTew5qACZiACZiACZiACZhAawTC0H1inD8sKnklMMwvSwecNTT1ff2QVB7RlxrWPJeKqrulkh71qWxgbSoowsiuXBKEZ8J4zdv4ykmBAKAQTRi8EQYQHzCwk7+B5Nd85hpeBxSM4hIz5KHAcVFUxAP65x4l4cZozr14GHCNUE9cz3p0K3k0R+aJoKE50g/eHxJSCKvEHPHmUMtZi6MAACAASURBVPJw2hDGihwS5OdQSCr64+8aJQCXWJE14me9LDiPECKBBIFF+TgQJ6jqT33wvUsqKq8Lj5amVLvy+XTAa8dGIu65afNCMSO8FOG4WBvP7rB4lvNCtLg1Pu90yYkWCgklnvIYUb+aJ9+zYX+dsHunyftGEzABEzABEzABEzCBvUHAOSz2BnWPaQImYAImYAImYAImYAKtEAgD9/g4fWZUDOS8rT85dZ3aO/V7XV0q7FqQygeVpopwamhuqEtdJj0a18m3oETTeC+QcwEhAMEALwI8KxAlMKBjvMYjAEO//g5QyCbOY7inYIDHgK/CNYQTcjI8k+uTcY/N9UeYKOWEQFT4R9Qjoh6aGzPT1fbQTJyjT0QNeUcgUCCsICawJpJtM2eEFHJM4IWBYME5PEJICI5HidbCkb6yIon6zp7HO4ECH0QLvit0lMJf6cWurMGftrBh7c1p7d2RgPu2FenxK5k3TKmIFcz9oaiIN/D4c4gW83Jj7vZDeFy8QMywh8VuR+4BTMAETMAETMAETMAEdiEBe1jsQpjuygRMwARMwARMwARMwAReIYGpcT+CA+LBiEiovSF1P/yAVHFg11TatyCV9CpJxV03p8LuhEfCMI+wgMGcvA9Lo2IsPyGqkkAjYhAWSqGSMKpTFEZIxm36wSDPdcbmvMQNDPsY9PGuoCAoHBwVYzwCBuMzLnNSzgXWkBUSNL6O9IOoIhGFvqgIAvLWILQSXhcIFXgvyCsCgQERRnkqaI/QkPWo0DiteSJk29IXfxOxRtadFTiy82e+eF4gniCWbEpVM8pS+eCYY93q9PjnEHNYMwwRYhBWEFlgwzPdY4JFCBT2quBpuZiACZiACZiACZiACXRIAk663SEfmydtAiZgAiZgAiZgAiawvxEI7wo8EiZGxUsCAaIi9Ti6KlWOKQixYmuEIypNdStXpoLSZam4EkM73gkICXz+UdTfRcUrAQM8QgVv+3MtKxKALRvuCeM9XhgY4nWUoV4hlxAzEBIwwpOzom/Uu6M+HxURQ+GhRsdn/r7AQ0SeEK09JhnUlYeBsREkGINriBTkhMArBNECgYB1IhiwJpJzD4xK+ChKNuG2/r7RUTkrsucVHkqeEQgtCA3LomY9K+S5whjZ3BjMp28qKS1MxQcUpX5vGZKqxiK+wB5PE9aF+MEz5FlOzD3b3HR9MAETMAETMAETMAETMAET2BEBCxbeGyZgAiZgAiZgAiZgAiawlwmEQRsD9/lRB0XFOD8y6sY04K39U49Du6aGDUUREirM4MO2pKIWOz0GfrwM7ot6T1RyPdRE/VRUklJnvQOyOSi4V9ckZsioLyEjm1eCz/qOQIJ4gfEeYz9H5ovoQV8IDidFxaCP90O+x4OECs1HfXMffSOYUBEjZPSXGMGi8WDAgwNRAfGCuejvGY2lteSPhfcGRbkg+MwayDlBH/LuILwVQoXCaTFedh3cpyTd3VJhSWEqHVSVxl07MpUNQEyRhwlteIY8Sxidn3vGuWn4YAImYAImYAImYAImYAIm0BoBh4TyvjABEzABEzABEzABEzCBvU/g3JgCiaQxzC9sMXL3f9vACP9UmgrKClKXcY2pubE+lQwoToVFf4/rGP0nRSVPAp//GlWJs5WvIRsWiRXqu8IeSYhQ3gZEAn3mmM13h6DCOQz6c3Nj4QmBOEJ/eEJg9Ff4qPyQTPm58yQoEEoJ4QAPBYz8GPjxdqDytwpj4oFBwaMDPqwTYQDRQmvhukJD8Tm7Fr6rj1xXLQfm+8+ocEBUQGjB24LPiCEIQnh65K+FuW6bX2FxzKdxc6ocVZXG/rAozT6dtgo5xXqeigobhBie8S+yE/BnEzABEzABEzABEzABEzCBFxKwh4V3hAmYgAmYgAmYgAmYgAnsRQLx5j0hlUhSTZ4DckJMShU11anPqwekprC7F3UtTIVhmy8duD7EigVxfUpUDOFfjDo96mejEo6JN/zxbJA4IM+AbFiorLcF1/l7QNf1t4HyPnA9G1IJIz2CAoIBcybsFPdgoKcdVbkglABbgkJ+Pgi+k+MBoz4eDQgQGPWZP54UeFkwlsJRMRflrEB8kJgRH7cn8pYAo3Vlr2XXovUxBiwZmzk8HRWPC0SUW3Pzk2cGbbJ5P5jDNhGksKg8FVQ9mbpOGpx6ny6BhXmzHkQlninP9ojcs265zcUETMAETMAETMAETMAETODFBCxYeFeYgAmYgAmYgAmYgAmYwN4l8NUYnjf5p0UlR8Ta1PvsLqmoqi4VxK/rmxeGIb304TCMIwZgbF8SFW+Ds6KOi8ob/xjK+d1eggQr0neFVcLgjgE+K2hIWMiey96bFRoI3UQoKvJsDI2KER+vBCpjIGKQt0HigDwNZOjnPOPrO+LA0qgIISuiKgF2/lwQLhAr6B8GtEXs0D3MV14Q9LGjtWT/9qENybFJ6I1ogfiAxwYeHIwxPved/hBVGFthsCSIcD+lIBWVlKbCPgWp1/HyUGFt9EMbninPlmfMs3YxARMwARMwARMwARMwARPYAQELFt4aJmACJmACJmACJmACJrCXCMQb9xj+N0VFDPhX1OWp54m1qeu06lRYui41125Oxd2fDfFiWFx7OCoiAQb8i6MiHOCZwXdKa14MWW8JDO14JjAWhnj9LZAfJjabswFxAZFiaVTEBgzweFbgOUBSbK5zjnlJUJBQQnvlqWB+CgPFOcItMe+aqHhUEHIKjwSM/ApHxRwlEiBq0IZ7EEj4zn0IA4Sm4j7KS60lm+dCAkd13ANHRAvWw5iP5uaHiIFQgkcJAgmfxYxnxljwZexeIS7Vpeoze6SeR/OdBNzMD2+N5VF5tnDflHvmuen6YAImYAImYAImYAImYAImkCXgHBbeDyZgAiZgAiZgAiZgAiaw9wi8LobGUE84p00tORHKh/RLzfVh9C7okSqGF6WyYc3hXUFSbQzneFPgFYAnAzVb5C0hjwqM75Rs4uxsngeuSUTIP0r84F4Z7hEmxkSVEIFHAsZ5BAQl7M7me+Achn2OiBn87YHhH8M9HiLMjz64zpo4T6F/mDA2a16TG0NhpxAruE4Yp6y4grihZN/0o2v5nhVaW+/c/BFbxGhyfCa8FqIJoZwQlCgIJXhacC9jMD7zYM7w2ZiKiqtTeU196vfGPmndvWNSUx3tyUtC//TDM0Zg4ZlfnevXBxMwARMwARMwARMwARMwgQwBe1h4O5iACZiACZiACZiACZjAXiAQb9qTjLlvVCXJrkllNQWp92l9IolzSSosqUgFxQsj3BCJoBEnCFOEFwDGc0IXyXsiKxYoj4PCLkm8kJDASpW3Ihs+SgSyIZU4Rz8Y5R/JzZXPCAoY9BEIsuGm6I/cDdzDNQQFjrRnfMQKrv076rLcNTwRuIZwQV94JSAGKOySwk4pnBVtYCFhAgGAOSlcFu0pjMn51v7eUV4OjcHY9IcYRD+c57kgzrAG+oIL80KcQKhAvJG3isJhFcUzK0hdD1mZehw3IK4jWMCDPmtyc2Hsvrlnn5uqDyZgAiZgAiZgAiZgAiZgAiJgwcJ7wQRMwARMwARMwARMwAT2DoGjYlg8D8hvwLE89b9oQIR/akpNW+tTw+bHItE2RvexGLmjEhIJgzcGe4zmEjqYPYZ6eRTwXWGZ+CxPi6wYgeFdXhXyOKCtEmhzjfYY7PGGwJiPAZ75YOCnHfPB0C+Dv0I4KYk1icERJp7IzQfDPSGS8DQgBBN9E86JZNcU+qNwnrEIG8V4fFfIJ/rG4wIhhPUjCCAoIIYoMTaeERSYSrjJnWo5SOjhPiXwxpMDEWhw1JrcvZyjZpN4M648MrgX8YjrnOf7ilQ5pjL1fxPzgQfhtLY92xc+a569iwmYgAmYgAmYgAmYgAmYQB4BCxbeEiZgAiZgAiZgAiZgAiawhwnEG/bHxJAHRVWIpi2pfHBFGLurU0HBltRctzZ1Gb86FZURtgijOW/3YyjnzX0KBnC+YxTHYI6xXJ4WXFd4JQzm8ijYkbeBhAvuU2gk+lqY6x9PAkQSRAuOtEFAYEyqvCyYzx25eUno4IjYgnAhcYP1IILURCVUEp4MElwQERiP/hEwmD9tuc5YrAsWFAkwiCC0IWzW4qh8l5gj4UaeF/I04bzC4zIWnxkvG04L0UTtJOpobMQN5QRhzggnzGdUKirdmnocNj8VdyF3BeIJ3OgfUUOC0EG5PZBbig8mYAImYAImYAImYAImYAIQsGDhfWACJmACJmACJmACJmACe57AuTEkBnw8DQj51DVVjSlsyV1R3GtjqoiQUEU9MHJj3MfTAGM6hm+M5BjxKby5rwTVGOiVwwLj/b1RCVuE0VxJtuVpIQFDAkf2O/3LK2F4fCbkEgIAfTFPxmNeiAcSS3QP/SHEcA/XEAKYO/cjvJA0nLYY/VmXkluzHuWyyIZyQmTA+wIxgFBRXONI4dzAqCSz1nhcWxSVvBlag47Ml6LvysOhnBR4rGgdtFP+jGxuDz5zH2IF6+MzhfXQD54k9NM/lQ6tTF1nwGxBbj48A+YHQ545z5494GICJmACJmACJmACJmACJpAhYMHC28EETMAETMAETMAETMAE9iCBeLN+agyHwRuDO8ZuhIiqVDWpeyqujNwV5b1Sad+mSLTNNYzvhFDCwC8PBYz1ylWhMFCIA9Rbov4x1/+NccSozn0IDSryFsB4zzyyfXENoUDhkjDOM79Zuf6V44F75C1AWKcVUREe8EpgzggJs6PiQYFnAYILAku/qIgT9M85PEb4zr0Y+xmbyjgIHNxDn/JmYH4KRcU9eGcgBOBZMTMqwoiSfLM2RAR5VSi006o4R1iprBih3BtxuqXoHrHKz/fB2GIKC0JDjcsdC+PZjUn9LkKwqMmtgTUyBix5rjz7xtxe0Jg+moAJmIAJmIAJmIAJmECnJ2DBotNvAQMwARMwARMwARMwARPYwwReHeP1jIphHmM+9enwrlidig8oTMU961JhFzwCMO6TZBsDvXJOyIsiG/KI6SNo4MmAgZ97ro+K5wFFRnf97q/v8s7IhkvCUM95xmMM+sPQflzUmtx3hY1CdFCibUQRiR8IGPTDvcx9WK6vkXHEO4P7lfcCYYJ+aKvwS4SdQgAYFbVPVPjkJwNnXbQbnbsXrwV4PRmVcfBkYP7crzBPEijkIZHvPZHN+0H/ynUhjrSXJ4i8KtSGo+ZYE5+7pL7nwWROVMQN8nngLaLnrWTi7AUXEzABEzABEzABEzABEzCBHAELFt4KJmACJmACJmACJmACJrCHCMQb9QgL/A4+MWfEXhLHrals0KOp99lDU/2zDanumRXxhj5GbgzeEgIUrkg5L5ixziFUYKgnHBIeFo9E/WVUwjEhBiBAyGNAK8W4Tl9U5aGQ8R1RgRBG3Md8ESzwhJCXg/JjYHTHK4Lv9IERf1BUBApEgSOiIkTQB33Tn8QRPmPER1zhM14ZzFUhmySmIGgwNmPIy0FtNK7CSMHgyNw8ERmYb77nRJxq6QdxQ1zkYZJN0J0NjYUwwvwUikt9yLtFf1OxTtYLv96pqCtjkMOD73iBIF7Ai2fO2tkDhbk9QZ8uJmACJmACJmACJmACJtDpCViw6PRbwABMwARMwARMwARMwAT2IIFjY6zpUTGOY0zHyF2Xus8YnupXrE9dJtambtOV7wCjP8ZujOAUfndX3oisAIDBnlwJtMdzg0TPGMMPjKpk3Vqi8lVIEJD3ga7L+4Ix+SxPCPpRCCR5e6gNhns8IpTXgTUp0TT9SxDhiMEe4z/hkqpzc2W93K85ac0SU+CkkhVelOODsFMIHydFJdwT3hXMW2NpjRI8EIEkzogn/XNOwog4IZjQp7xOsuGl1J+EC11jXsz5qHRCM2u9Pbdmko/Tv0QgxmAvHJtZnz+agAmYgAmYgAmYgAmYQKcmYMGiUz9+L94ETMAETMAETMAETGAPEzg9xuNNfbwByGUxLvU8sjRVv6omdZlelYq6EDYIjwJCKWEsl1ghAzuGc36Hl5cD+R3wqMDLgnBDvMlPMuvLoipHBUm4KfSh3//lYaFzWY8CIdGYfJdRnj4Zk7HWRcWLA68J5bTgiHcDORoQUjDe0zbrGUIbvAzIe4HxHqFFYgzt8UqAkXJ1MA7iA3NW4vDsWrgGL/o6IFfJZSFhgPln/+6R0KDk3PTPZ42TzV8hLw2uMzfWmu+tQv8KL6Xk58yTOQxI469jLTxXng39kOuCZ88e4Bp7wsUETMAETMAETMAETMAETCDvF3cDMQETMAETMAETMAETMAET2MUEIuQPhu4UR8QGPAvwfECUWJ7KB81LA941KJUNKUpbn1qQSvtwnXbcIxFBM8omgMZbAUEAozcGe3I5cB+eEORzUILnhfGZnBISLyQ80KeM+DK263u2rbwOJBggViCiUBlLNWvkR6zAw0LhqCTQIGSwPgQUvCBoMzgqhvys6MHcESDk1YC3BN4Y8iqRkCI+3M88FJKJz4ggSgq+PD5rfgqDJeGBOTInCgIRDJgfzOShgSAEZwQN7ucerombBJCs1wv9MJ/pqd+bxqYJvyZUFuxg8WBU5sQeYC+sze0N9kjLXnExARMwARMwARMwARMwgc5KwB4WnfXJe90mYAImYAImYAImYAK7nUAYoGXEZqxzo2K4vj8qhu/1qfeZh6Xmul6puFtp6joRQ71CFGEUxxCvIs+C7HfaYMznrX2M5xjDyR9xSFQ8MJRfAuM/RSGd+My8uF/jZY3v8paQQII4IpGCcEoY+wk7dUNUeU/QlnYU5sPcEQAwwCMgIEzwmZBVCAKToxLGSWGvlFhcnhgIGlStUQm+6VPz15E+EBNYMx4WEnvkhYGAorXo7x/lrWD+CBJ4fDA2wgRM8PJAyKBfQk4xLt4keLJwL2uUiKPwUcyHz4wvQYmk30+nimFPp8Hvh8GIqHhXSERiL7Anzo29Qiliz+Q+t5xwMQETMAETMAETMAETMIHORMCCRWd62l6rCZiACZiACZiACZjAniaA4b53GKBJwDwyKgZ1DNTrU0nvganLhMJU3KMsEjSvT0W9MF5jxEcUkAAhQ7vEBoVyYh0YzDGs85b+E7kj5zGYE25peO4cYkA2lJE8ArJ5LLJ5Hugja4TPho1SQm4M7uRkQGTJemjQD+NxD+tlLYyDmKKcF6yR+wmZJI8FCTtKvE0/CB2IBggRiAV4JSAcIDIo1wRz5V5yYCDeSCzQGvPXovZwxOOB/hEX/p5bB/1zDmGCMWgn4Yd78fTQPYgZ4qqE3fr7SqG8YBHPeVq31G3GhlR9Os8fFrCDAXuBc7Bij8Cka8GJDOViAiZgAiZgAiZgAiZgAp2PgAWLzvfMvWITMAETMAETMAETMIE9RwDDNW/ZI1xMiIqRnLfsG1Jp/54hWmyMsFD1YXIvTUUlR8V53ubH2E64JO7lTX4VhAEJFxjTMXgTdgjD/rSoeC9gtO8RlbwIGMUxhGPMRzjA0E/Jhm/i7wFEAhUJFcopkc1jwdyZz1NRMexjzJfHg/rlyByYJ+MzLvNjbAkNiAqMg3GecSTQMBaf5VVxY3wmfJIEEXjcmesnG84qK8BoHdlwWtm16DrhqXgmCp2FaLAstx548Z218RwQEvBaQazgHuURQYzIeqbk57Fg3ZTRqbBoYWpYW5BqPtwtlfTCi4MxWCd7Aa7sDfpmr0js0Fx9NAETMAETMAETMAETMIFOQ8CCRad51F6oCZjA/k6gsKioqN/AQUNGjRk/cezEydOqD+jbryDK/r7utqyvpKS0tN+AQYTicNlLBLr36NnL+3Evwfewe5sACZaPi3pJ1IOjzojKG/qDUtXoxrRlaWXauqwuFZTypj6eBxjyCbeEMZs3+GXcZx286U/h33aFTqKNEk5j+F7a0ve2t/gRM+Q5wb14Ekis4Kg8DK0lpNY4tNN1+mNsxuTcX6Kuiqrk1VzLJsWmD4z+rI11IGRgrKcolFTu6/ak3oxH299FRWxB9Fic6wNDPkID3iQINjDQ+pSbQoJLNq9Edi18Zgz6ZRwYIJLMjwp3WNI3wgHrRZyQl4j4c5+EHq7DQ2NoXMZg3Ygdi6IelgrL16Utj22NBOvj4zvMeE7sBfYEe4M9wl6ZlOvPBxMwARMwARMwARMwARPodAQsWHS6R+4Fm4AJ7E8Ehg4feeB7L//MF+9e8PSG+x57ZsuN985/4n9vuWfOL//vzgdunbXo6dtnL3nmo5/9yrcH1wzH6LNflPd9/Kov/fh3f/tnexbzxre+6/1wac89+0PbHr2qe//sD7fcPXzUGAyme60UF5eU/OVfDy/5wBWf/+pem8R+NvDp5134pp//5e//3s+Wtb8uBy8CjNfkbEBQeDgqb9dXpMpRhan7jKJUMaI0lQ/HGM51Cm/3YzzHwK9k1JznOwIAdU1U3vjnPnJCYKgnDBSeFnhYYAzHmM79CBW0U24H+pJhnfMY3OmTPuSFQRv+VsgK39xPaCaM+ogG3IcAgZAg7wJ5gCi5N3Om4D1Af3gUMM9RUREGmJ+EB3JWsG6uswZEG1ggHCAawOeCXB8KO0XfCieluSoHBeJGNsl4NkwU55kb+S/wsrg4KpwQGBSKCo8VQkPJy4VnSQgu2jFn+NMPz5O1UBibdTI2niicZ5xnU98LH00FZVviuddHzhK4swbuZU+wNvYI/eHV4WICJmACJmACJmACJmACnZIAf3S4mIAJmIAJdDAC0w454uh3fegTV3Fk6mtWr1r5v9dd/53ly5Yu2bJ506au3br3GDCkZthRx538qgsuftu7znndxf/55Ss/8t7f/vwn3+9gS33RdA8/5oRTNm3ciMGozWX6oUces3H9er0B2+b7OnrD408985zJBx1y+KaNGwgbs9dKzYhRo7vEpqyvq82Gjtlr89kfBj7u5NPPwqNqf1jL/ryGyFuhBNOEesLLS4ZujqtTxfD+qW7thlQ+AgM3Bnp+N8czgrfuMfBnPQgwtmPcp1IwrMsbgXYY1REBMITTB4Zy+sTQz+dswm3u5xyCAMZ6DOr0wRgSH7KeGLkhW9oPiIqIQN/8H8S/rXdFPSzXB2tWoU/WyvoQVRAelkZFFMEzQwmyuS7hhbwbv4yKBwTiBnNifsyTtdCnRJCsAJEZdrtIwL85EiwU2kr3wBqWCBLypOA74jYeDpyHMfNRPxzlZSJvFeaC0CKRgbXQD6ILHjN4V9CmJBWUDEiVoxtScfeyVHlgl7R+Js8ZBqyJftkj/FzPZu9EHguYuZiACZiACZiACZiACZhApyJgwaJTPW4v1gRMoKMT6Fnd+4BPfeU7Pzn6xFPPWPTI3DlfvOKyd7/zQ1dcdcOvf/7Tb33x05fnr+9rn7n8g8edcsbZH/vcV6/5+Be+8b3GKH+4/tofdVQOhHYaNmr0WNbbnjVMmDL94Pvu+vtt7blnf2g7fvK0GStXPPXkqqeX85bvXiujxo5vCW8yd/YD9gjYRU9hysGHHfn4okcf2UXduZvdRwAD/1lRJ0ZFCODtewzS28I8rZ9dl3qfWpwaN5dFjoOn45zyJtTEZ+5FZKCtjO28ka98DAgUvJVPwm3aIeRi0MfIjcEcIzmiBAZ7BAIM/tzDOQQN+sG7QAm14+N2r4vWxAquS/RQzovj4xyGe4mRiCzytFBIJOZEkacJogocONIPc5WIgIEfDwuOtFcoJo54LMiTQlwULivr3SHRhfUpqXdWrFFbxuZzTW4cmCDGKD8Fgom8TbjGedZHkbjDZ8bjuSlZOOdYH+IDIgzc8YbpmwqLG1Jh1aDUXL81dT+kVwgWrJU1sCfokz3Cv5f0OTM3lg8mYAImYAImYAImYAIm0KkIOCRUp3rcXqwJmEBHJzBu0tSD+g8aPPSyt7/p/NeefPjkBfPmPIg3xT9uvfHPO1rbHTf95Y+XnH/aMc8+s/Lpj1715W8NGDSkpqNyGDF67HjCCy1e+Mi8tq5h0NBhI7r37FU998GZ97X1nv2lHfvl4Vn337u313PguImEOUnzH37wgb09l/1h/IGDhw6r7t2n74K5c0hG7LIPE4g35BERyIWAYZowQxjQeRO/KZX07Jl6HlmaGjasjfBAGM4xbCNAYLTGiI+AIYO8wgzhzUDFa4r2GNDJ70BYJozrGMgxdnONqpBQiBf0ReVNfqpCIUFQBvhs3ofWvBfk4UE/GPTxQEBEYc6MhRjCGuiPNeV7a/C3B+3wWsADQcm2FeKK+1nToVEx4tO3RJosP8Io0Y/yVmRFF+Xc0PwV1iob2oo1wxSxRYIKTFgfbFkfPPms+1gL40mskfBBXwgaWXZaz9259eg5NKfCCAmVijanbkfE2IV4qdAne4K9wRrZK31ye4e+XUzABEzABEzABEzABEygUxGwYNGpHrcXawIm0NEJ3H3HLTe+9qTDJt32fzeQjDSdcNpZ5z2/5tnVL2eMf3Lpkseu/sRll5aWlZe/9X0fuaKjchg9buIU5v7YgvnE+25TwbuChg/P7lyCBc965JhxEx7eB4SaMRMmT33u2dXPrFz+1LI2PTQ3ekkCE6bOOIQG8+fM8hvYHWOv4AlTExWBAMM2humKVH1qn1TUvSTVraxPBT3wgsLgjQGbHBEU2mFQ15v7GNgxaMvjYml8xjBO6CJEEQz9XMPoT1+IFwgZfEfkwMBOHxjPMc4jaHAum6SaceXNkZ88m2v0ryTU9IERH/GAtTHO8tw5eSnIiC+PDQkaGOXJscH6NB6hpBQiijWzVuagPhBd+MxaJIgwp2yejexa9Jk2ra2FsXVe82MtykuBRwdcEUzw+MA7RR4e2b+huBfRQ/MgPJTCWJE/SsnBEWjWpZIes1P5wF6ppHewa4Ib/fOs2Rt8r4m6T3lPNTc3p1wtyBz53FotzJ1vOQLfxQRMwARMwARMwARMwATaQ8CCRXtoua0JmIAJ7GMEjj35Va++6/ab/68pystN7bYb//T7Rx6ekNz52wAAIABJREFU/cDJZ5z72vKKCgxNHa6MnTRlOpNetGBemwWLSdMOPrSxoaHhkYcfmtXhFvwKJjx63ITJeKPMn/PgXjdqjxk/aeq+MI9XgHOfunX85KkHMaF5D826f5+amCezIwIYwSUgIBJg9C9PXWeUp4bnt6bqUwakolIM40oujSEfIUBv6WPolgcBb/3zGUM7bTCOD8wNjEiAkR0D+dKohIZCBFBYI/rDOL5t/G1F3gj8TYBIIPGAa5zLCgOck2CR9SbI5sd4LDcu85CBX+MwZ9pilCdckvJQ0CfiBP8vydME8YXrEik0N9aAN4LyYmS9QLSW3NJahBV5QdAufy2sT1X/h0q44DzhoSi6xrjio77Uv/6mwkNDycWZO2uGP5421KpUUDor1a54LnpqSkMugwXPAgbsDXnIsGf2WMkTJPJFCAkx8o7Jftc5WMOG58K+5NgiWkXfRVEtXuyxp+mBTMAETMAETMAETKDjE7Bg0fGfoVdgAibQSQkMGzl6LOGO7rz9pr+2FcGNf/zN9ZVVVV2mHHToEW29Z19qN27i1OmrVz29Yu1zazCGtalMmHrQIRFBak7t1i0y2rXpvo7eaHx4liBkLZg7e68KNSSG7tGrure9AXbdjiLU1/p1a5/Hc2rX9do5etIb39k3w1l5/pviu5gGoZ0QDvQ2fxi7CzamsoFNqevkbqm4a2MqKsZgj8GXEES0k5eFjPkYuyl8V1Jn7iE3AsZtPBbwbpAggFiBVwBtJH5gTNfv/oyhhN70ixDAvZyXEZ72tMl6J2TDINEX32Wk5t/YqblzGKtlrMcIr7EQJfiu3BrZ8E18ljeJ3syXWKCQVtxPyKnsm/uac/Yc3grKq5ENDZX1wMjm2lBeP/XBNeW94DM8s94oMJMIwues0CGRhTk8GvWe3HNYGsdNqbjLsanLpKpU0rckFVbAWCG06Ie1sFfYM7u9aN/n1iJRjHUrxBdHmCt0FoIX3/EE0t7Kb89+lDCnEGQtScdz4kVWEGnx3HAxARMwARMwARMwARMwgSwBCxbeDyZgAibQQQmQeBuD9H133nFrW5cQiadb2k6YclBLmKSOVIqKi4sPDK+B9sTtLy0tKxszYdLUubPv73T5KyZMnj5j2ZLHFm7auFGGzr3yuBGZGNgeFrsGf0GU0eMnTcG7Igx9tvTtAOuOwtdE8xZjaRz5HbglpwNvf+e+y7C9/Y3wVkLe7IyBFcM5Y8iD4PlU0r0yrb6hKd6035IKu82JaxjEKbydT3u9rS5jNm/3UzAcK38EYaR4Ox+hQkZkhA68qvBgYH8QPgnDMvdhZJZhXW/E06dyTeitePHRd+WK0L0cVbmf9kpg/c/4TDgjqjw0EAlYB8Z4PEKYMwbtrJeG5iGRIJtoXMIIHhsU5kWR+NBaQm2tKeuBwT3620dr0fwlRnBEBJJQo/sREbLeGhI28oUOviuMFWIE+XuUSJ35EyJqeSquXpqaa6O/xqJUNpRnLkGE58gcJbbklrprDplQTS17PHqFnfZUa/lNuIYXCPlKFHKM3CJ4BHEvz5HrCBJ4+pDThPPsNdpwHXaE2aJNPsP857NrFupeTMAETMAETMAETMAEOjQB/ZLdoRfhyZuACZhAZyRwxHEnnYYRmDet27r+pY8tXNDU2Ng4cGgNCU87VBlx4NjxZRHLqj0eA2MmTp5WUlJaui/kcdjTsPEs2RdCBimMVzh6OHzRLtgEA4fUDO/StVv3uQ92PhHupfBlYuXLIK03+mWYxkiOAZmCkZTPGFZ5YxxRj3P8XiwvBAy1MhrLIL49bFBOLNouGIWO9FLTOy8uYrilT4zWXVPV2NpUfVppKqkuTUVdxsY5jLqMR5/MCQ8EhVqSEZwx5J2AURxDMfkrMCQjXiAS0BajOOtlvhiamRx9UnY0UeW2UKgjxs56CjAvjOlZA3M2fBTjYqCeFvXHUV8ddXbUbQnGUxqWu5f5yJNCokR2TupTnhc8TyUcR3ihKJxV7uuLDownQUbCirwhEFaUX0Nr5Zhdl0I/qWPNKX+eXNf+yoaIktDD+vB84RrPnT2A50R1KqoMVrFpqk8pSVsXb0krn+AZ4qHCvbRjz1yzowW+3Pk8LROdky2r+cOUcZQfpcX7ISp7X+IDc6Dw+wVCBN/x/oEfogQCBGtjXRKi8K5BnFHIRp7XsqiIVXhdKGcIfcjrp+VnKvPz1PIz9TI/Ty+3fF83ARMwARMwARMwARPo4ATsYdHBH6CnbwIm0DkJVFRWVk2ZcegR9/zztpvbQ6CurrZ2zbPPrKru3QejUYcqkW+75U39eQ+1PSfDpGkzDuWeuQ8+8O8OtdhXOFkM2kOGjRi14OGdCwc1/dAjjyHs0CucRsvt48PTY9XTy59as3oVhtUOV+DQlp+X7j17VZ9w2qvPJeTa7lwkCcxb9vTszrWn85nmx9yP6/KSwBCq8EEcMdRzxMCK0RQjsvIGYIDflgB7m2EdrwSuyWjMfRjHqbShb9X2vBmOwRahAeMvhumGVDG+JDWuK0lNdWWpsAijL0ZczZX2a6NiwH4it3YZ2pkTfVHpi/kQGox7T4w6Lipv9WtdMqTrd/6s0V25CBiC84yHtwZhjPiOaEHSbgkX+YZ7CTbZ/A2IJrTDy0NGbq4vzq2FdRHSL+t9kVviC0Is6bqEB4ziClGVFSFa83qQt4RCWSn8FSyU+4IxJU61JkhoTtn+s54lWQ8N8eM5StRi/nDDw4X1sv6hOaYNqaBwcdr6eEhUq4pSUS/WyPOVpwXPlj2w0wWDf87o3+JJFD8vrJv9zhgK60TIMPYJex+Ra3RU8nbwM8BxYlTECUQI9hXXR0QdFRUvTfbbpKj838yeo1/a0YZx6XtMVPYRY/OihJLD87PIXLRP871t4pKLCZiACZiACZiACZhAZyVgD4vO+uS9bhMwgQ5NYMbhRx+H58C9/7i9XYIFiyZEUEdMuq039dvjNYCXwaaNG9YvXbxwQYd+4O2c/LjJ0w7ildpH5rY/0fjZF150yZVf/vaPyBNy3ORhGKpeUUFomnnvXf/YmU7Yp336DRi47PHFi3bm/ld6D8LgtTfc+q/6uvq6b1595cd+9dPvf6u1PglX9ou//uP+gYOHDrv6E5dd+utrf7DTb0a/3JwnTz/kcNq0R7h7uT478PWskZPfaRWWCEOoDPMYjRVrH6MtwoUSUWPsx1iLIKGkzwrJw3neKMfrgft4m5zPEgDwysBoLWP4dm+LVnhiAMY4jgF/m9dG43PFqahbY2reioihMDoYqhXCSZ4WjKN8DBh7GY810R9hdzAMMzeEAPpHjMYYzJryDfvyMmAG+syRPpkXlfthRKEPfaadvAR0f65ZywGxA5ECbhdFDWt8OjCqwkHRDxxhmh/KScb/fBFAnhWMrbfzs+KC+mF88ecc68DgL08MecgotJT2Bs9fRSKHrslLQwz1PbtmrvEcFKIK/tl9wD7EOwGj/Lej8pz5jkF/SSofXps2zatPlSO0NuZNH+wB9kybS55HhUJ4ceTngnWydvYFR7w8YMs15sO+ow3fdY1nNz4qHPm5op0ElQnxmb5ZD9e2JRPf1gceNjVRH4jKPmU/0U5rJIE8c2DvImTAm/2rZON6Di/18xTNXUzABEzABEzABEzABPZnAvaw2J+frtdmAiaw3xI49KjjT9qyefOmObPuv7e9iyT5NMbs9t63t9uPnTBl2jMrVyx/9pmVbU5GSq6OebMf6HSx/ieGUEOIjQVzH3qwvc+tV+8DMIqmx3eByIMBH8+D9ohM2fl+5DNf/uaVX7mG8DJ7pfAz9v5LXnf2xg3r1jGXd37oE1e1NpHi4pKSbt179IT50iWLeDt9txU8q/g56KgeK7sBjH6X1Vvj8qBAgEBwUygo3u7mbW/eHKctb5djFMZIzD3E5ecNckIXYWStiYrBdVBUvFpoj8GWI/1igMfoisChPBg7Wp4M8fISKEwlPWLejQ2psIo+8GpQOCDmhjEYIzBiBgZ+KsZmjOP8283amBsGX84fkpsPLJg/a8aQLA+KrDdI1quC+Uqw4DNzoXAvYxFmCjYYk1fl5sGYKvp/hLwZfGZsjNasBQ8txpIAhKBCbgjWJuEla5TOFyv4ng3dxJjKDaFxW1uL5odIoL0hUYn7JFoo6TdzZW6M90RmbVkxivtgoDlo3hyzL39pPlmvDJhi9K+JigfP0twc8LCpSI0b61NBsdYJc62xvQZ7jU1fPH/2BcIcAhL7lb3Ls5B3EecZg/kpfBoeFQgOJ0TFO5GfCfa/8lcQuuyY3Dr4f5g+zol6elR+Lo6OihhzWFR+ZrRP2QuIHIge9Klr7DOEDHlaMGf2f4f7/STm7GICJmACJmACJmACJrALCViw2IUw3ZUJmIAJ7CkCBx95zAmzZ957d0NDvWKyt3no8nhtPCJDyfjS5vv2ZsPCKKPGTpjUnlwUGMoxmHfG0DkTpkw/ePmypUvCuYQ3ddtVfnrN164+/4RDJrz9gjMxWr2iMn7K9Bl0sDOCBQnTTzrjnNcsnPcwcfD3Wrnr9pv/77zjDx4/+/57777k0ssun3zQNg+HbEEEPOeY6WNOO2TckPvuvKMlsf3uKHickES+PYnnd8c89pE+ZXzGQEvFQI1BGCMpIgTeABj1JUQQqgaDOqHJEAAwWNMGYyx7nftpi2FV/65i8MVQT/98xtMBIy1GeT7zezTGYY4kMd6RoZX+MMRijMZoXJLq1zan2pUFqWwwfctzQWvBsK832pUngD4wrjMWBnC90S5RAEMxBmcMwBIoJAJk5yWPgWi2XaxAMMFoz9vv3K/QWaxTxnqMy8yLf1NYO/z0VjztETcQWThizFZYKVjDDIFH7BibtXJ/a14SXM8a/WkHO/qCgUprayGpN+0RUbLX9TeP+mVttJkV9aHcnP+cOxLWSl4njKX9IK+ErKcK15XrhL4lHEh4wBgPW7iyVljl5li4PlWMLk8FbImW63zgPvZKm/9vzySR5372qfYyng01Udn7U6LyHeHuyKin5s4hZhDS6YKop0RFdKAt+4mfJcQGwj4xb+Wu4J6zoiLwcQ5vDIRAclcopwpr5TPhytgP7GP2zmlRWRvneZ78/PBzS5+wa0kAHmvi56klwX2e90hcdjEBEzABEzABEzABE9jfCTgk1P7+hL0+EzCB/Y4A8fRJQH3jH3/zy51ZHDH2N0dcqJ25d2/dM3T4qNEYa+c+OPO+ts5h/ORpLcbyzihYsPaHZt73r7ayyrbDS2Dxwkfm7cy9+fcwD/qb/9AsQsW0qxDOqyqSccz697/ubNeNu6Fx6D5rP3bpW153w50PLnrDJe98X2tsyQ2zG4Z+QZcTp844BG+OhY88jIHVZZvRW/kqeHNcBnaMoBiKMbzyNj+eRhi6MbTTTm//Y5RVDP858RmDPG+KE6NfXhfKJYF3hgQD5bOQaKB/T5W0O//Z0I650hfzKkxrHyhOvU4sTo1bFNpJSb5ZA8bhpbn1YAxmb9EOA7KMusrHICO5rkkAyIoUSiqtecnLgHsxIrNmBAiFIeI8AgXzwIAOF+aO4CPDOqKAvFf4DBO9vY8Ao6ThSubMfHhWjI2BP+tVoNBNWc8F2mktCivFGPkJt7NrYa4YvulfHgSsmbFZj5hIbOF5IlixNq7zHDGks2cYk3Y8D9aHGMCclaxdYZfoU6Gl5DHAOYWhggX7jb7Egn3SIzWsDw+bWE7TBtbNXBgT0Yd1Kuk1899hiX9eJZDAhb2sHCsSSJg3XhQwYZ3yPFqYG49cFKwXbswfcYHnpPBW+s5ekKeIwqexJkI/IfQhOig/CGtAPGNOiGGIVfRHJbwfc6EPhUDTvmN8SjYhd3s9TXJd+GACJmACJmACJmACJtCRCdjDoiM/Pc/dBEygUxI4KPJXsPCZ99z59/YCwFMBz4OwrbY5rFJbx+jRq7r3pOkHH9Zv4CCMF7u08FY5HbbHw2L8pGktSaPbc88unXQbO8MA3cambWp2QN/+A6jzH56NIaldhbwoE3OJyttyI14QLxVeDNHhicWLHt0ZT4+Ro8fxpnsITjP3iYTpK1c89eQdf/vzH44+8dQz8tc8bOTosT2re+8w3wfCS1t4vlybKTMO483o9NiCR+a+XNtOcr3FsyEqhk4MvhhAMX5ipFUYI4kXGI4xuJ8ddWhU/p2iLUZcCkZmBAwEArxoiN9PO4RPBAxC45BYmOTE9MP+pA8ECOXBqODN8Fx/+QcM3eyRbYnA655uTgWlBal+FSKK8i4wByUoxrjL3HkLnfVx5M38bDgk1iSDOUZueVQoxI/mkO/5kRUGmD+G/iVRESYYB3YKC8W9JI1G1CBEFcZvzmF0Z66sS0nJeYuea8wdJvLcUKgjeR1wxPgtbxDGynpa0Ed2LfTPOeaYbcf6sgZt5WuQsV3rloAgzxMM5nhXbEuAntL8qDy3o6Ii1rJ/8gUh2MirJ39chZeiD3lfaP6MwXnm9GRUjPe02ZIqRvZItcubUnEPvivhOnukzd4V0VYeNvQvUYj9yX5lLJ4B+wTPC8QZniNH9vp5UfGoYGzWjdDAvzGIc8yV/X9uVH7noG9+b6Atwgj/LiM+wJznw88IXBHX+LmCH/uoJipc8cBgT1AZmzBSnIM1fdMH3hoSoPLDfcUlFxMwARMwARMwARMwgc5CwIJFZ3nSXqcJmMB+Q+Cgw448NiLQbJ43e9b97V1UvwGDhmBkJgb+y92LIf11b3nHe77/qz/f9tlv/OC6lzK6/se7PvDRWx9Y9PS1f7z1XzfeO/+Jr/zg57/blYm9x0yYPLUpyiMPP/gARvVL3n3Z5T/+3d/++Zmvfe9nGOdbW8v4KdNmrHp6+VPtyXmB0fl9H7/qSz/+7Y3/+K8PXv7pHTEi6fnHv/CN770UQzxZdmTMLywqKoLZzTMfXX7f4tVbv/ajX/6Bdb3cM2nL9XGTprYINQsenk2ok3aVC9/8tkuvu+G2e0aPn8Sb6TssJ55+9vm/ve2+ucz91lmPrWwtTBJrJO9IVjBija+96K3v5LkxVj6fsy9401uu+fkf/vaNn/z6T+w9vDM+eMXnv/qV7//Pb7/03Wv/96Of/cq34dquRWUa89wuu/Lqr+/o/lPPOv91n/vmj36+o+uzw2ulLDY24pzasIb/+fPt917xxW/+oLX7hgwbMer2h5Y8c8RxJxEKJcHlore/5zI4/+T3N915zEmvenVr9x1+zAmnsO5f33T37O/+8oab+RkgfwVtH1swj9Arnb3IeMzvshhGMaZjZMUQzhvjy6LikUVYGr5jdMfYrrwWGE1pw7+F9IHhFbECgyyGU4y1NVEx9GKIxZD/RFSMuogcSsLNc0CE2BbqqfXQUDKcY6jfVkp7xdv1ZQWpsBJDrTwzJFbQP+IEYxGmCQMwIhWG5mwYKiUXzxckNEo2rBIGZAkGyovBumAngzr/ZnCNcRlHyb3JXYCwghFcRR4S3A8L2PBvmEQMjOSMKYEBgzp9cB/PCK58lmiBkT4bwikz1PY393kmEgQkPmSPzFnPUqGjsmGxuAZP9ooM6jw3hCg8DtgfMNW8uVehoTC0a02ap4QVeY5ozjK2K7QT/XE//27wGcN/91RYWhZiRVEqqc6KLtojO3qm27nkvCvgxzgUngV7ibH4fxHhAWGN58LaCOGEJwTrJQwUa4UTz5y5KZxUTXyGC8+SvnleiBOIPOwNRB5Cf/Hzg7CHCKL+CWVGe4lBzIVny7Nnr3Odf8d4CYFr/KzxMykhhLHZ7/lM45SLCZiACZiACZiACZhAZyFgwaKzPGmv0wRMYL8hMP2QI45+aOa9/9qZ/BVDh4/EIJdeLuRP7z79+mNM/fCnv/TfBx9xzPGnn3fhm04/98I3tgZx7MTJ0979kSs/H1GE5nznK5/7JImeTzjt1ee+/pJ3vndXQR89buKUJYsW8BZs+v6v/3zbpR/+5OeGhiH4zNe8/mKM/a2NQzii9oSDwhj8m1vumXPxO977oWnB+G3v++gnh48aQ+zvF5U3/9f7Ptx/4OAdepJgXL555sLlRx5/8qvyb0YI+toPf/F7mD3473vuuuWvf/jNcaeccfbJrz6XGOKvuIyfvE2wmD/nwXaHYXpm1UqMeWnQkBrinLda3vGBj33qy9+77jebN23a+D8//PbXQv8qQ1TIbzwi2EW6lCoJFtUH9O133Z9uu/djn/vqNWec/7qLPnLVV7711vd+5IrsfXjoFAeg+kiyghC1fu3zz/ULzoNrho+sGXngmEFDhu1wXm0Bd+zJp5/1hv985/v0c5B/z5nnv/6i085+zeuLYhKt9UdoKM5nxTtEldWrVj49KDZka/eMGjN+IiIh7RDxvvuLP978/k989ss9I7n5+BCXXvOmS96RvY+xP/mlb/0Q4QYGjz36yFz28jd+8qs/TQ4+JALfFQnR28JrX2qTjWeflytCBlsZbTF0YkQ9I+rxUXmWvGmOsZZrGIT5/RfjM2GgMNhibMWTAgM+Agf/1vCsMRpjjMUQTDv6weCMcZ7vGHgR0BgDA+2ODO4Y65knht5toYcqRpanhg1bUkEZ/WEs5joGXeZFuSM3BiGbMLCzPnmDcF1vovM56zHB96wRXwmnEQf4zPj6TLi1xVHJ2YCBGgOy8n9grEbMYV4YkNnftFEYKQQVjNAUeblgGKct98KE8QixxJr4rHZKup27vYWvEorvaC0aW94jHPN5Zw3/LYkhoogTc2UM5shzxOuJPsi1wTXa8wwx5LMH2Cs8W9pzXsm8WTclO7bEBQz12fOsi2cvDwdEBPrk3IbUXLc1FZZsTbVspxYjv/YHzNsSEkoeRrSlX/ajRAg8Hfg/Cu8G9jDMEbxYjxK783xZOwICXkX8HCBEcF7JwpkTQhW/OyAusBdhQQ6Mk3LzZl/yfBEjGIv5w4GfQwQS+uJ++iEfBgIF/PFWYu6wRgjRPtGejVNOwA0EFxMwARMwARMwARPobAQsWHS2J+71moAJdGgCvcLIOWzU6LEk3N6ZhUw95HCMF2nh/Lk7jIHft//AQT8J74WJEc7nVz/7wbdJJIwIwRvxp7z6/Avzxz3z/DdczFvm7/2P1575w//+4lVvOe+Uo27+8+//d1e+BU7CbcSHj332a9fw1v4733D2KSdOG9WfhMgkmMbQnZ1Xn34DBiK6zIt72sIJUea7v7jh5orKLl2+eMVl7z7ziEkjGhsaGi7//Ne+w9jZPhAcph58+FF3//2Wv7XWN2G3PvP1711bUVnVZVGIOPlt8ODgrfqrPvKet33knW++4GPvesvr1j3/3BqFsGrLfF+qzdiJU6c/9cTji9eFsb+9fTXU17UY5RbnxKEXPesQiN7+/o9d+Zv/+dF3Lz7rhMO+9pnLP/iLH13zDcJIHXTYUcdm2+uZzJ19/31VXbp0/d71N9zSf9CQoe9582vOOGrcwO54v1xw8Vvflb3nMx9+91vffuGZJ3w08kWUlBSX/Ok3v/jZG8849uALTjliymtPOmzSpRed9yqEkvauS+0XzHuIXAapNQ+S0rLycoQq9nLvEFdaG6NLl24toZ0iBwzGte2lPrhJUMu/jz65HiLj3Vdf89PrDzr0yGO+8umPvv/VR04eeeykmt4ffNsbCcuyvVz19e9fe/aFF13y6Q9d+p8Xn33i4R9/z3++kXXzc4lQMn/OrJlNjY3//039nYXRwe6Lx5IyNWuYxjiKoV0ik96yJ0QNBup7o2IoR3zEmK78BBheMbDSF20w3v8uKkIEIoHe8OYehDL65168DRBDMPJiHMb4jSFYgkNrZDFo5z2zsJU3PNuYNj6IcRwPBQpzp0+M5/K8Ya9h0SYk0eNRMSbnC2oymMuIT1/ypuAahnOMwfCg4klxY1TWxpgYsPFAoTIXfsa4DwM769Kb+/QLL4zj8haQhwbznB0VLxf6WJCbg0QePAKZtzw96Ed5JeSpQP/Ztcg7QyKTQj1xr67leyKIdb6gwBphgCeFDOO0xWtDc6J/1iwGnKeNBAT2hMIWiTVHmLIWjcE6lDwbvogCCB2IQQq1tCxtfWJdatzYmDbMyg9zpWdHPy9XNA/2Mv8+IXqx3xEvECeYswQB5qexaI+YwJ7mudCGexAX4IAXhsJ/0S8/P4jhCH+0gxNH2CBKsTZ5zeB5gfjNPmb9/EyxJipeT/zfye8w7BdCUSlsFXNnztnnG19dTMAETMAETMAETMAEOhsBJ93ubE/c6zUBE+jQBKbmYtjvbEJljMpPLVu6hHj8rYHgDXDe5B4Yb9hf8f63X/yX315/He0IQdUSkuagQw6/6U+//VX23gGDhw7DuL961dMtb+fzBjiG+F0FmpwbCDVdu3brfnx4bnzgP19/zj3/vP1m+n/g3rv+gRdDRLqqmfPAv+/RmAqLNO+hlw+bxZv7eGlsjYm/4/VnnfTovDmzMV5juJ4exuVAMXLRI3O3Cw/jwoOhxXNg1v0YOV9UCCvEW/V333HLjfmcCZ30+kv+673/e90Pv/OH66/9ETfrzfuGgLgrmOHxcv+/7uTt7HaXsROnTA9b/HryTuTfTG4SBKPZ94fh/YoPvZt50+Y31/34u4R6QtTK3oOIURsbB88bjPB4R4SYdfQjudwaiDk8O1jX1W7F6Lm9kFSe86EvtNtL5KUWLQGJnBP57Q458pgTFMYs9IoBCCr5bfDMYE1rn1uDYbelcM/w6O/Pv/nlta2NfchRx57Iz+sZ573+oqNPPO3My999yRv+dsNvr6ctPyvZexAq8PD46TVfu/qPv7rux7rG3l762MIF7FX4t/vB7r83YHzFGIxRGYMpwgIGVcQI3jDHUIqh/5dRERV4K3xYVAQOjKvch4GUdspBQj+c5+eRPY7hnZA57G/C2GDkJaQPhm8Zadm/ylOCsX9z/Hg0xj8hElY4hzjA793bQi1tmrMlDfyvLqn7jJr4zl5TQnBEQ+bMv6cIJworpHA+CAAUeQUwbIePAAAgAElEQVTIuKv8CTLg851rtGOejM+aGJ8wQayfcamwYQ14UWCAxtDMXBWuSXkGZOyWBwV98XY9bZkf7eC+NNc/a8DojcABO3lSMBfmqRenMJYrB0lLWK2863zPGvW5V+tTyKc41VKy3+Vpwjn6Z54Y3jGMK08HwgtzhpEEHcQoJe2GGfepXxngs946nONeuHBeRd/hy3xpw/7JCUDN5al+fWUqOYB2iATyLGCstgqzzI9nzF5hLyMksD72KOPxTPi54Dr7mPN4XuAJIY8bCUIw0Frpg3/n4MazY04IZ+w/2snThWcJQ9ZHYb8y3pLc2PAgnBQiEPdwnjkrNJc8j/j5gYGeg0KOdTpxNsfRBxMwARMwARMwARPo1AQsWHTqx+/Fm4AJdDQCJN0ll8OcHRjLX2o91b379J00dcahf8gYQvPbf/qr3/0pwgRvukusIAa/3pZvzauAsD2EsSF8jUSLXcmV0EL0d/RJp53Jm/1/v/mvN6j/jWFc53N+UmfyV2BQj7BIL5l4OjSQHt/48a+iv4ICiRX096owGpNrACHmvrv+flt2PZOnH3I4b7hjiM9fJ/cozNHvfvHTF+U0eN/lV33p+TXPrv7vz3/yI7oXIzR5EbKiyM7yw6uE0EsPPXDfdvGmPX0hMsx9cOa/JUZk733/xz/75dAQKr74yQ+9O/uG/5rI4P6tL3768vxx8NAh8fdRx59yOkb4Kz/wX/8hsYK2JaFy4HmQL1ZwDa8Zjg/P+nerolB71pRt+8SSRRiZ07CRo4jt/oJywqvO2u7psKO8KPBZGmIOP4O6eVx4tLD/H37wxQIWuS4QXxCo3v3RKz//s+9+40sSK/LHj63Y832Xf+aL5Fz5QXgq5V/fEPGoODfrvrv/ubPr38/uw4CKQRbjL8ZljMJ6q5wQRxhxOY84xfPC44h/L/jM2+V85/dghez5a+46mDB0ExYKIzyGUwy3eEJgbKXw86X4/hiJeUuf78rRkP/WP2NSZWQPU/GW4rR+Zl0q6/d8qhihHAI8Y4z7vPXOW+vkKiFJOGtkzggZXMeYrJBHCrXEUcZmiRgYf/HYyOYD4BrnEG5YHwzpV6IKR+aqEEwKqaS3/vnO+NyHMRtjNfOHD/dwf01UfnYJAYT4iZGeOcioTf94ZLAWDNZ8Z+7MQ/lhsiKBhB+dk7E8mm/3yMh6aTDHrLcJXBEl2CO0w9sBw7vEIAQc5oNRHQ8K1qYx5BUizx3mos+MLw8TPrOXxIt2yunBs6Mf2iIYsPempYoDq9LG+ZHLpAIGMsxLnMn3uqD//CLRB+4IboxDhTXjIAwgKGjPIBIgJiA8KI8HghXzQsxDXMLbgTnAh2ehnEFco29Ysj/FG27sBwr8YECtiSpPFubAfmbf4Q15SFT2C54WzIVnwzzwIJIg5ygAOag+mIAJmIAJmIAJmEBnJOBfBjvjU/eaTcAEOiwB8iwsfnT+XN6Cb+8iXnXOa9+AYfWmP/3uBR4S6odEwCefee5rf/7Da76ut/+59pZLP/gxwhxhvMejIX/c++6641bOHXXCKae3d05taU8ILNptWLdu7Te/8KmPZe+JSEMtbzXnhz8aN2naQcseX7woX8jIH48Ey7w1/4n3vvVNeFZwHdGBNfOZPBD5fZBH4Ikljy1szdB++rkXvLFmxKjR3HPnbTdhAN1eEH14ftd+77+/nA1r9Nb3fPgTPM+/3/T/hZi2cGmtjQz98Rb+Xe3tg3VPmHLQwXNm/X9PFfWB0f2kM855zV9+d/11+Z4UrY0Tj6U7XgyPzp3z4Ic+/cVv/OOWG/9MeKds24FDhw3nGbV2P2GUMNyvCHeg9q7jpdrj0bAmEk4MGTaqJZeLCh4ix5965jmE0uIc3iT5/SA+4Lkz675/vUAw4LmST2b+nNkvEsf0PPCsWLP6mVXf++rnr9zR/C5489svxZvoe1/7wqfwaMpvF1rUQH4GdzYc3K7kuI/1hWFYb/xj9CQ5NQZbMcQYfWzUU6IiVGEQxSsALy0MuH+PSlga/i05OSrPXoZajKnUlm0RFQM8b7BPjIo3AoIIxlsMxhhuMUrnewNwrzw5FBZoawoHjFQ5Mtq2eCpJUOH3cuaknAB4qiEKUDH+YjxWyKPctLaLFDLmI1JQ6EtGcu5nDAkXzFF5NTiHIRphmHXXRMX4jRFdfyfozX+9kU//rJc+EHPoD0M498EIAzT5CTgPH9jJQ0HeEYgFEiLol2fIs5F3ha4pLBNtOKdE4VmDvoQr5kWRIV/zZywlKMdQDkcJEgqZxDwxylPkJaFnQz8Y/zWmcjRojsp9QigkeWZJ6KAt/JW/A9EEHsvS5keeizwWTal2Ff0gGtAPewShI1/00tqyR4lIWgvjsO+ZK9eWRkWYQEhAwOAIZ/YrwgP/3vHzgjBGW+bK3mZs2sGJfpgbQhTCBHtTXhD0gTCFyEGBs3Jv0BdjIlRwVNJtrvPvPucRbtjXrJf9xO81Wc8h8c1174MJmIAJmIAJmIAJmEBnIWDBorM8aa/TBEygwxPgLfwxEyZN3ZlwUBijz3vjW95OOKjW3tAmpNI7L/v4ZzBGf/MLV35UsEgkfMa5F76J74+FUJIfwobzt934p9+TjPj86H93QFb4np//6Jqv5ws1GJEZc3msKzs2yYxfLuk04gwiC2+/Z702EB1I8kx/rXmyIIYsWjAPA88LCrkt3vGByz/FyXv/efst+UnRX/2aN7wZkSMrBpEPAiHpy1d+5H1K6PxKGOJZgrF7YSaEVVv7Gzl63ITKqqousyN8Uf495C8hRNavfvr9b7elv/FTps+g/ejYr72qD+hz9RUfvDR7H+MMjFBiO8qlMi1yhJCQvC1jtbfNk0sfXxzRqVqerwqhqfC2uebLV13BOXJt5Pd70unnvAbh7q7bb/q/7DUEi0cefmhWawLWgeMmEgc+9RswaDBeKOFOImPyC7pHSIQx+/svv/vV/+SPzT4nh8Ujcx+a9UpyeLSXVQdpL8MuRloMnxg9MZwfGxVhCoMthlwMpRheMbDjgYFAiWEdTwNyUlwU9fioiAR42+DZcFpUEguTkJs9kTWiIyxkQwHpzXmJA1l8etMcgzjGYgy7BWnTvIa0dQWGYM5jdGZ/IB5QMPwjiCCYZHMTYNBW2CiNkRUxZOxmTIkW3C/vBoW6Yi16q18MOZdvJJZnCPdjhKdiVGbejMG6+UxfGMTxcoEp/fBzhpChnC/w198ecMCorTBEfObZsDYJAxI5ECT0Rj9igsQOGeZluJeoAZfsWhQCin6Ul4FxZCjHC4T2StwuDw2FlJIHSPY8z5/1yIDPnqJPxAjx1FoZn2vMl9BijLUlVY3vmcprilPdMxobJsyPdbwgXBwL2kFhbsxD4bb0Wc8HMYFzPBfWx36if54Le429f25UuPLzoPwXPFcKz45nxPzl9YMwwx7gmZFYW3uW/vVvHPNCHIIL+4JrS3Pjk1sK0QIuhKdkPjwLBBIYcK+8XCxa5B6EDyZgAiZgAiZgAibQmQhYsOhMT9trNQET6NAExk+eNgOj+OwH/h97ZwJuY/X98c3lGlIKoSjzPI+hlIooSSXNVDRIaaC5aERJChGRscwUGRIyZco8z+41X/M83um/Pqez/N97nOsOhl/ctZ9nP+973neP373PuazvXut7tkE5oYk98MiTz+BJMLBn12+84Wy03jufdegMqfF+i6ZPEqZHn7d49+N23PMMY2mwfjCQD+nX83v0D26pfmfNhMaS1Pd4LDDmMcN+6RdYlzkRkmj/3j0qWusgXzipjjhxfH1hMG/Vpl0nwvt889mHrbQcugkvt/zwUz3hvnrFkjhzph6n7zesXc2p1Dip/mNPP0ffPJSQTGcZ/avecfc9Myb/MRZiAkKk28BRE5q1fP+T7l9/0Xr0sJ/7JhWXYOXxkEiuKDOGd0JBebVA6APvgzoPNnyCcE7ekE7nGm8pETvhfZnylav2+f6b9hHbt2HgOpMKisYHhMa6VcvPEn9HMP2G3DflWfTP7JkXApPANrZv3RyGePV1WbOpZoGDpELUHeIKDG4UNiWw3kNPPPM8e23u39N8HkWaSkuYqPhIRLRMKMc+mzJ+NILOQRNhxtBpmTTutxFoZAQWUu2aYB5OFwOjy6RNNUjrqX+ICgzznKTHkKqC2BhiNfwTZTHgYoylLHH8MdBiLMXQyntIUE76Y3Rm31IWDwyMrBhX0bTgZDntUw/jKm3yjKzGcy+M3lP2GHr/NcBHHYl0GfLgsUH77EeMtfz+MhbCNTGGepIhLuhXQ+7QhobOUeO+15hO38xbDe5q+Oc55ZQUUKJDPQl0zN7T/ZT3Gu7pW8kOjNkY6Bk7YX/whuM9gueEdcPoHi5ZvRu40p6SJ1zVm4F7sANj+lPPCh2zEha67rRDBnPvmDT8ls5F/68DsUD/GO7ph3sIErBmzenXS87oeLQf2lOtB+4x0vNdpR3myR5gv0AOePFk3JAHeHCw37jyOauLPpTGpU4X4w7OpF32hIYUo132zDmT/IRq2CvdX9RnLBqiK8w/R+bOc/YMJAHhDFUjg34h8+gTjwsy5ZVAAxeyhgpjv0ICQnyw/tRjb0JOUA9x9RmSIT/IYMKVvc33kLmqFw3P+A6xhhrmjDbpSwkLubVkCBgChoAhYAgYAoaAIZDSEDDCIqWtuM3XEDAELlsEMIwyeNEYmJeUSRCep1mrDz7Fu8Ir5KttcLr8jlr3PTC0X69uCPvqc8IX4YUwefxvIzBabwjiVaBlIUI4Hd6k+ZtnvDOSMsZzlUXjYdP6NasI5RNYDpIk8JS+PCtPOU69x9fui2+81wbD+HdtW7/jPRnf6MVXW2Isnz5p3BjqblizKo4nRX7R08DQLloIcUSpIZIII6UhhQI9MzhhD5lBKCkEqH+btnAN4YUQEO/VpcMXFwIrxoDhe6lHfDwp7aJvslGEOQJDYFW69fa72EN//j5qWGLbKyn6FZTdLULsA37s+k1gvcLFSpbmWTDCAp0I3i1dcHHEpbdt3uQL+6ReNGhHVK9Z535II4iqXTu2b0V03jtmvguImQ/r37u7V7+DNUUzJL4wTQWKFCMckRsqhF4wXRDto9oddxOuyE2KB+Mqt9/JKX93sbxOEruu/8FyGIYxbGKgxfiM9wEGUr6/f0nmFDeGVX7XpkoeJflXyRhQ75PMPsVQShnagTjgBDzGXby2uNffW9aSMvTDKXgyBlqMsPw26el+NfDLozNJje0YalWzIcodFSePk9sgRDB+Y0TWUEYYhWkPYz6GY/rC0K0hf3imIYq8BnXvv+u1HyUbGAz3zFfJDPXA0PF5PS284/d6ZSgxw3ueY+zXU/FqFGecEBgVJeOlotodamBXjFQEXD02WDdw57mXNNEwW/pMyQza4VQ+p/eZE94fgWQHBnAwVm8KQrexhngLsG4Yx+mXMuwf5ufVrfCe8FcSQ7GH+GHvqLi4CkhTR9eFew2tBC6EHKNeZgkFtccdXxPjYk9peyo47iWYpOg5E3UZM2Mgs7chGFhnMuugYZpU/Fx1OsAN8l1JGyWzIGFULJ05K060w3PCWml4KNZuqGQ8w5QIZP/yvcgrmT1AeX53GRckNVf+PmtYMfYN/YAP3yklfeTWkiFgCBgChoAhYAgYAoZASkTACIuUuOo2Z0PAELgsEcCQi1YDRu+kTKD1V11+JJxMx0/efSNYSJrmb330GUbq3l2/bqvt4m3xzqcdOvu0GP760xcCJ2z9WkI7BE14DQzr36t75dtq3F3Ib4xOyhjjKwtRcoOcdg/WNwZn5rVi8fw4BE6REqXKYhyOT2uBk/WE31k8f87f0yeN9xETJEiFJq+0ep/nO8UjgDY4Ge8dW66b8hLqxAVqLzz4eKMm10rDiJLjjbImgCwpU7HKrdRr2uKtD2rUrlv/p+87trv/1tIFpk4c+9uFwIk2SparUDlDxoxXLU+GIDv1y1S8pZpoX8wKHM8tsqY8U62SxIwXwW3K/dCxbZtgHgOFi5f0hUqSKGNneVhAzBF6LNi7xPSdUBmIO8ooYVGnfsMn+Dxx9Aiftgvk2E15C8QJGdX01bc+IBQTxIO3fTDjczDcIJDyCdnGfpjw2/BB5xoXoaMgQoJ55hCGSgXBg71PaL5X+Hs9yY7RVnUEMJRi8MRQy6l3jK14W01gy0nOK5n9h4GbOhhO+7OMLL9kNAi4n+4vjwEVAzZ9QGhQHgIEUW4IEfrAAK1Gfx/kwmt6Dd0YlDFGY5hVj4LT7kRYendyC54eGJLVC0mN3ZRTjwuM6oSI0tPnqksQLISTr3vJvPOKcHux0hBLShgoUaKG8mDeDLSrXgAY6cP9n8EbsWwM2PSn/7dg/Nxrv+pV4fVAAH/eUxYM8EgijJdXL4J++axz4bMSIIoxfStuXPU988D4joFc2/T9hvv7hGwBf77HEKUQlXhXeet7CR/qMQ7Wknno/mJPMAdIJYz6cfaCfAYH3uMpAymC0X+vS3OdeKakTueij6pXI2XYI7TPnkkw+b0sVGMC8oC9wX7BkwSPDg0HBr54WNA2e5qxq6cOhJ+STJBBrCf/zsCjBzwpz96H3GB8jI3Puq9ryL2uG2Nhjnw3wJ12aQdCjmd4qEGqsB76/eE7Sh0NLaZeMhYOSkCxZAgYAoaAIWAIGAKGQEpEwAiLlLjqNmdDwBC4LBHACLxSwtYkZfDPNX/zXbwk0E1A+DiwboUqt92BlwJkw6ED+zFS+FJTMdzzHJFrDPk8I5TOufoe1KdHF4yuDz7WqElSxniusjkkNg8GW4nEo/G0zxRXke+5M+OG6ClcvHRZxhqfMPmjjV9ojh5Ir++++lwbw2vik47d+qQNTRv6Veu3WxQtWaYcHh2BxnaEj6mzc/vWMyGOCCP1wuvvtB7St0dXsFq7cvmSQGIoxw03Ymx0nT7/8K3alYrk7i6G/OQIp58Lq0rV7riL98F0NxJaDzQSbs5XoFAwTwFCkUFcrREB7YTa4T0eKoQ3wttk7Kiz9RgoU0jEWBDVDuY1AzG3evnihV5PhsT0m9gy6gUjEhoFqFOv4ZPPIHiuGiIbhbC4StTc8ZzgPcLZeCGN/KVPz0Bx99IVbqkKARJsHvkLFy0OaTFP9mdgvcCxQmxA0Bw7elRj/Z8pgvdT1mzZcyBAfnD/Pk6GW4qLgBo1MXJiHMUQilEW47qGPsKIzHeQ0+0YjcMlQ8ByIh2jLrhCaGC45bv9h2RICQyoGHYh8jAEsydon3eUxbCN0ReDLmU13JOGaZJHvoSxGKM6RmQV545xMccPu9jI/S4mGiMwotfU01BA3NMep+AxhNMHoZe+k4zhmPb0xH/giXyvoVe9EmgLQgYjM7jw+azwY/4x6Li9HhdqdMdgT9/MHxx4jvcC81dSAbLIm5Tw4ZnqT9C2kjeqPYLXA2uia0d5SA1vCCklEDS0kHpVqNHf65mh64BHF6f+GTf9Q1Qwf/oCD8bLVcXOlXjxEkJe7w764h1/G/nbRD32RyDRoeuinkAY6CmTQdb8iIs6fMSd2sHaq0YGe4M9wjjZM4lNuvcx/LNfaZN9iocgpDDrTIZc4u84pBx7HKKFv/sQeZRlf7D/IRdYC9YX4oLy4AXmYMOa8D2CnKA93kFCQEbgaTFFMiQh4aFoD+KCNYYIBjP2DmOB9PNpssifYNpkzD5iCcJPMsSfL1syBAwBQ8AQMAQMAUPAEEhZCBhhkbLW22ZrCBgClykCGMKvF6v3iiULEk1YPPV88zdee//TL4l7/1Wbd14LNnWMtTwf+UvfH/U9RMWLb77bhnj+wwf2/kGiIJXC22Dntq2cqo03YYCeO3PqpNslvM6FglmkKHyi2sKlnGWorSe6HGhXBBrZi8hp9XOFr7r/kScaQ2gwVh3n48+91AL9jc7t2ry7duWyJcx5x9Yt4YHzyHJ99hzRUVFRXnLn6RdeeVM0Ea4m9FERIUu2hm/C0BMnXSsT4cGwAb27XyzRZMIKYdQOZjxPaD003NjSIB4WEBk7t23ZfK6QRt72S5Wr5POuGDWoX6/4SIdCxUqUii9kF7oPq5YtIWzLRUnqHXNzvoKFCDcGITFm+C/9tLNNa1dzctihncL1jQ8/7wC51P+Hzl8HDqiM6H4Ew4xyRUX5netff/xOCKJzJgij7VvCfJ4fganxS6+9xbNg4bMSavdKfu81Zvq9GfRUu4biwZCMERmDqRpaOemNYRZDLCGjekmeJhnDK+UgAniHwRfjMYZYDK3qKfCvsfnf9tQAjNGbeyVHfMbWAOzRL6FNDPG0Rdt+jwQpGnNUQxFhbKYtCBbeczpeNTH4LcSwPlEyv4dqHMeArEkxUEM949BT9xiox0lmP4ZLxghNO15yJTC8lFqKuYIR46c/vBCq+sfJvNTDQcfEeBQDnmnoKeqTNGyTYoLBHwM93g/efigPEaJeGlpf11O9KpT80M/04Q3NxZpBNoEzzzGYQ5aAN7/NvGe/0A59KPHlH+6ZuagnCnuCMowVDw71GmGuXtJC56qhlthfGOQPClmVWcS2T7q945gL+LEnKEf/4BKv5o0OSq9+Lwv1MoKAgCCgPcYJMQC+PKd/QjNBzuhc6J/5sw80fBblIU6UjIFE0zWAuIaIUE8j2psrmd8vCBm+X3zPaJ/99bdkSA2+VxB/ECjUAXsN/xQjf184N8B3J9j3R4paMgQMAUPAEDAEDAFDwBBISQh4/5OTkuZtczUEDAFD4LJCoIQYVRnwqmWL4xWS1gmFhqZLJyLaXRo89dyLhKpp8cwjdYOF5aE8J8cx0GPo5jOnyr/9afBv4tEQ8Umr5j5PCQy7B/bt3RMsnFQgiPRXrUbNOngwxNdnUoCnHcqfFCu/tx6aAnhBDBSSwGsUV1HscaOG/Bysn3wFixQT2YH8v/Tu/p0a4CtVu/3OVq3bfTNzysRxPKcNcFg4d9aMwDZ4J9GKVKzUZROXC8JI9RYdCrQwEOTeNWY7hsA46RphLHgQefoUp0gveEJEGg8cEW0enpzG0b5AUFrDJXnbIISWOB3E0fI4Vx8QALyPL9wVug+Md/3qFZzijZPQFUEvg7BMyZlHYupAckkEswMQEojR7xGdjTkz/vpT6673a7UULFK8pMhbZMEL6WsJpwY+3vZla2YULY4yo8R7KVi/7E+ez542GUPxOZNE8sokwzpLo6XW/Q81ZK9TedXShL/7CfVzhb/X0+wYXjHSYlBWwzJGZZ7z3dW4+RhVNXa+ijFjQMVojJEfI7SG6MGoy/rw/VVxbv0uq56CGuGDhbFRLQrapX2MwX4B4ugYd3pXYZcmM8Zh+qQfQgapVwHGbPqnPwgYfpchR5TI0H69yxt4IIl5crK9m2T+7d9ecn3JD0rmt4nQU7QPaeD1CuBeyQFtkzKMk99mxLX5rAZ+njFujOc6fu+41HuEdiENIGAYP+sENni7sC4q5sy6QNqQ1MDOPW2Du46Je8ap2hcQ+/wO8YwE/tyz/njJ0Sb39AuWKngO7hAGtK+eHLqe3nWlP9pkDhjq8UJ4QDJETqCHh5JdjA1yhHFEu9MReVyqyBiXOlS9NVgHMCBr+/7hJ3zB0C9/0yioxAV7mfmR2DesO30wPsqw5jyHOAAPxgmpoYQL+PCbBwmh+wJsqKu6IboOSjyxXpSBoABL2oYIVBKIfaJ7iv60vpEU/oWyiyFgCBgChoAhYAgYAobAvwgYYWE7wRAwBAyBywABwvIwzIROnmN8f+vj9t8SEx+viQ4fv/u6V1TaO1W8Ngg1M/WPf3UUMCJ37jt0DF4Nzze8r4aGsRGdiJsChZgpj1FfHAuu8WpqpJLwTTEkCQ11IWDVfpW40DZffadNW7QBhvSNqymQXTQtKLM5LLjOR/Ey5RAAdcv9wuUFChcr8XXPgSMkxNPm1m+82Jh3OSSmEddgcyb8k5eIee+Ljt/vF0M2REee/AWJ4e12iQBG4NyF4/CF+pHqGdBnuBDYeNuoesfd94SkSZNm3t/TCMWR5EQYpmXnEOvGOB/YKF4B7B+Eur3vINciRAMkUP9Dy6jGyQaJgRTY5o033ZyXZ14vEQgO2U5RwXBN8kT9FTatW7MKEe2s12fP+dvQgX28+5X5sIX5zlWsWr0GBMbQ/r0w9MZJxUuXrwjm8eGGlgreHIkZ92lhAwMxhrh5+5Mvv0MInHebNsSvIZNcHK7AenoKnCvGUTVqawgkDdmEwR1jrhrKKa8eEtRTYoLvqobK45k3LJCGC9JroG6FF14M8RiH8ZJQLwCMvpHu4KwjLlvdzBIiKItLHcL4VNeBK/9OZwzqOUFoKH5nMCSrV4Ma0nWuXoM57/D44kT9r2LU5rS7E8M2Bmp+CwmRRQIH/T+BkgBquGfcGLp1nup5ghcUvwu0QVne44XHHDFW+7ryX9WLA4wZN0nDRvGOcpy850pbEKSEcYLgCNSQ8Fc/Q1Zo34orc+HvpfatAuPU47ed5xjKmRNeF+DLnLnnneKgxE2gHoXuFQgnvGuYfwXJ/O2hLbD17g0lUdRb5rSLiUol2iUx7vjmSHd8LeNgnoo7YwNz9kySkp+0oG/GAdbqYQEGPGeO7CvW0HcYwN8378GR7wUkDGUhV9iPeEmwV3X8qn+hbVLWS3iwJyhDP7SlHjLqZUN5MNF05vvjeWa3hoAhYAgYAoaAIWAIGAIpHAELCZXCN4BN3xAwBC4PBDCeEnKJ0+CBI0aYusY9det/P2Dk+B+Hjv0r0zWZM7/1UqNHvnjv9ZfiIytoA4Mz14PiPnGNHCXvOeT3ycVLl6vYpmXz59Sgz3tx2EgXLLb+B+06de/366RZ6BVQDm+Dh5985gWEgSETLgSyojewiRBMBYsVR4zVlwjBxKn3If1+/F49Q/SdSA/4TuPiERKsfw0xxZyLlChdtvfw8dOIQ9Hi2Yb3K0HDfKkrGstn6Qmc9JANCHfffe8DD3/z2QetmK/Yl31Gut07d5xFWCipU1DCHd8AK6oAACAASURBVHnHVa5S1ds+/7ZnfzwzzgevJ5o084X8mjV1EnH4k5TYP4Rx8q65t4Ft4WEbCXWFroM+Z60HjJ4yp9XH7Tt5y6I3Uqxk2fKEIYtvEJBpvFMtCW+5EGEA+JwhYyZf/HbCQw3+4+9FOr8kTewchQkZBgmWTUg3Qld5i0IQbBddCkKHoceBpgl7MLC58pWrVYd8Cka8UJa1RosjMWOGJKlS/c5aeEdRHiLki84/DiAM3D+zphO6yEV4dFMS02YKLqMGUBWIxujKdxnDK2QERlRICDKGYX3GaXBOy0MGYIymHIZfjLjqQUCb5Gj52SBrrH3i2aiBPBj0agTGWK/6ArR72h2eG+WOrj3mYo7gWQGxQDgo3zaQzL/T1Wivhvc88uwpyRiG4wvur8+ZB55MtHGjEBUhkuvJ/XuSEZqmD8YDwcwYz2gIyL16pKhYtZ76h2gAJ+rhraB6C+AMYYFnGt4iSvB4PSNoS0/Y06eGoFJ9BOZYQnJZyRCaYKRJ11Xnpp8ZF4Z5bZc5j/HPBcO5huEKDJ3FPOgHLxHIgWBYKpnCGJQ44arC1XjKgCNEAH8Hvd4g1NGwVFzZV5AwUS7mhAhtHwtxx5bzd5LMPMHGG16L9Uhy8ms/KPnAvqcd9rnqs7A2fBf4twT3hI/Ci4Ir3i2UY0wapkz3AfsTPEmsHX2wxpTlu0R52qVNDTem3iLqAeMrL2PUfUY75/reJHn+VsEQMAQMAUPAEDAEDAFD4MpAwDwsrox1tFkYAobAFYYAJ97f+OCzr0YP/bkvBlEhEiqsWbF0MTH3xakhMyQBwsVF5ZQ4XhUQDpzm/qrN26+N/Llvz8QQBoR9IiwSItQPP/HsC7TZSYzvE8eMGOKFExFnjKkvvfn+xz2/bf+pvkPj4q469R7qPWz8tPBN69dyGh3j99vNGje8UMuBl8PfU/8cX/Pe+g2atnjrA8SrH3m6aTMMvN06fP5RYD8H/cLhhMMi7E+V6nfVerRx05ffafbMo4v+mT1zT0SEj/D5uMP3vbNky5ZdImjENn/qwdrhG9YRX9uXNm9av466Dz3euOmC2TOmzpj8x1h9J24DGzDWd/zx55HM/ffhg/pPnzQe45jDu4Sr6CafZWiaPH70yHc//7rre5937NqjU7tPCBF1f4MnGoEr2gRHpL/kYsb6YzzHS+CL73oOwLtk+5bNYbsjdmxHpFkiVfmEdTmln0FiWmWQsFbXSZyntELM9O3W6ctcN+fJxzsIl0HjZy7s0antx945jxkxqP9r733SvlOvQb8O6vND58zCdL3c6sNPESBv98Gbzb3jzlugcNEMEt9o9YolxDcPmtAH4UUwTxP2MHsS/RU8ViCFjh0R/YgeZ+tHJBcv6q1a/q9GxjRZO7xBAtvaK4LrN+XNX3CKrFt85EvBosVKHjq4f/+zL7/xTg0Rxm5c/25i+vsSBBTfySUL5s1OzDjHjhg04F3ZG136DRtLWK97H2z4JKTchN+GD1q9bPFCdGFEv1vD6SSmyRRXJkCYVyO+6cl+DZ+kuCgBpafo+e6qcdobZojyXm+x5BpXi0k74ZIhGyAaMOzS1gkXfSLKpRGO4tDsdC7rfTo+fg8oB3HHv9VZexXrZjxqCNbQRcHGxTNO0VeXjLG8pv8zxvX8kjG88572aQcDvobBAh/q8AwCBeM0xARXjNZghcaLEio8Q3+C3xqITYzWGO+9XhuUpS01XqvnAuQH9ajDOwzfCJDzO8r8vboYuk66RswRskIN5xjKEX7mu8g9Y/ISLj4tIf84uAbDjTFoOCvGqMSKtzzvEfGGsPCOE/xYK+//rxgrYwBLxpnVnVwf6k5t3+92j1SCinWgLvjwLFwyeybZya9rQf1o+TIoUaTeJBrGjPdeDxYlbVQrRPHRMirSznPV7dA2tKyGuPK2yzsv+aNC2sn9PiUbF6toCBgChoAhYAgYAoaAIWAIGAKGgCFgCBgCyUSAk91d+48YN2/D7hOLtx6ODZZnr4042mfUxJmIAqtuQFK7a/Hux+3+Xr3j8JiZS9ZzojxYfUSXeT94wsw4Rmg8E9797Osui7Ycipkftu90z8FjJnMiPqljSKg8YZumLg3boxj0/23ybMJRxVfv004/9PXixbjU+4GQTt0GjpowZ92uY7SD7kOwdvBY+Xv19kOt2sT1IODE+7Tlm/fR/je9fhnlDVWFgZvnHSXEVLA2G73YopV3XBPmrdryTLPX39ZT9QnhEN/72vUaPDZ3/a7jC8L2R8a3V4I9HzDmr7mc5Cf00LyNe05SptvPv/6hWGl/kBk/jZgw3dvGxPlrtt16Z617A8eExwnl6tR/5In4xgs+CzcfjEavIliZlq3bdtS+IFBy58lXILnYxFcPQhC84lv/Lv2Gj/1ryabd5/J8QdCecU5fsWV/4Hyr3127Lu0n1nOGPcB3WefNd+qTb7r3YX/h9cTzBxo+9eyFxsHa84VHShUkXzBoYie7qyV/J3mK5HWSV0teJHmz5NmS58TOKTkudu+fq2QcAyXPlwxxt0PyMcmbJB+XfFDyFskQzScln44nn5LnkZK5Hpa8WXK4v50xcp0neYPkvZIP+N/T1n5/u/TJ/Wp/X2v87Wz3j2unXMMkL/WPiz4YK+Pj+Vj/Z8ZJu7THWLhnHkck7/aXYQzMlfFMkLzHPy7q8o6xU5/5Bs6ZOdKmzveo3I+Q3ELyT/62tvnrefvXOvpMr972FFt9pn1rWeawyz8X7nmvmAeuC3NlDqwBeVDs7t+Wxi66Z7Jv7f/dA+wF9gR7gz3CXmHPnPFqu2AbMpENyTjj+24E+77E5+mTyN6smCFgCBgChoAhYAgYAoaAIRAXAfsHpu0IQ8AQMAT+wwikkWPV9z7U8MnPOvXo10uEnReJEDReB4QvEtmFsAulFZEYCDBuBwuNQ6ggMW7Eii72GTHqxLSXlDIY1ctUvKUaoZ4SIzyOoDIhr/A0CBZGKzF9pw4JCYkVLQPm5i0fn3YDZdp06NqL8Y34uU/PYH1gfM9fqEgxie61fZ2ITl+o9YM8Ypx4uEAwpBc3hzNX0c3A8M179DfwANm/Z/cuvEh0jOhKMNf4whsR6okT/zluzHUTIa8WzZs9MyoqUk/hnpkq3hWIVa9cumg+OhDBMMDzAC+Vcwlrs954FOAhkpi1Sk4ZNFsk6lfQsCsQUyKbEYVAd3xtg2/ZilVuJQRaoLcIuhsFihQrgZB7YscGxqUrVK4qy5VRHJZW4SGjdfE4Gf/rsF/iC3WW2D6s3KVHQIzOnMIn9BCizLUkcwJ/tWTIXbwJ8JbY4/K8t9/l/+Iq0bHAM4HyqhuhIZX0dDxXTveT+G1SUWc+U1ZPsus7fpfpg9P7YZLxSOCeK14TnPonFJNmPI7wbFBRZE7M4zGAFwUGdPUUwCuAPqjPnNQThd8FdG3wENB2vDoQqqFAqCoIYz5v9JdV4WlCNBGCCDFrQi7Rl3pVeE/ue/vEiwCx7QWSEdymbcJDQYx6PQXk4xmNCfXY8P5/SDHUMdOuekxo3yq8zrzVy4V2SSo4ruvCepDxWJkpWiW53IFJUW7JveCpYt9c0e0AM/CbJBnPvSWpavrCOVkyBAwBQ8AQMAQMAUPAEDAEUhQCRlikqOW2yRoChsDliABG7o/af9eDUEvCVWgM6ctxKjZmQ8AQMARSHAJCWjwik0bw+R7JeIehF4B4NonQRdEuR8NjrtjAvS4knQpDo/WCoVxDNUEwQFZgIIdc4J2GtKKdwFBW+g7CAmJOxakhKzTME/V4jsEcwzjPNawR4X8gDSBQMMJDGnCP4Z05qFA0/5dQ0kKN8xCNqguh4Ye8YZzog79leO1RbrTkpv550R5zmyb5VsloA/FZCQT9v4v3M6QKc5zobw/C5EHPOL0khIqTy+sz+Hlx5Lkm5q06FN42IEoUfyUmeK/lvQQJZBHrxTpvdzGnNroF1dK5I4vQvGAtEesmQc6w9mD+p+StQlYE9dbzDtDuDQFDwBAwBAwBQ8AQMAQMgSsRARPdvhJX1eZkCBgCVxQCiBM3e7J+LSMrrqhltckYAoZAykGAk/4YtJdKxusA7woM7JACaFVkc7uGx7g9wyEC8L5A6wJyAjIBIzjlwiVj4MYrguT1plAkvYZ3NezjFZFNsupRMJbN/jb5fwBeRBAIiFxDWmifGNmpg+6DajXwDtJCdR6UNKAsbaneBgSIimCrBoVXw4A5QFSUl4zhHsKDZ5ArKuJNKDg+g4N6NnjJAxXd1vHyGeLiZsmQBODm9ezQuqpPIa/PYKhYBWoqKBmhGgzUZayQCupB5u1Hx6li4eiOoI8EthBOJ9yWDmmFrID8YU1YexV9Z0+wN9gjtMM6WTIEDAFDwBAwBAwBQ8AQMARSJAJGWKTIZbdJGwKGgCFgCBgChoAhYAhcIgQIfzRV8k+SCVs0XzKeA5y6x6shXPIhd3CGilv/5X8OEYARHiM5hm28GjREE0Z0DUfkNczrlLxGeIzllOXf/RAA9I3INcQFzzHwY+jnPWVpm7Hsk4zRneeEa9LwVIzD6+lAn2rUV2KAqwpO6z3l1NBP+xjuIURekoznBmHQIADwkMCgz9gYr7avhIASMxr2irpz/XXw3EBfBzJAx6LkRrArbQd6behcAokSsIdQwSuCtvmsY+Oq5AxlwJQyeE1QHiy7uI1tuKqwNmvPHmA92BPsDfYIe4U9Y8kQMAQMAUPAEDAEDAFDwBBIkQgYYZEil90mbQgYAoaAIWAIGAKGgCFwiRDAsI0nA8Z/Tttzkh7dBjwS8LTIJ7mg2z99vYuJwuiNER8yAcM2xnPIAspgQMcYrl4HapDXaaiHgNfTQk/w42mBYRwiAKM+/aBXAWmAZwVZNR1onzEzDsgJjO8kxqteFN6+vGGflERQcoN+eE8YJX2nIZVoi3d4cEAwMF/CQ0GmqMFeiQf613YCiQQIgSKSCbPFfJgrOHk9JPxT8F20voaHUoJGPUx07JRlrF6iBjzVW0Q9SyhHG+ptwZxVI2SH3OORscateHKGf44F5cp6svZgoBoe7A32CHtFyRDvuO3eEDAEDAFDwBAwBAwBQ8AQSBEIGGGRIpbZJmkIGAKGgCFgCBgChoAh8D9CACP0XtEkwHC9QTJi25ysV00IjPKn3Yl1Rdz2HqvkHnFswiphfMc4jiEf4kA9JbxhjZiSEgbqaaHEgxr4Ocmv+hIaBopwSzkkYzTHKI+xXsWkeacEB2PA+E/GWA/Z4iUg1GNCx8HVKzitnxkb/dAHdQh5RD+UpW1IGTLkBeGRqvr70v40BJZXC0OJB66IaxNmCkFy5sWcNSyVelAwFk3MRXGkHMQBcyYpIUE9cFfsuIKHtqflNASU19OFd8yV8YPtBLdrcEW5IqgOGcGa4xnCHmAvsCfYG+wRNECOiPaJJUPAEDAEDAFDwBAwBAwBQyBFImCERYpcdpu0IWAIGAKGgCFgCBgChsClQECICjWc090ov4G6klz5dzgG68WSOWUf69a1wOiNwRpjN0QHRm0lDDRUESf5MYir54MSBJAAGMMJrQQ5oLoSGOZVEBqvCoz7GOfRysCLghP9lNf28MLAy4GwTTzHuM47rupJoGGeNAySvDoj/M29Gu/VEwOCQAkAFQ6HWKB9DVeFpgWZsTJ35uP15PCSFartwXx1nBA6EBV4PqiXiZI3Xn0K7ilLPSV7lLTwiol7w2p5vVbUM4P3OhfmrN4YrBntK7FDiK+x/rnRDmvNmrP2jI+9AGkxSvaKrx32jP/e98CSIWAIGAKGgCFgCBgChoAhkJIQMMIiJa22zdUQMAQMAUPAEDAEDAFD4JIjIMZnDOxOrhi1Cc20TjLhgiAPykmGDOA0fhG3qTUhmSAWwiVriCMNp0Q7EBh8po4SG5zyh4SgfcS71SOB+iT9N39Jf/94cGDsx7jOqX7IC/UmYBy0QXuQHzzHA0FDIKlngnpX8M7rXQARoH3qc/Wq4DP90gZXCAbqq/EeEW6eMw/GSJ9eTwolHqjP3Ji/kgxekoY2GYeXdGCelNH2FVPGqu0G6l4o0eN9Tt/alxI4ECzaF0QM3iMIbqPHkcZNSYVnBWGrwJZ1Y81Ze/YAe+Fa/95gj/j2iiVDwBAwBAwBQ8AQMAQMAUMgpSJghEVKXXmbtyFgCBgChoAhYAgYAobA/wKBcX6jNYLMnLQnDBSGe4zeN7iwLxDAniIZw7d6R/BOvQEwaKNxoUZzykBYqOGeOalYtxriVX8CozqECeLP1MOoTxgliAue0Qdt8Zy66ELQnxrmCW/kDaVEP+r5Qb+0j3eBemzgqYFRnrBWeFls9Y+dPqjHM/V0YPwQFMxfwzMpCaDeC/Sh/XCF6KA++EHk0IZ6tKg2BaQGHiJ4k+DJQMgt1RRR0kVxpo56U6hHiNfLgz6V6FBMKAcJQVgn2ibMFlfIHkgSNEPwnSBkFevIWFlz1p49QF32hCVDwBAwBAwBQ8AQMAQMAUPAEBAEjLCwbWAIGAKGgCFgCBgChoAhYAhcOgSmSVcL/f8Ox5sCYzpGfkgDjNl3ualpIQnIGL8xfHMynwTxgGcBQtMYzKmLkV71ITDOQxBgGKdNknoocE/7lEf4mbqUhaigb+pg9Md4zzvVaOD/CxAJeAxAPOA9oG1q6CPa1lBVjAEig7JcaZN3eI3gTUB9FahmLkq0aH98Zr6QEdTnuYp3e+dCnyTa1+fqncCYGRuf50sO949ntX8c/8gV7wevvgXYKmGhVyWJ6Mfr6cE981DyhnFC/OCpslwya4aXymG35D6Ikrskg72GiwJf1p5xshem+WZiyRAwBAwBQ8AQMAQMAUPAEDAEjLCwPWAIGAKGgCFgCBgChoAhYAhcKgQk5I+SARi2IR7yS8boXloypEGUi4m6ykWfXCT3EBYY7kkaTgljOp4KSnSg9YDh3yvODcGAdwPJq9+gBnr648R/AcmQA2QM6xjUMfJjvIc4UCO9ej4QxkjJE21bwyV5NSY0VBUGfdrQ9pkvwtq0r6SFenColoXqQtCekhmBXg7+qZ3BhRutryQDhAD32t8vcv+ZZDwy8GrQ0E7alnpOBAp78z4wTBPt0oa+w3MDMmaYZNYF75hVLvp4WrdvAt4kqsvBGoM9aw4W7IEY/57wzsnuDQFDwBAwBAwBQ8AQMAQMgRSLgHlYpNilt4kbAoaAIWAIGAKGgCFgCPyPEBgj/RJeCYM8ZAMZAgEjNobw0m5rp3lyXSoZ7wmM7youzZA5zU84JU75Y/znhD9tkQmnBGGghnvqa/J6FKz11yU8EfczJKvHBPoR6mVAXYz7tO31KOC5V6OCz9TRcaBHQXnGiHcBn/FAgLxgTGT1ntCwUnxWTwsN6aTP6Ms7Fy8Ro215BbEhWfgMOQD5Q8gmRL0hZSBzeK4hpHQu2rd+1vmBsYpo6zwhJsIl402RRTLEEtoUlIM8inERAyAyIClYU9aWNdb1pm/2AHvBkiFgCBgChoAhYAgYAoaAIWAI+BEwwsK2giFgCBgChoAhYAgYAoaAIXAJEZAT9egXYMzH2I1BHy8JSAkNpxTutv+Q3cXGYHSnDM+VhEB/AWM5xnQM3kpoQASokR8DO1oQkBzck9TAr7oNEAgY2atK5tQ/Rnz6Uw8K9ZxQLwuM7uoNoVoXKjbNeCjPlUQd7tHLgPzgczbJECI804RhX/UplAxRkoCrjoF3jD++uagnB+W9uh2KXwV5fqvkMpLzSUYEW8XLPcM5I1auY1CdCtUL0fbBYaNkvCeYJ/eQE7pGu1xM9FG35mVIiXDJqinCGrPWrDnrGuLfC94x2L0hYAgYAoaAIWAIGAKGgCGQohEwwiJFL79N3hAwBAwBQ+BCIJD75rz5a9dr8NiFaCult5H52uuypJKU0nGw+acIBEbJLDF4L5GMUV91J/BGKOpO773RHZyClwWGdZIaz/UzxnG8LCAaMOTjQYDAs5aFrMBQrsZ3nisJoGXwNtgrGUP+3f6+lBxQYsPryUA9NC8YN8QJhAP90C5XNehjmCfEFHXxKFAPBa6QFhAJGP0pr94R/qGfGT83gf9XiW8u2obOj7HreCBKeF9CMp4QaEug4YEnCnPwEjnqleINQcWYFRMlYtbLM9aL+mBO++CyWTJrstvtHsza5ZVcVDJryrypw1qz5mDIHrBkCBgChoAhYAgYAoaAIWAIGAIeBIywsO1gCBgChoAhcEkQ+LD9dz1atWnf6ZJ0dok7+bhjt58+aP/tD5e42yuuuzRp0qYdO3v5ppat231zxU3OJmQIBCAgJ+uny6MFktVoj2EfIz4n8LO7mJO5XHiH0i76BELRGLcxeKtoNt4OnN6HGMAIjkEdA3xmyZABZOpwxYCOFgZt4w2AMR4ig3vCFGG8x9OipGT1fvCGg8JIr2GZ1AsEDwEM9PRJO4xHPSWYD+OkrIZcUg8IJUHUk4OrkgEa8kq1JORVHFFsHQf9UEav3AcSMXymb/UEWebHgGeIh9MXcwBzr0eH9ul9xr1qWIAlBM+PklVjBAzwVoGIgERK7U7u2OZWNgLPm/zvWFPaoD/11ljg3wP0ackQMAQMAUPAEDAEDAFDwBAwBPwIGGFhW8EQMAQMAUPgkiBQ8776Da7PmZO461dUuirT1deUq1T1tuWL5s+9oib2P5hM3gKFigicmSNPn8LoZ8kQSAkIzJRJQh5g/OYKycD1X1Ho/ZOLuWNL+Pc6xm4M7LxXnQjwwSBOCCfIAQzrhCUiTBReARjHldCA1OCeZ3y/IBmoB+lAoryKSKvxX0M0KSGA8Z9xREhW4WrKUg9PA96rbgSeFzzX8arngnpP0Q5ZSQ68FBgfhECgwLY3PBPtMH7K6Pj8Uziji+HVuaAMREIdyZAKeDvgSeINN6X1eUZ5rwi4htjiOaQDmiI/ScYjBQwgeiBBwARSiPXY7/aPR3S7ur89cPCura41a2/JEDAEDAFDwBAwBAwBQ8AQMAQCEDDCwraEIWAIGAKGwEVHIG/BwkWvzZI1W9j6dZwUvqLSbXfVvi8kTZo0q5Yt4qS0pfNAoFCxEojTuhVLFv5zHs1YVUPgskFATtivk8ESlol/k2OMD5eM0R/jPYTCEbfhg3QuOpJT/V5PBAzglMcYfp1kDOYY1/mMEV3bw3hPO5ThPe2qeDTkBeGReI4YNHWVnADDQJIBUgMCAlIBYgRPBW1PQz1pffXs4EpSLxL/Rx9xgsF/h+RwyfxtILSV15vDG/5JPSWUFIFw8Ya7CtS70LqQCSQIFfCDNOcZHiCKs2Kp3h989npwQGAwNrw0GGch/7hLyZUwXEpG/Osdc2rbXLfuTTxXIImUTKIv5qmi4Lv8a+8fnl0MAUPAEDAEDAFDwBAwBAwBQ0ARMMLC9oIhYAgYAobARUegTPnKiLq6NSuWIjR7RaX7GzzeiAmtXLrYCIvzXNnCxUtxatmtWr544Xk2ZdUNgcsJgcEyWLwntkhGAwHvBDQSMHavcwemnXDHV4eIiDOeBRAQKhYNwYA3BcZ5hKQhDwgJtUkyZTGSQ1RgJMdYTz28BDCkQzpo2CQ0Hjb4AcNQr4Z7JRnU4wGDPAQLhAieBNTTUFBe7QeICJKSGNzTl3pX8JkyzBPiYqtk+oAUgEwg9JWXOFHPBw3fBFaqH8F8eK9eFeqNQh8a9oqx5fKXgagggQ910dmgT+1D+1VChLJKXhD6ibJ3SQZvfvN5BmkB7plcTNRhF/FzVRd9lDmAFWvIWjJX1pY1ZvysuSVDwBAwBAwBQ8AQMAQMAUPAEAiCgBEWti0MAUPAEDAELjoCJctVvIVOVi27soz62XPemKvq7Xfdw9y2bQ7beNGBvMI7KFqyTLn9e/fsjti+DaOeJUMgRSAgJ+0xZKsoczW5x7iO5wNG+eKSs7tdg4+72FiM8hj1MbZjYMeAz7/lISowgvMML4CbJUMuYLCnDm2rdwYEBmQBBnXeqbYCngfUUWJBCQD9rORFeSkDUQH5TFuElMKgT0gn1Xlg3Or9Ibe+e68mBuOHzMBrJEwypAcZEoQ2lPzgvZdAYT7UQ2dDQ1hRhvaYP+QNc6OO1wMDzJg/9WgDIgfsCNtEOzpHJVpoSz1HmBfzIdMPpA9j5DcKnNVbA2+TTe50xHYX9iXPCD/F2lGPtWRNWVufDol/zeXWkiFgCBgChoAhYAgYAoaAIWAIBCJghIXtCUPAEDAEDIGLjkCJMuUr7tm1cwf5ond2CTt47JkXXiEcFF1G7NjGKWFL54FA0RKly11ppNZ5wGFVUxYCrfgZkYy+AR4SGNcxrEMOiDrCnFTuZNhe8bLAIwCDOsZ1wjNhGJ8lWU/xc9qf9xjNlaSgBYzyGO4x5Ou//ylDP7SFAR7yAc8LJQyoR1n1jMDYjsGeOhj7yYyPMgh30x7GfL2qHgXjYKwapol5KbEAMQIRQJ8Y9vFawNsDwkD71zEooUA7vIeYyOJvC68PvB1oDwyYD3gSbotxMiayinyrCDh9aDgp32+5JNqC0KA8zyAtaId5V5QMCVFAsuqKgH1B8aoIdyuf2OaiDzEmEtjQH/VYU9aWMbHWlgwBQ8AQMAQMAUPAEDAEDAFDIB4EjLCwrWEIGAKGgCFwURFImzY0tGDR4qWuNF2C9BkyZGzw1HMvAt6xo0cOky8qkFd44zlz5b4ZnRPTArnCF9qmFxQBOXHPyX+IhxKSISHwlNCT/pHu5PY0LmrfKXdiQ6yQFvz7HYM7BnXqYWCnLMZwvClUuJt3quEAIYDxHWO7ClbTDiQAVwz0KjbNb5lqSTBeDQnFM/UwUA8O+oWsxahPfxAF9EOIJK7UZTwadon2VHsCgoF+8ayA8ICEQBuD55AnzEvDMamouOpw4JHBePSqmh2QKtou7+iXMXuThn1SIkTFxCFOIHUgJyjDXPBAgXjR8FcaTgvih7YZY1YJBTXZbf22sjv4N2PiGbiq5wtryZqytrP8ax0wJPtoCBgChoAhYAgYvFluowAAIABJREFUAoaAIWAIGAKKgJ4kMkQMAUPAEDAEDIGLgkDBosVKQlpcaYRFw6ebNst09TWZVy9fuig0XagKy14UDFNCo8VLlavAPM3DIiWsts0xHgRGyfNykhHARtgZUgLDd7QLyZDWndqRzaXJnMHFiF09Nl2UCwmBNMCjoLpkRKUhDTDOo5sASQBpQBn1tMCDYbzkPJIxyEMcUJb+eIcRnqREAQZ9JSu8OhaUQcNBQ03hwYDRn/7xAGEs9M1YIAFUzFuJAgz9EAF5JRNWCSM/XhVrJZeW7Aub5G+TvpSYgABgPmT+DwNZAjnBcw3ZdL3cq4cHYa70/zpgEJh0PFyZq3qcQFBs9/fPnMIl3y4ZvMAOYgjMmFs2IZBC3JGFZd3GNowHfQvV1KBv8GUtaQ8yhDW2ZAgYAoaAIWAIGAKGgCFgCBgC50DAPCxsexgChoAhYAhcVASKlCiDAc6tWLxg3kXt6BI2nk7cK555+fW3x/069Ofo6Kgo01w4f/CLlS7rIyxWLFk0//xbsxYMgcsPATl5j6F8hGS8DPBywIiPwTvEHV0e6U5s3OaOLDrmoo+kcrHREBUQpfxbHqJhuWRCIalgtXpfqN4FxnOM9hjeCU/EqX8IAoz1eBRQV70XNCRUoFA2oPIOkgBCAQM+/TFutCQgKPBKWEJB/3MlRiBQSHyGhEH/Au0O5kk7kAt4WhA2kPeQHEqY8J5+mYu2gYg1XgsQFepxQuglJU5UX0LnEGwuqqvh7Qcc8O6AcJkiGYyr+vsGU8gRxsj4KbNEQnVtcSsegsSgf7DUcFysHWvIHFnTEf419k/DLoaAIWAIGAKGgCFgCBgChoAhEAwBIyxsXxgChoAhcBkikLdAoSLV765d93IYetGSpcvFSlq5dBGxya+I9Gjj55tfe13WbL06d/jiBgllZPoV57+sJcpUqLRr5/Zt+/bswvBnyRBIkQiIQXuuTBzyYYVkTvdDBkA0ZHIHZmZ2qUKjXdT+WBd7OMRFncQIjiEew3kVyWgnYLDHQI7BnxP/GPkhNFSsG+8HvCPy+5/zeaVkjPB4AUCEqCHfK7yt66FECAQIng5KmDBG+pojmfBO6iWB8R8CAjJD/9+hpAXl8OagLoLZeHmUkYyXBonyzIFxQBRAejC3Gf4rdQgpBTHAuLR9iAM+K/GiYaX8zZ658Jz2uEK4QIwwVjLEBdhoyCwICsoomUKfp92JrYdc+BcH3cmdhIwCZ4S2/yWZ/l071pC1XO5f28Ax2GdDwBAwBAwBQ8AQMAQMAUPAEAhAwAgL2xKGgCFgCFxmCOQvVLT40D9nL+3Sb/jYAoWLERP7P53KVLil2uZNG9ZdKRoPhIFq2uKtD8aOGjJwx7Yt4ddlvT67aIljOExUKlSsJCFPLAUgULxU2QrJDRuG9kXv4eOnfddnyOjUISFxQr8ULFK85A+DRv9Zu16Dxwx0Q+AyQWCxjBPPAcImbZSMAT69S5cj1qW5KlQ8LCJd5K5jLuYIoZggBsiQFZSjPIZ6jPtkDOwY9vEUoE3KQXDgzVBJcri/H4zzfHcohxFfDfW0peGggE9DJ9GGilVDVEBI8FlFvHlGPQz5jI921EuCchoWSrUtICsI58RVwzgxfsgKiBEIFQgAjP+EZcrlL6tEiGp1MD7VrAgUHad/TUpmaFgr5s/cdS54RjwjOa9kCBTa5J6xQVzgofKniKFXcDv70xZz5J3W17VgDcGdNbVkCBgChoAhYAgYAoaAIWAIGAKJQMAIi0SAZEUMAUPAEPgvIXB15szXogkhGs+H9u6O4NTsfzZlvOqqTIXFQH8l6RI0eaXlexkyZrzqx2+//Oy6LNmuTy0psV4BdR9+7Okhf/y9OE2atGpc+8+u3aUcWK6b8uTLfF2WrOKFk6xwUA80fOrZClVuu+OOWvc9APGhY08l6YdBv/1ZpfqdtSrdejux5S0ZAv95BOQkPh4PeKSVlMyJfU77T3OHZm9wp/eIATz1IRcdFepSpQp1pw+lczExeCHgyYDRHWM+Rn88DwiZBKnBVT0nICMIW/SHZLwW8LTIKxnD/UJ/X7SDtwGZpHUhGry6D/RDwksCgz3hoPAu4J4+IBnUKwIChAQpoJoReC2o8LUKZCuxoV4ZSmhAUEACUJ6QVPTJeHR81NP/1zBu9apQkgLSg3vmQta6EAyULyAZQoQy4EkYKPpjXCTVoCDcVYyLjUntwj6+z614bI18Zh6rJENO4CE2TTJrxtqxhgv8a+pvyi6GgCFgCBgChoAhYAgYAoaAIXAuBIywsP1hCBgChsBlhsDSBfNmP1C9bKH7qpTIe+jgAQwk/9lUunzlqpx4X7Ni6RVxuvT6HDfc+GTTl18f2u/H733eFXKyH/AP7t/HidsEU90GTzTauG71yqioSDXeJVgnJRQoUbYCJ71dcgkL9d5ZMn/urDUrlp3ZayEhadKEpkuf/vTpU6d+GzLgp5SApc3xykBADNyTZSaEV4KU5nR/PndsVSp3ercQAGJ7jz2d2Z3aecDFHE7tok9kFAIDUgJxZxW6hozA+I4xHqM/hnd+r/ACgMyoJpmT/2rYx4sAAzuGe0JGQQhQVvUhvGSF6kFAAqg2BaGs8DSjDoLUEBe5/Z8hQyAqSPSn90oaMGb14lCvDUgPPCQYO/VVyJqQUerRoOQJ5ZSQ4JkSwjxn/OoVojoeXi8s9bTAowK8IV0gi9DIIJwTYZ74vYYkQfMjlYs6cNodnh/qtn6LtwokR2XJjJcEzuDHnFi7Of619L+2iyFgCBgChoAhYAgYAoaAIWAIJISAulwnVM7eGwKGgCFgCPyHENi2OYywH//5VK5y1dsY5LrVK5b+5webiAE2f+vDz06dOnWyd5ev21JcokNxAteJswuGrXMmvCoqVLn1DjOcnw1TiTLlK6FzsiqZOid/jB4+OK24Hf02dGAfLxnE/aO1qpYWjfSMhCVLaI3svSHwX0JADN2dYyf7DOeQCBASN7iDU9K7jEWvcemyp3Ix0WldzNFIlzo0REz48m96sdWHpFXdBP6ND2mgh5P0HtICozoGfgzuaszH0wAiAWIAYzteBpRTPQslFzREFJ81hBRlICcIE0WiDHUhSyAbSOpV4Q0vpW1TXskFfa/6GerdwXvKMS9+d5VAUc8K9cTw9uXv2udRoeGhlOSgPnPktxuyAeJFQ2WVlXvwUp0OQmpBxtzook8ec4fmhLjwDjtc5BFIIfCkb0L9QWpAXodJxktlo6xhPx2EXQ0BQ8AQMAQMAUPAEDAEDAFDIHEImIdF4nCyUoaAIWAI/GcQKFW+UpXLJaRQ2Ur/EhYb1qwi7vg5U0JzukrEIxJq42K+L1y8VJkHHn36ud4itC38BAYsR2gorsePHcXwdc50c74ChUJD06VLjE4DBvbM116HMfE/kdCIKF2hctWcIjB+rgGVk/W+IfdNhKRJUipZruItmzeuX0uYsyRV9BcW+I8MEa+XkydOcBo6TkLI+1xkRXL3lThvpCHkVHLGa3UMgSQgQOgmyABO7R91eyeuc3tG7BRPiygXe0yIhdBId3xjahd7IFa8LfCYIEwT3yN+LzGkQ0xAHPBvfiUSVKQarwrVbeC3TMvwPcILg/2tHhRKJChB4PW4oA/NhEKCNKFviA+8EzQsk5IFTF89KbQP/S5RHoJBxba1HwgH5sQ7xqaC3/p/GQ0txXudh4aA4rNXeJt71fmAqIG0YNzF/H1QHrKCeYCl6nlscyfWR7iIn0Pcwel4ehDyCi0Q2qA9PjNu1oo1Y+0sGQKGgCFgCBgChoAhYAgYAoZAEhEwwiKJgFlxQ8AQMAT+lwgUK1Wm/IDRU+Y8+szzzYON47FnXnzlueZvvut9h8hz++/7DGrVpn0nNbBf6DlANjz85LMvdP/lt4nDJ89d3rZL759F3iF7qXKVbiFcUnwaD4SLek40If5csHb7vI17TnbqPehX9DkCx3f/I080nrosbI8alzHmv/vZ110GT5i56Ls+Q8fkK1gEQ9NFTa1at/2GMFBD+/fqph3JUH1jjY6Oxnh2ViolhvjvB4wc37nvsN9bf9XlRwqgt9Cx58ARX/cYMPzTTj/0DSac/kXnXgPbyZp5G0SH4aeRf8z4e/X2Q72GjZtKeCp9f1Pe/AWpM2Pl1gM/jZgwXRw/iKkebwK/5m9/9Dl7aZgIuL/23iftg+FOA6zP5IXrd/b/bfLsCXNXbe74488jIVQCG2e9e0vfTZq3fI93iJO3bN2245iZS9aP/OuflYH7UuuzB4qVLFt++eIF887gKsA+2viF5p916tHv8WdffDUpxMB1WbNd/8aHn3cAh5dbffDpuXBIzr5CxJt9Pm/97hNTl4XvrXr7Xfdc1I1njadoBOSEPpoIP0iGJCXUUgZ3dMl17tT2ky70+mgXfSitS5PxpDu1X3QVThd2kfsgLRCvxtjOaX/CBmJ0x5C+WTJeASQM8hAT/F9AQzTxHIIAQkAJABW15h2Gfm84JS2DsR6tDA3HRtu0Q7/c62dtQ70m1MPCq+lDWdqDnGD8zIM5oImB1wI4oNfBFSJGNS/U8yNQaFv/r6MEifczv2PgxXjwkICY4DddPSUYF3PYJHmhOxl+tdv4UTYXMZjyhJAqKBlvCvpGCwTcWCPG9oN/7ZizJUPAEDAEDAFDwBAwBAwBQ8AQSAICFhIqCWBZUUPAEDAE/tcI7I6I4ASnuylPfkKExEmQBhhqCYPTt/u3X/GyZNkKlXsOGTsF8Ws+h6YLTdf+w1avXMh5ZM2WPce3Pw3+rXjpchX/njppwpawjevr1H/kiSIlSpWFIFk8f87fwfpjvB1/HDji9pr31ps09tfhsS42tna9Bo/d88DDj40bOWSgt06J0uUrokcQExMdjXH+x6Fj/8pxQ67cnJy/vWad+5dIH2Eb1q6+kPPytoWYc+Xbatzd8vknH0IPQd+lSpXaZ/wSg3rQAwBFSpQuC8myb+/uXQJTTtYmnVj7c+fJVwBD/Yljx44KDGcJcJcWLxqvUDlG+3eEoDksmiUSDmxTxarVa7zz6Ved327WuCFC3h992aXn1vCNGxbO/Xt6jXvq1sfY37vrv2GrAhPhl7r0Gz4WggHNiKio6ChICTwGvv3io7e95SHIWrz7cTt0IaZOHPvbXXXuf+juex94mLH1+f6b9t6yWa/PkRMBctGB35495425IFXwKpk7c+okcSxJ/9r7n34pocGWzZI94q1XoFDR4uwTJSxo5/sBI8YXLVmmHGGi6jV88plrrs2S5cfvvvwsofUtW6nKrZBBtEHZ8rfcevvEMaOGblq/BkHcs7FI4r4C9679R4w7sG/vnkF9fuh8T72HH/ug/Xc/1Lu19Fnfx4TGau8NgcQiIIbvfyQ0VD8pX1vyNe7o6hwucn86d3hJWpcxfxoRgM7oYqMi3cktx1yGPLlcFDb+kI0uTSikpmpAYMjHG4ArBncM8xjrMbZTASM9GfIVw70SB5AZ6iGh3g7qbaGeC5ALGO7RbKA/6kCaqgaGej3olNUDQvUlvJ8pQ3mIFcgSyAnITHQiKEc4KMYO2aDjoY56bzB+5sg7JTG87etc8ByBwOH3HKKBuSNITvtKQCOovVLCQOVwx1dlckeXxbi9YygDrpTj72pRfz8qZs51Imumk7WrIWAIGAKGgCFgCBgChoAhYAgYAoaAIWAIGAJXLAKcjF+89XDsI42aNgucJAZe3nGan3cYyifMW7Xl16kLVt9R6956f/yzeuvE+WuIw33BEn3Q/jQ5aQ5hoQ03ebXV+4yF3Kzl+58E6/Ctj7/8lvcPPfHM87znFD3tvPNph86B5YdOnLWEE/7Mf/ycleFTl4btqXzrHXdRLrMoXyflBH5SJ49o8++zlm3sOXgMIrhxEmQJc8BQnlC71B80fgZirudMeEfQZpsOXXtREKJk4eaD0X1H/fk37yA8eA8Gjzzd5KUFYfsjG7/02ltg4COI5B3eJ8E6yXlj7pumLd+8b/LiDREY87UMe2bmqm0HIS289VgL2lNvDtr/qnu/ocw7sH2IBcpWv7t23UHjZy6cH7bvdM26Dz5COTCcs27XsWBr2+Cp516kHuTIVZkyXY2HDmOkHT6zb6cs3sjp6nMm9gN9zFqz8wgET+6b8+YHm97Dx0/DyyhY5aTsqxulwekrtuzHI0XDdT3+3EstGHtCHi0Jjd3eGwKJQUBIi/qSv5M8OnZx3T9jD8ycEbtr1Ga57og9unZH7MFZEZK3xJ7aszX2xLalwmHsF85vs+Sjkrlf4L/fK9fjko/43/8p18WS50g+Jvm0/0o97k9KPuXPfCbzjue0c0jyQskT/X3wmee0RbnIIO1Ql3Yox3vapzyZca2TvELyWMkdJC+VvEnyYX8+6K9/wn/VcVKXthkDz7Rt7Y9+uAeXjZK3SF4rebvkMMm7Ja/09907NvJw39gji/+MDe/QU3AfIHmM5G6SR0r+XfLrkof41uTftamfmLW0MoaAIWAIGAKGgCFgCBgChoAhED8CFhLKdochYAgYApcRAsVKla3AcFcuWTg/cNhCWJTnGSfhub767sdtJSpP5hbPPFJ3+qQJv8/7e9rkbHLy/EIa999v26lb3oKFi37QoulTXo+A0UMG9tHxLZk/d1bgWMtUvKXak01ffn3YgF7dfx3cvzfvxUAUS6ghOfAfJ7wSIX4wOM+ePmXiR1927plRjNjPN7yvxj+zpv9FvUMH9u+j7sVaxmdffuOdG8Ra/VWbd14L7EMcJjiJ7MSO7/NgOVcqWqpsefFoSJCwIOQQ7ezYuiUcPD7++vveu3Zs3/r6c4/WQzsjTZoQH6mAkfy9zzt+/3Grl58b0LNLRzDIeeNNPo2JvXt2EUYmTsKjo23X3r+go9Hs8QdqLpo3a4YWWDBn5jRCOOW6KQ+x18+kG+WzLEfUnl07fZ49J44fP/Zu82cfmzH5j7GB7RcvVc63N6vVqFUH8qHt+2++PHncbyN4dvrUyZNoSbCWgfXQZDkl4hPrVq9c9mH7zj1y35wv/8tP1r9n5pSJ49CmWC/P8QaB9IgPX/Yg4cROygCbNKhdHT2L3bsidrDXK1S57Q7hLgjdEicldV999FWXnngFvdn0iQdlGQhR42R5fKGxJCJY0JBg8Y3XnhsCyUFATu2PlnrDJIe5feNSSWiom8WPILOLOZnWHZwa4qKPZXCxpzK5mFOpxNviGhdz5ICLjmRv8v3limcAXhB4QODBgG4DZCB6DGguFPeXI9QSHgj8ruJ9QRm8Mfh/A94PhJLiSpu8p728/nYIDYWXBe/5rcIbgr74rdRwUng/qGaFN8QU/VKWkEpo+DAGQlnxu0b/hGdaJhmvC3QneEY7jIOyZMbCOL0eGCr4LY9946V9NDvwrNAwULyjLxXinuWiju50p8KulhBQad2Gd7bIO0IPEvqpqmTEtvm9fEgyWiB4mAzzrxFtWTIEDAFDwBAwBAwBQ8AQMAQMgWQiYCGhkgmcVTMEDAFD4H+BQKnylX3GXYy4gf0XLVm6HM8IuZNfwuw82vj55u0/bNlcZBeIv+18otYXUCQYQzDhiKZPGj8GMsE7niN+8WSM3csW/TMncKxvfPB5B8LqdG7X5ozeBkZnvAfWS9ggb3k8ATA8p5OwQpzYf7Vxg/s2inX7UuBP6KYmr7z53uC+PbsGCyuEAZ9xXJOAQDahkSAYli+aPzehcRfwExZrVi5d3Pil19+6QViEFx6te6cKfefJX6gIbUBAEJZp3KihP2ub+QsXxeDotoWHbQzsB42R8pWrVW/3QcvmG9bGFUEX0XAMfy5Q6JsQVHhd4GGhpEV844cwg5h46PFGTcf/OuyX34YM+MlbFu8MEdUmXEqchM7HquVLFla/q3bdex9s+OTHLV9+brV81kISMSs0MvK0ROI6qeK/ceoLz3Ltdz8NEUNuqlTNnqxfa+3KZUsocJ+0BUbsQSHrpgT2m5R9hX4IWhXs1+1bN2OY9KUi8p1D1wRiJaF1tfeGwIVAQAzis+UUf2Zpa41b26KBK9zlZpchf0aXPl86lzr0pIvcG+1Sbwl1IRlSu1ObY1yanIddSE5IA0IfEQKJ8GXoLxAeCsM+JCIEOARDWckY9wnnBCnB7xvvCaOkdSECIA95BzkAOcH3mueQDxomiivfWZ5zr2LajINn/F3C+K8i2pAVtMWVdiEn6ANigP4gFyAbIBoI1URIJg1dxf9nqKPkhdzG0dpQwW0NUcXcuIdoIBQUBC+kMyQJ4/pXe+PQ3ze7XYPSu50DISvwooPM4B19MWc+g+1IyZtZGzq2ZAgYAoaAIWAIGAKGgCFgCBgC54eAeVicH35W2xAwBAyBS4pAmQqVq64U/QC0EAI7LlK8dNnwjevXYlgmDNPalcuXjBrUzxdWiJQzV+6bMUBfKG+EF994t02MpM7tPvaJLHtT9pw35OIzhujjotPgfVda5kAIpf49On/tfffCa+98JHbzw9MmjuMU8ZmEQVukK6IRSB47YvCAQA2Ei7kArcWjQ7iXgz06tf04WD8yXIxX7tosWTGqxZs0/NLShfMSNGgVKFK0BA1FbN+2pfFLLVoxZ7QptHGIIu4hdrp1/KK1t9NK1arfyefAfjDcP9Ps9bfD1q9dPXJQX5/4tzeph8ipU6fikALz/p7qC4NFeKZzzQ/tCvQ68II4sG/fnrbvv35WyDI8Gth/3nbw6kAwfa1oZLz96Vff4Qk0Zvgv/bxlcuXJlx9dlPj6R+A9T/6ChT96/YVGSlYwX8KSUQfPH10nbxtJ2VeNm73+FuLxEFfaBgRbzXvrNxg7YtCAc2Fj7wyBi4AAJDDG+b/dutcWusjdO1zMiRMu+shBl+7GVOJxkd6likntTm4PcVF7MrjThzH2402BcR5CYKZk1ZXA8I4+BCH91kleLpnfAdWQgCRQIz1eDdSnb4gD2uAeAgKyAeM9V9XBwLAPOUAbeEXQL+1CKmb3l1VNDUgJ6tMuiTHjweDTo5G0wtMW46Nf3lGHrHoW9O/VBVKdDBXjZg5obkBiMDbGClkBaUHeKnmn29HviFvV5KiQFcyNseSRTN3t/ivlwAWNJvo+i5j3j9suhoAhYAgYAoaAIWAIGAKGgCGQRATMwyKJgFlxQ8AQMAT+VwjgZUD4nJG/nG1w5l3h4qXKTB7/2wifIVU8EV587P67IBR0vHnlZP7W8E2crD3vVKhoiVJoBiCoHEzsGj0NOvEa2rXTBxo+9Syn5TUUFM9fevP9j+976NGnPmnVvAkEgXeAzAsDNKf/v+/w2YfnPfggDZSrVPW2ex5o8NiRQwcOHDl06KAcmD8s0ZAKoB9B2KpS5SpViYmNjYkVPDntL04ux08I25ImbRqfYYxQW+caF54N+/fu2Y1IeELjJyTUzm1bN999X/0G4tyQNnDONe657wHa+PqT996AyPG2V+2OmrU58R+xYxvGtDOpprSFpsOnb7/6fGAdCl1/w40+gonwWt56UyaMGfXu5x27opXhJb8C54DXBx4UPO/TrdOXgSQVZIU4SoQeEBC8dUuUrVCJvYunQpas12f/snWrV73vEYsnTNUfo0cMDoabiF4/CpnCGk378/+JLjx/EGenzrJ4vFoSu68QEL/ltho1+//wXQe8m2iTMXUbOGrC5rAN6/rJ84TW1N4bAhcSATnJf1C8LPhOtJB83K16YbYr0qWWmOCPu8xZUrmQ60SI+1R6F5r9qIuJjHant4vB/UQBlybrdpc6Dcb+GpIJE4Whfa1kPBYwvuN1QUgnvNwQk4ZsxrhPSCbK8E5DO/FboSHe+B2EAFCygN8lPlOWZ3gocMV7Ae84vMQK+/vXcE3esH4QBLsl4+nBPaGs+I3VUFGMSb0q5NaXlLDgbx4ZooJnSsxATPAMrwqIU36vKAdhw2e+2/tdTFR6F9GnkFv3zh4XfWi1PEP3CbKC+UNWQG7gJUKG8KCNwayJDuRCXOVgAT+NnC/whs/yYuQVHA/EQMNt8Zw6NHYhhmVtGAKGgCFgCBgChoAhYAgYApcEASMsLgnM1okhYAgYAuePQJ4ChYoQVmjpgrNP6RO6COPuyiWL5jd64dWWEAnoEmivCFOjAzDzr4njzn8kzt1Zpx5xu93YkYMHBmsPAoDnwQiLqnfcfQ8aCBATGJVFh6FrtRo163T/+ovWo4f93DewPYluVYpnv4unAToIF2L8gW1g9K7/6NPPqdHd+/7Rxi80J5+rXxFffhVyY/a0SX/06NT+k8CyeJQsnj+Hk7jnTFioCgoZtGD2jKkIRw8b0Lv77ogdGMl8KccNuXKXFWxXLFn4z3wp420MnQ/wHOLxAtD3dR9+vBFhiwjVFGwAEFB4IXj7ohzEzJB+Pb/H++WW6nfWnDfzX4+LwIRmBc/w7hk99P/1S7RcgcLFfF4j61atWOqtW6psxVv4XKZ85arghleJ9z1YgMm6Vcvj1KMM+71Vm3ad8Cr65rMPW2k9vDxebvnhp4wdDZDVK5YsCj7nxO2rW6rXqIkHCaG3CI/14GONmrz50Rdfo2PR/KmHamtYsASW1l4bAuj0nPFslm19hkxODjR+0qKj1P1AbPJp3cYPN7pcTaPc6VynXepMmV3UkWMuU/Gr3bG1B12qKNGgKJjaRR2KdWnEAyM0EwZ/vBLQpuC7yT1EBh4GjAvPCMKcEXaJ/ytgnIfAYPx7JeMdgeeBGtB5DiGg4Zx0ntSlDOQEZAPeYbQLAUF/3Afq/6iHBu1ryCfIBMgUxgPBAHlB24qh9ue96js17KtWBvV5BsHgC+knCYJ3jzu9u4DbP3GvW/3SGPlMuCrGBinDOAjDBdnCWLgHEwidjrIWPiLzQiQ/QeEjW+ReyRavx4h6tWjoLV0Drl4Sg89gwLPUfs9KLRvIXvhIDf/4fe8gSy7EfKwNQ8AQMAQMAUPAEDAEDAFDIDkIGGGRHNSsjiFgCBgC/wMESsspf7oNFlaosBireYd9ChZ4AAAgAElEQVRBv1Wbtt8gSu0d4v8bjM82/CZnKtXuuLs22gBT//j912D1q9x+Zy28OwLJlZw35r5J9KvzTvh12KDPv+3ZH68KtBlaPv/kQyoW7m0Pr4psEl+KZ0NFSDk5Y01MnS5ffvI+GS8AyJ1uA0dOIMzT+680eQK3itSpUqfGgoPh+iqJY3R15szXop1w9TXXXguxgJE8VNSsg4WGoj2IhOEDev+Q0FgIbcScb8h9c570wp707f7tV946dRs83ogxeL1T9H2t+x9syP1Uj6cBn5lTFTG6g28wHQjGLnxB9SVChAULFzawZ9dvnmzy8mtNmr/5XvyExb+C20P79+omYhMY8uKkwsVLlmE/BIqOl5RwXxTcLUTHgB+7fnNWPf++DkZYvPjGe23wfnijyeP1vfNq9OKrLW/IfVOeiWNGDKn9wCOPb1izihA3cVJS9hXhvPbt3b0LjZjO/Yb9jnfFpLG/Dv/ivddfUl2RhNbV3qdsBDxEhWooQF5g4I85H+LCbyhvLd4WtV3UwVi3+ZvMLnJ/NnddzdMuNEdGF3VMDNaxJ0V4O6s7tSXEpc0moaLE0yEyi5Aa10a4kDRKCkAmYAiHcMAIj9EabygM5Xg4YOzH0E/YJu7JGPzxUsCYT3n1rlBDuWpYqHYF89XQUVzJ6g3BBlEDPM9oH9KEvhkXBIESKXhdaNgo9aSgfjADuz6jHO1o+Cj0OHiGx5uIlR9dJloVFdyeMaFu7zj6reQfD+8ZJ/UgJSBe8Mbg+TTBP452E4NIbvLvEfUKUW0QsCMrbjzXcJA6JyUbIH+4V1z5Hdb/5+maaOgsJTbUW0a9YRg+78Sh8Ayc9GMeGsldWKtnCBgChoAhYAgYAoaAIZAsBIywSBZsVskQMAQMgUuPQJmKt1TjNDmx9AN7xyDMM07yL5g7a/ryxQvmecvEd8I9ubPg5PvqFUsXBYb+oT0Ev8kIOweGdypTsQrCpa5pi7c+4ET/T993bNe/R5eOaFcEGwv98BwR5vVrVp5leE7u+OOrR7inR55+7iW8FV55+qE6i/6ZTcz1cyYwh4R5vM5tvjBYgam0hPHi2RJZmITaKi3MAWWKlihd7pc+P3RGmNxbBy8QiCJCNQW2dc/9Dz9KSKdAr5YiJUr5tCX+mTXjr2D9V6x6Ww3ez5zyx9hg71nDYf17dX/ulZbvgUugKLpvvH7Bd4ioYG1UvrXG3eEb160JXGd0JCj/Q8e2bTTckre+7mvZSnE8LAgxBVGE1wqi71oHQqzJK63e57lwd1sgYPjOBI4pKfuqrOzZrNmy5/iic6+B7AdEwYN5DiW0tvY+5SHgMUJjiMb4TiZxst8XrkjK+Iz250lcTBTSglBHJd2Ovutd2uxZXPo8MS79zftchrw5XMypTO5E2F4XmjO1O31Q+kt71IWczC3B7E64kPRq9FdvB4zYGOTxLmCMeGHw/wVIAwgLvDMw3q+STJ8QHMwLA7kSCepxoULYtI2nGKGlKEf7xSTrez3xD6kAWUGb6nmhbfGO/r2EiNZTo31gmCTmRtgmDQ3FPaGs8KigvT3u+Jqr3L4Jdd3GT8dICCh+fyEk0Pog/BXzwkMLDzJwYVwQNSsuFFnh2SPSrK9fEhgwVzJkkpJBaCUxJsYAjkpwME/Whed4oaiHjIau4j1ED5iydpBHtMN8aFsxpzxYqjcKY/ERUn4y+4xXkHlg+FfKLoaAIWAIGAKGgCFgCBgCFwUBE92+KLBao4aAIWAIXHgEEKuOz+iNARYi4345gf9Tl6/bBvaOkDMGhzUrli4+35ERluiqTJmuji/EUYOnnnuRPhA7Duwrxw03ipHMuU6ff/hW7UpFcncXQ3V8ZAXlMLZznThm5NDzHXdi6hOaivBHCILPmfHXn4mps3dXxM5M11yDMS9oQncEIgQR9ITaoyxlokVoAs8Gb3nCbN2cr0AhjOWBWhMIXuOdgXcFhIa3HpomfI5v7R96vHFT9kYwEkTbGdSnRxe0LwiHFDgHQjahWYKgN/oZge/TSVymilWr1whsHy8IwpRt2xy2ceyoIUFDixUSJmTv7oid+/bsIlTNmUSILtrt9d1Xn+tDxvFJx2590oamDf2q9dstGBP1ghEhSdlX7HfxDJnfqN6dtzRtUOd2IysS2sX2PgABjM4Yi7liSCbz72+Mxxio+ZzGGy4qmQgOkXr/SN7oNn+10B1ZsMdFHkrljq3e5Q7O2utO783kog6IAHeEaFqIPMTpwyHu1NZYF3k0nYuNgWiAfCDUEuPid4jfXkI/oQXDe0iWjZIhUTH2F/CPk/FjBOcZYZ7w0oAY0M/MlfolJUNcZJEMGUB7/FZRl3v11FACRL0vNCySkhHqwRXoUaH/p9FyXGlXjf28pw+I480y55Vuz68ZRFg7xK1reUzICkJOMU5+LyFW1LDPM8a00z9/MAbrC5kghPCMYJ9wTwYjRMeLSwYDNEbIkBaQPYTVYg0g9RkvnoiEr+JvLBiDE2vBvApJZn2pR3n+XtE+z1lv9iZrTduKHwQI7XBln1JGyQ0IjBD2LCGsPN4YUsSSIWAIGAKGgCFgCBgChoAhcP4IGGFx/hhaC4aAIWAIXHQEJApRZrwWls4PfkofDQLCEe3YuiU8mFcAHhbbt4RvwqvhfAerYY+2bw5HQDVOQmPjQTGA8zBYGB+JdoTRxKHNEMw7I7C9oiX+Fe/+K57QU+c7F2/9fAWLFPuqe78hC+fNmpEUce+9YhTPmDFTYBz2M00Trmvj2tUrg4VKChx/GSGleDZx9Mgh6EF43xMOis9/jv11WGC9mnXrP+LDKYjnxfX+kFoS1QiDW5yE50ANke+YNXXSBIS+48MT0gBdlNtr1rk/sEwuEfNmfy5d9M+cYPVr13v4MQiusaJB4n0vQuY+7wrEvIMJgfOuUDHx5Fm+9CwNivsfeaLx9q2bwxiTtik6Ii3Q2ejcrs27a1cuW4L2Cd+HYGNK7L6SKF/p0DVBLwTdkAu536ytKwsBjLaejDFXT8ljBIYIwEjMv7sx/qqHM8Zg1Sc4L9JCTvxj4IdkXSH5iNvRZ6lb3XiNO7Ziv7umfKTLVHSPS50xUogLIQmi07vInZHiXXDMHZq6U8qcFOIitYSO4oQ+hnOIBcaKoR6PBAz9eflKSsYwriGENBQUpAXkA0LZXsIUIzd1CUXEPPGk43eN3wra9panP/4+MQ/IAkgPiErao6yGjFKvDK/uAveQJRouiStzYQ1oE68J2hrvTm1b7PaOPuRmZEntlj180h2aQ3+Mj79NlKfcNMnoVSixxDMwAds//VjL7QVJ2gf7BHIEIoGxQFSAN96T6IygqZHLPyYV/F4vn5k3ZBAkE2sHkQHpQn1C9T0gmb8dfMarAhJECQ36UUKIe/XOYEzsWYgQ9ihECuPjORhpaC3ueQZxQT7zHZBnlgwBQ8AQMAQMAUPAEDAEDIFkI2AhoZINnVU0BAwBQ+DSIUDoHLQLliw8W3AbYWGMxoxmYK/vOwUbFYRFMO2L5MxAtI59YSsw1AfWf+Wd1l8ghszzVUvP9rC4RhgL3kUG0TkINhZCDW0N37SBnJyxJrYO+PQYPHoS3hJvv9TokUAvhXO1gzEfozZETrBwXRBNgSG6grUHbgWKFMfw5EYO6vujtwzeAxALGPaDkTd31LrvATwJ5v09fUpg2xLtyReG5oQwRIHvnn/9nY/SpEmb9pfe3b5LCKslQpbhgYJng9drAU8G6gZbI/bs0y+88iZ1t4RtxLh2JpUsW6EyH4Jpl/CcMFvohQSGoIJYklf5f+nd/TvV3KhU7fY7W7Vu983MKRPH8Rwss16fI+fCubNmnM++Sup+TQhDe3/FI4ABn4whl39jY6RXzwrVcOA5v5GcfsdAzXtIAYzQkbKnTyY3PJQY0o9LaChICwz8lV1sdAYX9kU2CQcV6TLfUdTFHDrlUqVP5SIPbHOnInL7QkSdWJvKpU53xMWcvMqFXJ3BpU5/wmXIh4EfQ3iYZE7kM2YNHwSRoFoW6oWgIa+YFwQBp/UxhCsZoAekML6DQx7J9AEZiSEcY7mSDLSBgRwSgiu/X/QTKCgNxj59Bcm0D5EBKYsXYTX/+BkL4wbb6W7Jfesk/BOYY3BnfBAAzIe2CFOFNwJjpy1CWGn4KvqHsJwtGJ+l0SPPk5X8XjWQDMwZjBkLc9JQW/zd4287OJAZU17JkCeMA28K9dThOfuIPcdvK1nDeIEPHo+Ex6Mef4fpD+8Z+sfzAjy2+Otr2EmekehDNU4oD/HE3xP9f6R6w/j0L/x1TLTbD4RdDAFDwBAwBAwBQ8AQMASSjoARFknHzGoYAoaAIXDJEShVvnIVBH43B4nHj0EcwzCG82DGX+L9kzetW0PM8fNOp06dxJDlIEq8jUGqPPJ002ZiNz/Ou00b1q4O7Oy4xH/iGUb0E8ePn2VA95ZHLDpfoSLFxgz7pd95D/ocDVS+rcbdX3XrO+SouJ+8/NSD9wjMGNISnXbt2E48dFe8VNkKs6dPOUuEldBH0zxC2BjhhWDKF+iBglYC6xgh2guBYuUY9/GG4KR/oK4Fug142OAlEUxUe9+ePcSgd4Rf8mqKoEfxaKOmL/8za/pfXk8FymLsz3T11dds3rQBI54voTiOcHagN4TqTEjUKwywcdLDTz77AuHKnnv4ntsC35WQOTHXYBoTlGV8XNFC8dYtXqZcRT4rCQTZ9HXPgSN2istF6zdebMy7HAI612AeRUnZV8ePHfHv1wyqPZDofWEFUxwCGGtVU0CFqfmt5KQ/ib2EMZd/e2N8xrhMeCUM9pxkpxxlMOif9V1KLJp+g/pUIS743rwpOYOL+CXCHRAJmxuaZHGZqxR2qTNkdWkypXMh6VK7dDfFitdFVndsXai7unyskBcR7vCCvC5TicMuff6CLnVoqHz5Ccn3tGSM/UqyQDCovgLDUwFujO0Y+PnOYLRWnQk1Zit5ASmAwTxcMqGm8CbgVD+GcTCAGKcdyBEIBgzt3CsppFoWGvYJYzseG7Q52ddGTPQxF3sigzu+4Ua3a2BZISsgMPDsggTAKA/BgfGediEvuPJ3i7koCUPf3QTXOHpC8uxCJPUagVQBN/piPhATZMbB7yBeESR+yylLOYgk5kJ5sGYeeGJASrC38BBhjSCUlRRiDfGiUK8O5k/bd0kGa7zsIM3BATwhJnjO2CByWKdtktlbef3ts29pD7JFw1CdVm0WeeZM7wIULBkChoAhYAgYAoaAIWAIJAUBCwmVFLSsrCFgCBgC/yMERIu5OiFp9ES5dxgFihTDSOEw7AfzDFDBbeEzMICcd8KIHRUVGXlHzXvraWMY09t36zv4sBj7OREPaRGos0BZNYCr6LHWR5/h82979s+ZKzeGO1+CrOD0P4Lb5z3oIA1IFKNrW7Zp902PQaMnRezYtrXJw7Wrc01qXxKZCCOOQ2MksC4ERGqx9GfI+K/XCWRFr2Hj/mrToWuvwLLoPPDsjzEjhgSuc7nK1arzLhghVabCLZwmPmPAD2x3zYolvpBKeGHoO8bRrmvvX04J+9T2/TeaBdb5oF2n7v1+nTQLkoN32SSs1MNPPvMCXjrocXjLFyle2qczks+vlaHvSpQpX6lVm/adRg8d2CeQgAGWYiXLlj+XHkTh4qV8QvJoXHj7k6hiGN/cQWFu0O7oPXz8NDxQWjzb8H4lmySSE8ZQd8xPkHnrJ2VfEbYMIjBwvxLiChHyZ19+451A7OxzikVACQv1oMCATHgejL0QFF4tCIzAGtaHehjnITMw1IdeAD0L5zewd5b2Jkje507t3OfC265zm95b6Q7NOOCiDh12J8MOifk/q4s+eshlKnnYRR2MclFHcrrQ629we0be5A7NzOVOhMtIdxAKjr8fkAQYyNWzgXBBXsFsxs/8lajQd7opICNUBJt3kN7gVEQyvysY2nmmWcNoKXEBZl6tDJ6TmCdeYniEMIZoGXNemef1LvzLm9zuQfnczp/5Pw/EKcb4uf6+CJ1EG9ovV9qHOOIe7DpfJLJCMdGwWuwBCAoVQee3F0ICfCijXhjL5R7cGSfP8XRkbcL9z+vKld/OmpIhgfi9ZD1qSeZvwL2S+TcDRAhhotibkDGQITy/XXIdyQiN005h/zPCS+WVrNoZYFlJMmMmTBjeHqwXa8f4vOGiAveBvLZkCBgChoAhYAgYAoaAIWAIxI+AeVjY7jAEDAFD4DJAoGDR4iXF7jy/bZfeP2NA/faLj97WYRMih1PvI3+JG0ZI3ythESxcUXKmzqn16X+OH1Pr/ocafnBgX/ewDevWPP3Cq28Swufzd1978XYhMlKHpA7BiBxoeJ88fvTIdz//uut7n3fs2qNTu08IuXN/gycaVal+Zy08Do6IxVnHpCf3A43dyRmzt07jl157C3Kg/C3VqguPcPWIn3/qgQg4JEty2lYCp0SZChhv4iQcEiA07qxz/4NChmypVffBhvkLFy3+0mP17g4sW6biv8TDuJFnC1Br2CVCHgXWEy6Bk8EuXNYh2PjxRMBL4eVWH36KB4ZIY2xr1vL9T/IVKFy01YtPNwgM1UQbeITcVafeQ72HjZ8Wvmn9WvDCM+HtZo0bBvaBgDX6HHUffuxpSDUIq0q33nHX8y3e/nDnti2bvXtV6+aVvgmjtdpPpgQbNxoUPA/0xNkTEeHT9vi4w/e9s2TLlp2w6c2ferC2d/6bN61fh0cSguILxCtlxuQ/xiZ3X00YPWLwU02bvwFBgTZGucpVb3vkqSYvodfy6duvPp+cPWN1rkgE+De1nphX/QrC82BY5qoGXYzDGM3xJsBIr6GN1LOA0/N4ZmhonWSDJYb2Xf4QUXgNPCb5Zndk5SF3+uAMd1WpOi7djalcxgIHXKo0oS5qf1YR4xbDdvQJly5/qLxPL+Gh0riY4xmE2Ih2UYczu9BcofIs1oWk5TuIYRqPBYzRjJ05cYVUCPRIwmDOO+aKgZsykIrMESJHjfac3qcs5SANwA0sMIBzpRyEhPaJBwG/iRjWhXiJLOliDoZICKy8UuxqIS1CXOT+KBcxeLuLPsh41buF30wM9Iyf8dAPHoiEUaJ/PA3wKtkqGOJlcLES82eujE1DV/GM8eEFwvwYI6QB+P4fe+cBH1XRtfF9pYNilw6hd0LvvfcmRUFQmgp2VBRRiiJFAUGkiRRBAUF6772XBEjoJTTpVXr9zj/u8F2W3WQ3yZJscsbfcXfvnTt35pm5S/Y8c84DVqR24t8qIkSoS8QZ7zEIDtYP2PL9iQh3aApHKURSsOaIquC4n71d7gsZAh7oZ1Cowz2ZRzYMQG4g8A32XFdPDKJjgb0+dVnLRLhwf9Y6ERq0DSEUqm8h5b5GW9gR0xdFQBFQBBQBRUARUAQUgTARUMJCF4gioAgoAj6AgGz8P1KuSo06OMc7tX+zibXLiSS/0rhfB/cXf3iIs6G8lCIFux9tYTmHPYXg5z7dOxNR0LhF2/Zci1N5wLdffYqAMgLM9DVVmnQZHPtE1MXgPj2+6vjN9/1+Hjsl1IlMVMPA77/pNHH08J+twtSkOSJdkGNKIE/76lgf5zuaB0QrjB028Adn4uCe3AM9B4gECBpn1w3u2+Mrohne79T1e8imT9q8Xj9g8/o11rqIO+fMW6AQfXI23hSpUqeFCHCMNqCNixJpADG0d9eOQFf9/lYc64PHTZ33hRBF1EFgm/RXpJhydg0C2bmkP03fevv9dBkzZdkmWhD9enT+ZP+eYHb3Piw47VOkSpMW3YjSFavW/Kbvzw+1N0gz9fVHb7eEOHC8h4nGOH/2TGi6KmeFKAwIH8frlwuZsm7FkgUFi5Uquzd4Z2C/Hl9+4qgRAvnUrWP7Vj0H/TquSMlyFa2EhafrauzQn/pWqFqr3odfdu9NPyEHVy1dMOfXgX2+dSYI7sna0bq+jYA8diaqwmgo4HjGcct3rkkrZFJCQVTgnDa6FtZ0QKSh47j5uxwBbpy7UUFa4HAPFuICfaNqYrVtt068Yrt/Y5vt+tOZbZfX7rfdv51eyIt7thRNk0mUhaSFSnbbFv+5+LYHMpQzU6+KaPdLtms7/rVdC7xmi5/yjC15HtE8SJxA9DCO2OLFp9+MlfHhKCcCg/GbHfZmTIwXBzyfcWrjwebVpM/iM056iAra4zhRDvQfxzlYGOc6hALtnBN+5Y7txsE0tnhJc9vunD1ju3//Oduto3dsD+4klNRWiSUV1kkhK+gj1zNfOPZpj+uJ3sKJD6FDGjnmiqiKhUJUmHmTj94pzK/MM5gwZhNtwmdDHpgIE3CCuAgRMwLhRCNCXNB/yAhICIMZ4+R7l3bBFCIiVD9KysMoRnkPQQQRBBFiyArqMH+hfzdIIQrDFIh2sDQR+syHSVHF3PNvkCFciBAJEUO7iDGFpvKCuFDSwoKovlUEFAFFQBFQBBQBRUARcIqAhujqwlAEFAFFwAcQeFk81un8MmUJFEc3TlxPupxQCA2ROcjgSivAk7asddkhTyonnMM4so0+AqmW6svOdhFy/slVX9NmyJg5k6R8Ik3VPnHEO+oicB+IBaJCopqwgFigeIpjWDhBOEAaOKZLMtcwB+ByUTz0zu6Lc77Wq6+1WLFw7kyrzoS5XrifjGhIOCMsiHzIkde/4M5tm0lz4rKQxoj0UczXDqlLWq/w5p5rGBepkZzVLVS8dDlSMn0mkRqQHxWq1a4vWbwS7NqxbUtYznzWThYRGA/evm2zq3mADCEV1aH9EddeeSpevHgP5AbWSJ+IrCswJgJGhpZw766dgRfOiWNUS5xGwE5W8Hc0DmScuLzi9MWZa0SNQ1OTSYHEwAHOcRzwOKRxNpMuip3zvOc8TmauvytfUexmj9IipAX9aWi/L/cmXRBOa9L74MDnO4GUP3eEwBD6IWVqW/yXztuSF7ppu3f9Wdsz+SVl1KWnbEkyX5EIjByibXFDNC+S2Z569qwtfmIc6kRCmGgBgw33MNEn5ncH5ASOcogDjllTSEF40IZJ/QS2nAcPQyLclxRXq203Q0pI5McF2/1rct8HZ2wJU+WQ9FZXbTePJRRC5oLt6GAhM/aBOWmTDFlEdAht0h7EMdEAkBiQI9i0qBTWDm8CZR0ZAgKcWD+kJYRIgViAIIBwMETQUjtupey4+ckrqZoYC+mwGIdJ0wQZzfUQD+hWcB/HEiIHaIMCacb8W4kLJ5c8cogoCq7j/qzdP+xtMLe0xdpeLcbaAHOT0utBVJBx4XVOzysCioAioAgoAoqAIqAI+C4CSlj47txpzxUBRUARUAQUgWhFoFmb9h993r3vwOpFc6Y7ffIEjk8tikCcQMCuM2F0GNgJDynBLncIZZzDoYLtUnBEkz4Hp7lJQYRTnvM4pSEOeM/zg9OX629726Er5AXaMxnEcHDTf9L+0A8/MZzmOJxxdOMIh3BAZ4JUQbzHSZ3clrxoMlvK19MKgXHdlijDZVsSvwsSnZHC9lQ8UgxB6uFohxCAhCE1EaSBIShoh7FCTEBQmPc4tXGAm4gTExlxw3bvrjjkHySw3dx/1nb/VmrbnfOJbPf+lfoJ49kSSlfvXo5neyrp/2xnZ962XVgYYLu2G3KI6AOIDtojiiLE3pcd8sp8bBY7IiSFywg1Oe+1Yl9HYGP0H+gz+II36wYtCdYJeC22Y1nfjhmED4QEhDLXmGgLjpPiivFCGrDGrGWefABn5p75oRBlwlwguu1YWK+0x3ow69lahygK1jyRL+vEiNgwJPcKeX/A/hlCxURlGB2U0HZcBCg66YoeUgQUAUVAEVAEFAFFQBGICwhoSqi4MMs6RkVAEVAEFAFFwAsI5MjtX4A0V0pWeAFcbTLGImCPrqB/OGlxtuNsJlc/Dn+cujiBcSCbdDs47nEsm538XEvaIwgDUilRj7ZwUNMOUUFEWXgUTecJYHYHfaAQFzi0ceajA7FSzKRsol9ETCBMzbjQyCFaAUc3/Upgu7LpgKRjSmJ7ocpN27NFk9tuZohvS5zhli1R+n9t8V+4KMQFBI4hC8CDzxAW3JP7cF8ThWIc2FYdELC4JGmekouWxjnbjUMXbAmeEy2Fu8klzdNt24O7CWwJX7lpu3MlnpAT52znF/5re3A/vu3sdHGQP8B5T7TIf238pwsBKcQY64htFLsjOMz0BLeormtPCwUhYKJbIFggGEz6qmB5D4HDcTAjRROEBCQHr1zH9ZBBEAfMG6SDESpnXUGWgQcFLEjtRzusUyPiLWm+HhbWI3NkCmScSVvFGnUs9IO5RLCb+UTvgv7TL54NIkO22Y+x7okoImomVNhCiyKgCCgCioAioAgoAoqAIuCIgBIWuiYUAUVAEVAEFAFFIEIIkIoKoe0IXawXKQI+iICdrDDphXAasyv9hBiOdowd5DhrcRDjpGdnOrvmiWjAsYtD19TDkWzSJUFm4FzmWo5FeUooZ3CLw/4vIS24HxEROLqDxIyANn0h7Q/OchNFYkgUiJr8EuWw23Z6UnKxy7an8963pf3wZduDtYltT/snt8V/+SlbvCRHxZ6yJUyJo5oIErQNwAEyBCxwoBviJ1TnQOyO7faFfRKtkc324HJ8281T52wPriSxxX/Rz/ZvwFVbvMRJbE8lkT4/uGi7uutpEQK/L5EWd22X1l6y3T4JbvSV8UBKEJ3AfZkDHPHMV0+xZTL2J4KxM9wdjoEpfeGVuYAYYh0RzYBTn/kw2LD2iGQgIoYIEQzSgogRyIQG9jEeklfwRUiciJntYmiYQKgRoUHbFMS5HQvrc68YUR4U2oVws5Ia1msgPiBIeA4oRNjQZxNZBEHBWmcMrAOeC8bKfbxGyjkZlx5SBBQBRUARUAQUAUVAEfARBJSw8JGJ0m4qAoqAIqAIKAIxCYFEiZMkyZw1R66Fs6ZOikn90r4oAt5CwJ6+B4cxfz/jeMXxjsMYRziOVxzEOJhxlrO7n/fskDcpWHFKs1ud3f441VmtCw4AACAASURBVNGywKlLO7zSBo51r6eEsmJkd9wvEuJiixz3s4+N/kAqGKFlLmHcOMILiOGgZkc/O+8hZx7Yru6MZ9vTTsiB+C/aXqh4wPZi1XSiKZHalihtPFvitLdt1w/ss73S4I7tqWdSiAbFadHIyGa7f/W2EBOCaTyJfngqke32Pzfl5Tnb3YuZRZ/ilgiCX5fP8W3X9ySyJc7ylO1/8XGGP2W7f+9/Enlxw3b7/FnblbUJbOfmEPlB39B8AHd2/DMHC+2YQlqw4z9ExovDPMYUe5QFawN9DSNWTl+NNgrpmnDus3YgEvzEIAAguZgnIjIgxCCcIA+oB06QFEQ7cAySwxSIBSPCbcUBHaTiYhBIhqww51mvpM8i4gaizrGwhlnXmCmkh0LDApKknBjPCf1gnPRRIyycAKmHFAFFQBFQBBQBRUARUAT+++GhRRFQBBQBRUARUAQUAY8QyJ47b35ErTXCwiPYtLKPImCPrMBpjBMZYsGICuMox8GLUxanLhEDOGIhMnDk46AlqgBHL07pfWL8/c0OdyPYzQ50yA6IDkN+PHGk7I78h858ITAYL9oOOLHpP85vxmkEwxkrGhc4qzlGkbHfPWO7sCiL2AXb/+KllOiKxLan4l+0xXvO33Zi1L+2eEnF2X7/eSEqDtterPSC7eres7ZEz1+3vfxaNtut48klSuK27V/JVJTwpYS2xOkS2e5cTGBLkvaG7VrQXbk2iS3RK/Ftl5Zdt/0zeqbt9jn6BUnB/ekb84JoNSmscMDvknHF+F38dtICJz4pnSAtWAcIYPNKlA7rjHNEXkBUsF6IYmBNsY4g0ALESHsF0QSRgYYFdf3EiK4whfOk53IszLOrAvmDmXkOo+rDU+hvUJ91tMzeP04S5WIVYHenLa2jCCgCioAioAgoAoqAIhCHEFDCIg5Ntg5VEVAEFAFFQBGIKgTyFihcTJy4D4IDt7LrVosiEFcQwPmKk5gIAxzIEBiQD1nFcA6zc533OM5Jp0R9nMM4e9k1D5nB7niu5xyOaK6jTZzRHIsRxe7oDxLiAtFk9Daw3GLoH+AYhwhgtz1jwIGOKDc77EkXxfjS2x7cu2e7dYIoDMHpCHWMgx1n+1nbxSUQOxA68W1XAs+JgHdyW7K8CWxPZ39gu3nsrmhTJLY9uHNVIjIS226fumG7uCzIducceNMO7XE9kQT0Bcc+ES2QRAhp4+z3mWLRszA6IoYUM0SMEdgmRRdEABE6RLlQDy0K8K8oZgS7iSpZJAZBQWoscEMQu7AdlPnyWsNDgJjb8AqEBKQLdbnfKrEQMdY964N+0H+MvlNfiyKgCCgCioAioAgoAoqAIvAQASUsdDEoAoqAIqAIKAKKgMcIQFgcObh/79V/r+Aw1KIIxCoEhIsz4zHaAXyGnDDC2DjccfxSkTROfGanO05ldsZDPmAcw4FuIjCox2ectURk4MzHuR96Q3Fa48CNUcXu+CcVEUbqKEiKymLVxdBSIMUP2BjdAj7jVGdsjNGkOeIzBQc19YnMMJod92wXl18Tk/E/Je3fh4CgHt8v3I97Q/rQFo55cOLekELzxJZIP0379tv43gvzL2vPaFqgPcH6McLkrBGj9wH5BWEGQWaEzcvY8SHChDRQRPMgMk56qPJiRhMDkmO6HUPWKpEQUVmYI1NMZAjRHhAnkF78/iTNFfPIHBvB9ajsg7alCCgCioAioAgoAoqAIuDDCChh4cOTp11XBBQBRUARUASiC4Hc+QsXDdi4jvzkWhSB2IoAznScrziMTRoniAec6JwjcoJd/efFSEvEZ+pxnpREREvgEOY8O/9xDLP7nTaIEMDRbISfccDH+NRFTLSdGJguxAX6EIg2d7CPg/5vE4O4gLQw4t1EOkDKGKICx3uIGA5s3kPgQGzwXkge0ab4j8yA1AAX2gIrdujjfDeYdZf3O6U/nqQpYggxughpcc9OWjAuE82Dgx+yAmw4RvQCa4wIBtYi2ECQgQ9EALoWrEWIDaIaWHNEXJB2CiIEEojjIWJ+YkbTwoh/c6+IFtY/88l8E51TU4w5ZG3QP97TF5P+jP6rnkVE0dbrFAFFQBFQBBQBRUARiIUIKGERCydVh6QIKAKKgCKgCHgTgRdfeiVF2vR+mcYN/7mfN++jbSsC0YgAZANkBY5znLtmdzt/O+PcNambcCrjRMYRS310KKhjUiNBULDjHScxhXM4c3FAG6ctbfmiw5Zx4xzvLwa5ADmD8DPRFTvE0JcgIsWIkOOw5hjYcHyrHZMi8grZAXGBEx5iB6c2qaLAiGPs0EcvI0iMVEgQGZAY9CHWFSEtyLgHuQCBgEMf5z7EGSQAuiJESzB+sOEV7JiDQmKsNbBmPUJYoD3CeUTViQYCWz8x1uECsVIWAMP6bYhYt1VU2xXu3AMBdOqzzvlMf1aIsTaYP+bVF9e8qzHrcUVAEVAEFAFFQBFQBBSBKERACYsoBFObUgQUAUVAEVAE4gIC+YuWKM04A7dsWBsXxqtjjP0IWFJAMVgIBCOwDWGBoDEOdRzChnAgeoBd7CXF1ovhfMeZXECMc5AcOJw5HmL/jNPY6FzgiOYeJh2OzzlvJbKBPpOSCbNJxAX4oIsAGWElL0hdBDboXnANDnZ2/JMeiIKDnWOQH4gzk/4JZzsRK1aSAid3fLlvjEubZR9HlL7YSQvWh4lAgJzhPWvH6KdwDALApN3iPedZf2BKfeaHeqxLzvNqCAPWM2uUuQBXCCXmEYKEdW8ta+RDYzFnOitmTqkPuYRxn01ik+z3h+hDb4QC4UK6KJ4Rn9IaccBEPyoCioAioAgoAoqAIqAIeAEBJSy8AKo2qQgoAoqAIqAIxGYEChYtWebK5UsXD+wJRuhViyIQmxDAwWsIC9Lu4LQl7Q7OV1LdoJPALnPICpzEnM8vtlEMJzCfSc1DdABOeXaz45glAoMd50bzwmg0mOiKBziofQVIIXgM2WKc14wHhzefL8hYLsgru+shMsApqxANRAMsk8+QGZeNKLZ8Bttn5TPOdOrjNN8vn52JMccJssKsA/uaINqCdUkxmiomDRbYQkbwyjnwgbCACDCi6KxbSAjWIKnJIM3AGlIBEo3vcdY067c2UyDGWuUaiA/WchUx5g0Rb7RLHAvRGo4FosREFhFpBGEFaeFnvyfPhk+kQXMyNj2kCCgCioAioAgoAoqAIuBFBJSw8CK42rQioAgoAoqAIhAbESgghEXg5g1r8aLFxvHpmOIsAkazAkct6XcgHDD+XsYpTGojcvuzmxzDSYwDGJICB3F6MUiOEDEcyghTQ2bgEDbi0hAexvlsnh9fJCtYJGBhUmcZIiHUAc1XgzjbQ9/biQfIitBiiAnLZ3bYP9xlbyc2zGl9BbP/J7NC14zgC5ljoi1Yexw35AXvOW9IDNYixAHrmHUNoQapgb4E10IksHYhMCAZWKOIdZPey4imQz6xttEtgnTIKQaZQSEKBjKEV0TnaYc1z7MBccX9ibqBKPGzX8f9mXP6qv+O2IHUF0VAEVAEFAFFQBFQBBSB/xBQwkJXgiKgCCgCioAioAh4hMCKRXNnrlm2cJ5HF2llRSBmI2B2ruPkZce/0a9IK+9JC4XDF+cuTnqcujhiSQeFc5YIDHQqSHNDah3y9FOPHem0Q/5+2k8pxt/enKOtUCFqH4ysgKRgDOBCAS+iSCAtcJQzNpzq92VsRiDbXlVfogIBwTUUYntbJgID7A2RQQXemzRSpi6aFswdBIMh0XhlPUMokJbLCHdnk/es6wAxUn1BYKAhQmqoVmKv2ed6uv1eEBMQfKTyYs1DSLAmWPM8E6wXiAxDfrBuIE+UsBAQtCgCioAioAgoAoqAIqAI/D8CZoeXYqIIKAKKgCKgCCgC0YAAAtbPPv/Ci4kSJ05y+eKF82dOnTxx9+6dWJH2JGmyZE+n88ucZW/wDkRi3S4JEyZK1Oq9jl+OGzGo343r13GwaXGCQNoMGTMfP3IYh6KWSCBgT7djIgXYgY7DFqc7jlciJHC0sg5xwEJAsLOceuhVEI2BITJMihuzS51nOJP9uiXyijMYZy7X855d7Nd8yaFvTwNlCBfGj8PZ7OQ36bA4DnZG8BnM7ppoi0hMk17qAQL24Ddnv/OM1gWvmFVLhXljflOLGYINIor0UKxrCAvqQGrkE+PZIIpmmhjPDOubeib9E6moWCOsAdJ8QfRNYd3b70s7kBwQW0paeDC/WlURUAQUAUVAEVAEFIHYjoBGWMT2GdbxKQKKgCKgCMQoBCAnajZo0ry1OOSffubZZxMnSUKajYfl9q2bN1ctWTBn8rjfhm5et2p5jOq8h5354IvuvYqXqVClQYXCpA9xu1SoXqfBux07d18wc8rEI4cO7HP7wjhUMW+BwsXGzVq2oWm1Uvn37dpphGzjEAJRM1Q7WWFN0QRxQcob49hF3JjzEAw4YEuIkdPfiArjhIWw4DzvcehuETPkBLvJQ8RwDOOUxQHMrnIc/b6Yvx9c2KFP//kdQdQIuDA20gFB5jA+xmmiVtjlHxp1oeXJIOAQgWG96V37modQsxIaJjUTa5JoC0g6UjxxnPnl3ymT+gkSgnVtNEuuyHuE0ok0Yl1AXlCfNU/qNNo7JUY9zvGsQHCZVFZPBhS9iyKgCCgCioAioAgoAoqAzyCghIXPTJV2VBFQBBQBRcCXEUib3i/Tu5926VG1ToMmCRIkTHhfypTxvw0LObh/77+iYC0BFkleTpEyddHS5StVrFG3YeVa9RtNmzB2ZK8uHTvcu3vXJ9OqZMmRK++FC+dw+HpUMmfPkfv+vXv3Tp44jgNYixMEChUvXY7DV69cxpmoJXIImN3maFFg5O2HuMDBimUWw5HL3804ZFmXHMdxu1YMQg4nLEQHznx2oiNizDUcI1LjvBhOWo4ZR+19IwNjdzBHbhRevNreT3AigsJEoTC25GIQNjil+Z5C5wOMeI+F4ibXa5SFF+fHk6Yd9TC41iJHBEFB1ANREcwdz4FJGQXxBOHA/HKe5wFijtRnvGcNQGIQacR5zkFgQTrTDpEarAnTvklf5YvEnSeQa11FQBFQBBQBRUARUAQUAQ8RUMLCQ8C0uiKgCCgCioAi4AkCT0n5uMt3P7zW6p0PSPn0+/BBPxYsVqps/Hjx4/f5+rP3HdsaPqB396w5cuf95ofBIxs2e6tdIiEyvv6oXQtP7hlT6qZOl8Fv57ZNGzztT27/QkX27toZSLSJp9fGlfp5JMJCuKAz/xw/GhJXxhzV47SkgjLpjSAbcJ4iQkwUBY7YQmJEDrAWIR1WiZH+iR3kpMQpKgbJgSMXpyzzYSILiDTgGNoWOPVx5OKspfhaChyTMovfDhj9Py0GaUOKH4hJiBnrDnoc3LEivZ19zmLti4Uwg0SAwDDRFzwPvGfdEjVjommohh4Fa5sCgUeqM2tKNdYGpAX6LxyH8GI9YA/1N2ItqDowRUARUAQUAUVAEVAEFIEII8CPDy2KgCKgCCgCioAi4CUEkj/3/AukOBr6Y89vapXMl2nkoB97Zs+VL//KJfNnu7rl/j3BO99uWqvito1rV9Vq2PSNanUbIW7qU0X4mPgpU6VJd+qfEzir3C5PxYsXz79Q0RIb16xY6vZFcbBinvyFiu4M2LIxDg49qoeMM5a/h3Gg4nQ1aW5wvhNpsVXM6ITgzIV4qCCGfgWRFyZ9FA5d0ujwmTZw5pIailQ45Opn9zkOfCINQoW2cRIbi+pBeaE9kzKIpnnPWBBSRu8AYodIC5zTEBZodyDYzHGMYwntGhhe6Jo2GdUI2NcnaxR9CdY9axrCwoirEynB2j4gFmJf40QOQV4RScQrERU7xCAyOAbZYSI3aA8yRKMronrytD1FQBFQBBQBRUARUARiAQIaYRELJlGHoAgoAoqAIhBzEbh04fy5OqXy4dgMLeWq1Kyb7Omnn1m12DVhQb2bN25c/+qDts1nrNy29/1O3/RcNHvqX+Lw85ld2a8IWwH5cPL4sSOezE7mrDlyJXv6meTB27dt9uS6uFT3JQE3Rao0af8eP3p4XBq3l8aKwzR0V7kUnLCQFDyvpHTC0Q7hRn5+HKxEXrCjnKgLcvMTWcH1pIjiOhz4kB8m1Q0RGewyp1DfpEjy0lC82izEDjvkGTMYvCgGWUFUCk7orGKQE+ykBxMIDI6DBWQO12rxbQQMaWXVvmBuTUQRvyuZe+rxnrVgyA6eHwgNPkOEmGfOtxHR3isCioAioAgoAoqAIqAIeAUBjbDwCqzaqCKgCCgCioAi4ByB8tVq1SONz4G9u4LCw+i0iDigc5E2Q8bMBYqWLBNe/Zh0Hoc6/TlxLAShVrdLpmw5c1P50L49u9y+KI5VzFewSHGGvDNQIywiOfU4WiEUrNEB/G3MbnB2j+N4NXoMpIUiBVQuMaNfAUnB9ZzDuGa5GAQHO8zZUU50BfV93UFrnNQQDxA5YMQzCiFpCAp23xNlQrossDP4Eq2ClgEObC0+iIA1GsgSfRFKPIgZvRIICd6TCo01D2HFZ/MMQVr4qti8D86adlkRUAQUAUVAEVAEFAHfRUAJC9+dO+25IqAIKAKKgI8hII6d/5WpWLXmmmUL57nb9fkzpkykbslylaq5e01MqJcipZ2wOHrEI8IifcbMWREkP37ksEnDExOGE6P6gH4F0TbBgVs1CiWCM2PRryBCgDRPOOFziCGYTWoj0tlAKuJkRasBRytRBThgSfVESiQIC7QuSAOFPgXHcd7jnCcFFNdBWODADY3ksAgeR7DnT+YygrksZnbQc3PGDxlD9Ai76CFsGCuvkBmIj/M+nRhps3glEoPfHIhve+W3h2N/mV9HezLIxdm7WMk9E1UBgQGJZUgLCI5Qi7Mo6cAVAUVAEVAEFAFFQBFQBNxCQFNCuQWTVlIEFAFFQBFQBCKPQK58BQq/+HKKlOtXLlvkbmu7dwZu/ffK5UtoFrh7TUyolyptugw41U8c84ywkGCSrKdF9+L27Vs4urQ4QQCNj5AD+/ZclYWhAHmOgIWswHmOU5V0TUQF+IlBPJBzHycr6aBwvuYT2y5GJAaRQ0QRmPQ3EBprxNC6wLEP8QGZAUlB2yZHv8+QFU4QtUZXECVBWqiUYpA1nIOgIU2UEWVmZ70R5wYzBLlNmixrOiEnt4r0IaNJQkO8N/N0355SL3Q+1GkeaZwfacAi2m0lI5SYiFqYtTVFQBFQBBQBRUARUATiDAJKWMSZqdaBKgKKgCKgCEQ3AqUqVK1x7+7du5vXrVzmSV8O7t0dnCZDRoRsfaZAWJDS6vatmzgv3S5p0vtlOhZyECFXLU4QQBckV76ChRfNmTZZAYoUApAVRvSXCAuc2zhYiaKgEC0AIYRznnRskBdoWBBVQWooiA2KibqApCDSgr+tDdHB+9B0OT7uIDfaBRAwRKQwVlL+gA1kBVhBZIAXabH4bHbcgxFRF5wHC28RFiYKhHuDO5/pK++JCKEwz6Fiz0JeICatgs92YPRFEVAEFAFFQBFQBBQBRUARiEkIeCUsOyYNUPuiCCgCioAioAjEFARI67QjYPOGa1ev4sBzu5yUMIUXX3oFQVufKWnS+WU8evjgfk87nDaDXyaR+DgU1nWFipcuR7SKp23HhvrZcubJlzhJkqRBAVs3xYbxRNMYzC58HNqkLzKObbqDeDSEBGmhEN7Gwc3zClGB43unGM530j2hV8ExogvSi+HAJ8qAaA2iMExu/9iw09yIZkNWILQMecMrJUCMKAowg8gAM35jhNjPP29/NboW9o9R+mJEwcGefqCbQXQHc4tBrNAPCAz6lkBIi9AUVfaImyjtjDamCCgCioAioAgoAoqAIqAIKAIRR0AJi4hjp1cqAoqAIhDnEcBxiuaArwKRVZy/T6rvzyR/9rm8oj3gSToo07drV//9N1HixDhAfaZkyJQlm6eERSJZUC+9kjJVWIRF/ddatvltyrwVQ8ZPm+8zYERhR9GvoLmgwM0bo7DZuNYUjnN217PjHpKBKCCTzojICSIk0LBApwGDpMDRzTOIox7nPKmhcIxzHQ76M2I484lC4O9rjpMGip38sYWwgLTB6c/YIQwhdCACeKWgV8FxiAxEyM1xroHkAZ8oER93orEB5hATEBYQFZBFaGtAoHBv5oq5hnjBqMNnLKGduHio22Efj74oAoqAIqAIKAKKgCKgCCgCikA0IKCERTSArrdUBBQBRSC2IPDFtz/+3K3fkFG+OJ5aDZu+MWnBmoD48RPgtPR6KVKybAXS+Wxcs3yJpzeTrEo3EOz29Lroqg+mqdOm9zt66MA+T/rANdQ/EUaExQsvvUzefNvhg/v2eNJ2bKmLlglptvbtDt4RW8YUTeMIFcG2G98BOLgReg+0H8P5DjGBY5t1aSIucNAjJA9JgeMehzj1iNSgHaIx0MTAOY9sgs88t+HMA6QLYzaEjIlSgZhBz8KkYeJ9bjtePKuQBuh5UB984nkBE6tuBf00KW/pK+QEc0e6KuaFPmWzv5o0YNQxacHCgUFPKwKKgCKgCCgCioAioAgoAoqAtxFQDQtvI6ztKwKKgCIQSxFImDBRoiq1GzSePWXC7744xFqvvt7ioHh97969gxPO66Vo6XKVbly/fi14+7bNnt6MSJY7PiRCnc4vUxbImZBD+/d6MtY06TNkpP7xI4ddpoQaM2RAn5WL5s3yNHrDk37E5Lq5/QsW2RO0IwAtlJjcTx/oG05qSAuIBTbw8D0A6YDxGW0K0jwFiU0VqyhG5MB6MSIyiDZgNz9Ob3bps4uf6AsIC6OP8SCWRFcY0gW8IAF22XHys2NBFArPLingIAUgByB8eP5NiiawYc2CuzfWriFMSNEFKWHSUDGfEBbMDzpA9M8IgpsIDMgKDLKDvtn1ueXdf8cQ6Q79oEURUAQUAUVAEVAEFAFFQBFQBLyPgBIW3sdY76AIKAKKQKxEgNQ0yZ5+Jvm2TetW+9oAiQAoVLxUuRmTxj2x6JBipcpX2r5147qIOJqTJnv66evXrrFL2SdKrnz5C9HRkIOPExYvvpwiZcrUadK9Iv97OUWq1M+98OJLpMt65tlnn8uSPVcervuq109D70tJkCABvFgiXkItUcJE/xPX4XstGla/c+c2jtM4VZIkTZosU5bsOSeN/fWXODVw7wwW57tJDWX0GYgW4DiRQRikBOsMUoM0UU/bDeKCunzGIU8dxKYhK4zYdGwhK6zo4/zH8U9kSWoxtDsgZyAEiFYh2oT0WXxXEZkCcREiBpkBqWEIC2ubUfme/kE8mSgL3hMRQ5+JqkDXgsgkSKhcYqQEZM6Yc/pHv8/Z+0m/HhJPUdlJbUsRUAQUAUVAEVAEFAFFQBFQBMJGQAkLXSGKgCKgCMQxBHDWhxVVgI5A1hy58hINQASCK3iMczkocEu44r8QG6LDgDPLo0IaJHbqR8TJH9aN0N3AEx4U+GSEi9Fl8MuSLcecaZPGewSAvbL49F85e+bUyfCuDW9ucXiTXgoyILy2InM+R578BZkzmfZnG7Vo8y7aHZmz5cztlzlrdtaCtW36wtr498rlS9S/LZEkaHYIH3ELUkI+3uI9b+5IYfPzwb3O1+VTUiBEzp4+iQ5BlBZvtm3taLz48ePfv3fvnnWLtzmfI7d/AZ6HnQGqXxEFk2tSQrGzHmc7fxOzO99ESODshoyAlICMwJltojJwZOOs55wRmYbA4DhtoVsRBV2MUU2AFxgROUHap4tiPGeQABAEkDu8BwOiGFLY66K1YrA0It0mFVNUDdCATf/oB98xJmIGsgTCwhBJEBjZxUhbxfxuFTNRH+gxHbWPi3XAdbRzx/48PtQiiYXzG1Vzoe0oAoqAIqAIKAKKgCKgCCgCioAioAgoAopAXEUgRao0ab/p+/OvCzfvOb561/FLIyfPXf72x192xSntDJOK1es0mLx4/Y6AY1ceTF22KThlmrSkO3mklChbseqKnUfOUwejvlVUu37TFq2H/DF9wcDRf82avmLrnm1HL9/vN2L839gPw36f/GXPfr8kTZYMJ97DwvUbD569WapClRocxOHa8p0PPxs3c+n60dMWri5XpWZdx348+9zzL3T9YfDItXtO/su1bT/4vItjnTfavfcJzvCw5l8CE3BOhRac5r+Mmzpv0JjJs8dMW7SG8YEZff9x+LgpPQYMG4NT3RvrqVrdRq9xP//CxUpGpP1564NDwhKZdmduue/stTsOfti5Rx/Th/JVa9UbNmHmognzVm1xhrGnfSV1Ve1Gr7ecv2HXEbOGth65dI+1MuC3CdM//LJ773pN3mjFOgNrCax43qrN8fPYKXP+nLvSZcqsFu3e70i72XPny++sb6+1eueDjQfOPKL3QXoq1ubKoKMXZqzctrdAkRKlzbUQJO936vr9gk27j81Zt/NQzrz+BV2N2Zttc08IwKF/zli45fCFOzyDYORszTP+tBkyZvZ0brT+owjYRZYTy+vTYonE0om9bH//grxmEysrVkgslVhRsRJiKcWSimUVyyT2kt1oIz76DAhC+3pxFLWWz2hPgE8pOyZ55PVVsS/E+omNFBsg9qnYm2Kfi/UXqylWXCyHHcfn5DXSukGW/oH3U3bsk8jr8/b7cD/mr6IYc1td7EOxrmId7f38xt7Xr+S1tf3Y2/a6zH9msRT0V4z7hM4tpkURUAQUAUVAEVAEFAFFQBFQBLyHgIpuew9bbVkRUAQUAa8hkK9Q0RKQCRWq1a4/a8qfY4f269kVAqP9p1/1SJrsmYdOetOBt9p/3Kn/yD+n3ZC0QpPGjBiMw/OdTzp3s3YQZ/N3A0f8zs74ET/17rF84ZwZWXPkzvtlz/4P089wX9kAngA9BdL5XLl08ULKNOnS4xQmgiBt+ozkCH+k0AbRDOLkecA9hv05Y9EnX/f88XkRT86dr0Dhxg6kA6mCxs9evrF6vcavz5k6Ydxeydff9klDFgAAIABJREFU/rMu36ZKmy6DaZhIgnc7dukhfMQju/WtN27w+pttV+86cdkQKDi52d3Prv2XXkmRkigToknAIoPs/PfLlDW7NBtpR5qzSS9UvGTZmzduXA8O9Fy/gj6mkBRKrqJd3Jlb+gQJJJrWD+cH8uCnURNnZMuZxz9VmnQZ3urwcaeICpDjbP/iu36DF2/d/893P434HTJs0expk9s3q1e1bO50zzcoXyhHx7bNGvzcp3vnmZP/GLN+1bJFjEeCKi6yLgxmWXPmznckDKHuM6dPhUZOWMdhxTtfwaLFJQjjtmmT9Tpx/uqt5avVqsf9IM/6DB0zifRSOfL4F5iyeMOOek3faLVl/ZoVL7+SItVHnb/t6+qh9WbbhUuUKc+aZw1OGD1s0E0Jb/qq98Bhjn3J7V+oyOWLF86Lxgfi0FoigYAQZUQMsHs+NCJCjB31pCxilz7HiBIgqokICr4XSPvEZ15JPUQ0BhEDph2TXioSvYrRlzI+fjdgjN9fjO9kIi7Q+yDKgegGtCPAjnrgyb9HRGOQVgu8wC8qI7zM9wdzxnzSNpERZo5IAcXcMndEwTCXiKSjw8EckhoK8j6J/Vr+TaEOpCARF+hhQMJzTH83CQhaFAFFQBFQBBQBRUARUAQUAUVAEVAEFAFFQBF4BAHxLWckouKvhWsDSX9jTv42Zd4KdpA7wsUuenZl40gmrQ3n+/36x9TJi9Ztt9Zllz71atRv3Mwc7yBEQbuPvvjGsU3S1rCTveM33/cLb3o+79534KZD524R7TBw9KSZW0Mu3m3etsPH7KwnGgSHvGkDhzmO2zW7/7mCQ5njEB70i/6ZekQqcCxrzjzkIH+sQG5s2H/6+qzVgYjAPlZGTJy1hKiC8PoeVeeJaGF+ItJe0dLlKzHWWq++1iKic8t1kFu0w859E6nQc+Cv45gDol6IdvC0fwWLlizDuGgXrFt1+OSLJi3bdeCzmT932+T+XOdsvZk2KtWo25A6kGPO2mVNmznn2VgScOAUxhqi/rhZyzZwfd3Gzd9ijfX+ZfQEQ2gR2QEJ6Kq/3mo7tbAvRH/QPqQS9yeag346zgljCyvSxl2std5/CNh35ieUVwjVZ+y76dlRTxQA0Rfs2OczRiRFMjGiK5KLPWt/pQ5txKod+CaSwP5KdAV4pBerJ9ZCrJlYFzEiK8aIfSc2RKydWD4xIhmGifW2X5PTjhPRELT3MFqBe3haHPpnsGceiYAhMqK0WGEx7ltSrIBYQ7FO9r41kde6Yh+L9RJrIFZb7B2x5mJNxd4QqyRGtAZrgPkP7bun/dX6ioAioAgoAoqAIqAIKAKKgCLgPgK6U8h9rLSmIqAIKALRjgBO/u79h46W4IA7Hd5oWP382dPkVrfhdGY3+crF82ZZO4mYMWmj9gbvCPy20wftjHaBBDokvXv3HrtfHxaIED6cOnGcHN6hZWi/77uOHNT3O8eBk84nYaLEiYO3B4Tr9C9Wpnzl7Vs2rqv9arOWZSvXqNPlo3Yt/vxt6EBx+jxAJ+OWhB6Y9lu+++FnefIXKtrj8/fa7AnaHsBxojJ4vSehH6ZeoeKlyyFCfXDvLsRTHyvtPuz0NUTItAljRzo7nyNv/oLB27eF2/eomPBnn3/hxYwilAwGEWmvcInS5bluq0QBRHRuuY55uC0CFldFL+Kjr77t+/f4UcO//vjtlswBmglEO7jbP9YVBNioqQtWJRcn+2dvv/Fq/XIFs48Z+lPfTNmy5yIKgDXnbnvUy2InFfbt2vkIkWZtI2fe/IXQuzjiRMwbEo1ImX+OHQnhmi++/eFnCIBPWr9Wb/+eYISAbSaC5Ou+g0YsnPX3pK8+aNPciJmnFObgvAiFOOuzN9v+uu/PI+jXJ21ery9TcIH783w6rnkwJ5IpePtWlymzPMFb60pIwP9HWfDdwu57EwHA38cJxdhZjzedqAB28Jtd/Hxmdz66Flx3R9oKFdlG2yCW6RsYvQkzZp4RohUQ1DZkMzjwXYzm0QkxIhpOi4ErOBLZReQK0Q9ga0TOI7wMDc72V+bIsB688m9K6LyIET2RxX5vP3kl8oJ5JT1fWbFUYhD/RcQQEufabfYxICZOBEkeMa4lWoS+Q1BBvISmh4oI4RLhgeuFioAioAgoAoqAIqAIKAKKQBxAQEW348Ak6xAVAUUg9iDA7nXSx3z5XuvXDVnB6IqWKleRNDeb161abh3tm+9+9PkLknrp49ZN65IKiXM4X7OIqPaG1csXW+saZ2motkU4LlFIBa7duW3ThrDQfU7UoiE3Jo8bOfSDL7v1Gjts4A8LZv490dk1OJdbv/dp57XLF89fPGf6FFMnuz3SYv/u/5zOFP9CxUri2HYmHg3xUqdxszdJ+US6LMd7kRaInes7t20Os+9RtWryFy5eCqIpcMuGtRFpk8iIEHHQn/rn+LGIzi3XQfIECmnSqccPg3YGbNnYp+vnH0SkP8znL+Onzn/2uRde6PVVxw5TJ4z5FcLDtFWsVPlKrEMIKU/aNyLu+3cHuYxyyFuwSPGggC2bnLWdXhS9ST22J3hHQMFipcpWqd2g8bD+vboxVvpBdJFkLMNxaeNYry4dO5h2IJV4To6HHHKaaslbbRcvU6EKES+DenX94sSxI4f/f83nK/DP8aMh14RdMsdy+RcszHsh2pSw8GRhhVMXkkGKSVFkUgrhVDei3DflPceN4LY5Hrq+7ddHYY9iXFOME9KC8UOkQeoQ2YYzH+c/5/g9AeFNXUgMXiEFSK90TgyCg/RRvCfFFmRCVBf6wdwwXxALaDmlsfeByKWcYrzSJ8bAK9fQH/qPYDj9Y0wc4xzpoiBdIGcYE88j7424OmOwkiVRPSZtTxFQBBQBRUARUAQUAUVAEYiTCGiERZycdh20IqAI+CICEBLtPu70zbqVSxeyO9w6hpLlK1fHeW/dxU+EQZM323VYvXThXOO05RrS4aATMefvieOsbWxau3IpnrsylarXCg8fHMLnzpw6iVM1rLqG2CCyQnavnx4uDmRX9V99o/U7pI1Cj8PUYQwt3/7g020b166y3iufOK7373Hu2H77ky+7smN94+oVSy6cO3vG8X70nWPbt0Ys4iE8bBzP5y9SHJHaBzu2blrv6bWIQOPId5xvT+eWtEcQDZA12XPnzU8EC1olnvYHvQ+E0olEaFqtZP4p438bZiUrWFeka9q0dtUyT9vOKiTavxLm4WpNkbYqT/7CRXdsc45j5uz/CaYTmfPBF916HT18cP+YIQMeCoyLhkkBNEzQEvlaonys4y9SsmwFrg10sSa81XbLdz/67NKF8+cmiq6MwQv8Kteo9+qcvyc88nzmEr0X6rgT1eQp9nG9PqSDYGC0KHCm4/Rmpz1RFIbE4Hm5K3XvEZlhIirALpZFVLhaDibiBCICMoBooH1iOPDRjCDK4hAYiUEGEJkApjj+IRAgC9KK0Y43iplD7s975g6iBKL7uBiEIFEgRBASCcIcQ0wQEQIJuEmMuYfU5N8IzjH3kDT8O0JkCW0zfsYABrzqbylvzKa2qQgoAoqAIqAIKAKKgCIQpxHQCIs4Pf06eEVAEfAlBKrVe/W1F0Ut+neJUnDsd6kKVWsgKozD15yrUK1WfdLITBoz/KEzFGLjy579fpk9ZcLvjtEY7OAn6qJi9doNnn/xpZcvnj+HMKnTgnZBwKb1a8LDL1uuvAiz2iTdTrrP323Z+LaIdbu6BiKFqIddO/5LM0UqqB+Hj5+CFsGn7Zo3NNeR85/Ijf27dz2MuDDnZJN99toN/9N6gKhxdi/6DpERlrhzeOPy5DwRFqQwMhEsnlxLRA2EgCO55Onckm6JKA/m4a/ffx1CxIYn/TB1P+vW5ydSLrV+tXpZ0ks5tlG0dLlKHNu0dsVST9tnrYSVRgriBuKFKBFnbUvWLdK22ITXSwhJxJoxUUUcL1+1Zl1ex40Y1O/k8WNHrG2ULFepGp8DNq5b/aTahtwpVrp8ZZ5nkxaN6CA0Ko4cPrCPaCRrX3L7Fyxy9vTJfyAKPcVW67uFAE5uIoWs+gTG+e1RtJBbd/OtSiYtFk58HPUHxIhIgISApCB6AYFqoiuIXoAQIFqJKAyiFqgLUWAiFYjWeBiVFYVQQJBANNE2r4aUJT0Vn0l7B8EAKUEaKEgNUg/y3cFvIsgJBMSriM0W4zqExBHgZtwrxSBneAZZJ0RjcE8srq+RKJxGbUoRUAQUAUVAEVAEFAFFIK4joLuC4voK0PErAoqAzyDweqt3PyBdjkRCPLJ7nR3ZODodNRJKlKtU9fy5M6c3rFmxBOKiY9de/Qf//vfczbL7HT0LZwPHScru/WZt2n/kChgcrYhab9vk3Llrvc6IHeMgXzpv5lRXbdJehkxZss2d9tcf1CHF1V8L1wUWKVmmwqftmjU0GgScM7vdnelXvPNJ527sxKeeqwgKnNkBm8MnW6JiYRAVk8u/QGFXO/fDugfREHUaNXtz6fxZ0ySQBafgw+Lp3Jp5IKpg7NCBfSM6tqw5c+fdIloazsgK2ixeukLl0ydPHPeUDGLOiPzYG7zTpe4FGi1hRapAeHDvKrUaNIb0WrZg9nTrOKvVbfQa0RUTRg//2XqceyNMzxpzFd3hjbbRFCFNFWueNG2vNm/19l+L1oWOv0PzBtXQFrH2M1feAoUMmRfR+dPrXCNg0UQwWhS8PhJNYY/EiIswWnUsIB1w2GcTQ5sCZz9O/QRiRFn4iRUQg5wmhRKaNBAYFEgDbwpWm/RMpD+kL5ALpKqCoCC9E/2FeCDaAtIFcoUoCupAthBtAbHyvBgkDJ9fEUPvgjRYkLRcY3Q4IDl4Hx8hbtW0sM+yvigCioAioAgoAoqAIqAIKAKRREAJi0gCqJcrAoqAIvAkEEBsl5Qw0yeNG+V4vzIVq4WmcHJ00JP6KChg6yYEqOdv3HXk9VbvfDDipz49PmzVpA76Ds76vWnNiqWkX2r65tvvsZvdWR10BELv54Ymg5ALobve/xo74pewNA1MmqYbooCMkPOISbOXsuu8ea3yRRy1NkhtRJshhx6NEoC4qVqnYdPjRw4fxDG9z4kWAloFYLl9c8T0JDyda5zw6CqI7kKojoInpeM3vfpTf/iA3t0dr/N0bo0+xIpFc2c6amF41Ke2zRo4E2E3bRBhASHmSZvUzZg5Ww6Isj2S78jVtfkKFClOFJFobuMwfayQJuzCuXNnSlesWnNY/+8fST0G2QEhtnzhnBkIglsvRhOGiCKwcXlvL7TNHEIo5siTr8DMVQH7vu4zaMS6FUsWvl69dEGIF2tf0HeB1Nu9cztiwFFSAo5d8abjOEr6qI3EGAQggfn34CUxIhNw3Bs9CtIsQQ7y3BNpQD0iFSAGiFYgHRSRFryH1IBM8DgdnQdIGNKCvnAfSBOjbcEr6Z+miUGOQwrmF4N4wHbbXxlnCTH+/WK8/HtpIkIYH6mtsovxbxHvGStj099VHkyUVlUEFAFFQBFQBBQBRUARUARcIaApoXRtKAKKgCLgAwiUqlClBt105lStUb9JM85ZIyxIoySZkzJhpeXaBbOmThouTlzHnfrOhj5qcL9eQ/6YvqBe0xatJzrsRqc+jmF2f+/dFcTOWZcFHYmMQiKQlmf+jCkTwqpL2iTO9xgwbAx97Naxfas50yaNt+ojmOuJJrkmXmtHfYp3P/myGzvQb0rnzpz654Sza+k77URUANvTpWLInR0eCnw3btG2fbkqNeqMH/nLgEP79+yy3jcic4vIOm04EyH3ZExhpWyCMHo5RarUGyOQDgqnPf3YG7TDJWHhX7hYScfoItN30oSBy/OinC3SJgFrli2aZx1XfVnLfF40e9pkx/FWrd2gCceWzpvlNALIW22z5knx1nPQyPFEK7Hmt25YQ8qZx4rob+BUFX2OwEgTFkJU4FTF0fqcvGeXOQ5enM9GXNmkt3kkxU2BdMgSaImDCBgxayILWCcQD6whSDWEtFOJmZRLaDqQlhBSAgc/zvzqYhzne4yUUoasMFEbUQKpg44I/Dj3h6yAlOC+ECdEXdBX+g8pQUorxmNIFMhQPhMxwjnqcIxridJgcwDkc3oxCAqMyAzGgs4F94oyEe6cefMX2r0zcKunABFRCTGvEVmPIyfQED1jk+yZpAeLskK6RXS6rGkIo6xxh4aIyJOMmclckffeum9sbZfNOXduy3/yt2psHaOOy/cRkD9vX3Gmy+f7I9MRKAKKgCLgGgHdCaSrQxFQBBQBH0DAv1CxEuTdd8y9T7RB5mzZcyHceyzkEM7H0CJ+YxxFtrlTJ42vXTpfZkSG3SEruAZRb5zkxsnrCA9O+N07A7Y6IwSsdTNly5HLiF+Hp9+QIlWatIzhs7ffeLVemfxZcay7av9lSUl18sQx0nY8LFlz5slXtc6rTYeJYDfOXVcEAX3nR2lYqYeicjnkK1g0lNwhMsDddgsVL13us269BpCi6Je+33ZxvC4ic0tKI/RN1q1YutDdfnhar3iZCuR9t21as9Jj/QrmDH2TQwf2ssP5sYJmCSmyXBFNeQVnLiK90+gh/XtbG0ALRSJvmkjwzlXWtvUcjp9KNeo25NlwRcZ4q23WfPD2bZtb1KlQrI1ogrgiK+hv9lx5QwmLKFy36A2wcxxD8wWNmCJipcX8xMz5FPIeSwzRIWZzZZ6uF63vUwhAYkEA4IzntwNRBnzm3xyc+xDqPIP8u2NIDFJG4fDHcOYj0A1xQX2c/N4uRpOEvkNUIJqNrgYkBk7rCmJERkAy8L2DZhNjQJeCY5AQpLXiGvrM2HhOeF54bogagcQhzRXjgdQgEoXrIh29RETlhHmrthAB5ilQP42aOKPNB5995el1caF+719GT+jef+hoV2MtW7l67ZVBRy8Q1eYuHvyd8/fSTcGNW7Zp7+41kan3Rtv3PlkacOAUDszItBPd10LWo10W3f3oO/T3v8bNWrohuvvh6f35+2XSgjUBlWrWe9XTa7W+awS69B44/NOuvQfEJIzQMFuy7cCpvAUKF4tJ/dK+KAKKgCLgbQSUsPA2wtq+IqAIKAJRgAA75J2lOGryZtsOsqnv5E6HlEPyW5tdorb5M6dMPHXi+CPOfXe6g8gzTm6cqo710UPYtSP8XZ85cv+3a95RS8DZ/ekvTmP0Gu5LCauPL778SorzZ07jfHpYPvm6549EmBw9fHA/u0ut5I21XjYhNg7u3R0clvi3O/i4WyeP/Lhwh9wx7RUoUqL0z2OnzIHgQTTamVaEp3NLhAC7ShEhd5UKzN3xhFVPCIvKEF1Et3janp+khCKVFxobzq41kTGuUnn5S8onrjtx7MjhZbKGrG2gT5Hs6WeSr1oyf7YjnjgDIUMcr7Fe7422SROWJGnSZAjfBwVu3RQeXoZwikw6r4drLF1yni8czWDN7njS96QWwymLQ5lc/W+LdRKrL0Z0CmQUzjF/MXaX8/2C05od5pF2zoY3fj0frQiYyBv0IHDws0YgAHD8E3ZzQQxnv3UdoPnAGjkmxk52CFvWHeuFdWe0H7y9dug792PnNMZn7s2xvWKksoKQMJESEBnUIwUUESSkj0Kvg2MQEpB3RgODf4NMpDrtQXQwHo5FelyksZN2bCZdIu/dKeji5PYvVAS9K3fqx6U6YJNf/o29esV5WkGwKF6mYpWn5d8LRw2hsHAiQjCZXBRWu1GJM05LSJLr167yHPpkYQNCrYZN37gn/+hH9wDAU/axQE76VCGVJps9SGnpUx2P4Z2tLATQyylT8jdRjClEGEsU4f8ksIp/f7QoAoqAIhBnENCUUHFmqnWgioAi4MsIpEqTPkOAg8g1KXiy5czrL7+tn3UkLJLbdwdG9EdYoF3jAaLEmk8fwW3u55imyBm2OfL4hxIWkpd/QXjY01/y+YdXj/OE7589ffIfU7dMpWq12N3/Zv3KJTNmzY5Qqs1RA8DUzZQ1Ry5HrNy5Z0TqoJdBSi50E9y5vlGLNu9+3r3PQCIh3m5au6Ir0sXTuTXzsHb5ovnu9CMidYhswPk/868/xkTketKXHHYRXUF7EmFUkvXhKkrIpN6aMXHcKEfCq2L1Og1oY8ncGX879q18lZp1ObZy8fzZrvrtjbb/fw5vueUkIVrp0L5HU4NFBGfLNegO7BdjRzivOJ5x1vIKcYGDFicIDl4c1UR4sPsccoNz7JrHYcvu8rVi5yTyAl0DHNfsOscJ9QjxqCmlIjlj0Xe5iRhgTkmPxJzjvIf0gvAi3RzOepz+rB2IDNYNZMURMaJ1IMGIsODaQ2JRmjrJGTQOKaLuS4oo1jp9pK8YRL6fGMQb/eUY5AREBREU9BWSjp3268XKibGmuY5xU2gTUp91T7osQ8bEQ4Bb+hAm+e6s3+YY0Xm8N4RpWHWt5zJkypqdqDJNB/U4YkSk8vdDWH8DoDslvPdBTzY1sDGBuz2pvy2IKCVqE60ud9dFTKvHjnH6ZE1lGh19JI0lf6sFTZ/8Z3TcPzL3zF+0BBGRtsP7nUemRqbtuHotv6vYxHJ4/z6n0b7RhYtJC+ps41p09UnvqwgoAorAk0BACYsngbLeQxFQBBSBSCLAj+y7d+4+IpT9ebc+P21cs3xJ/iLFS+3YtgmHSmhKHFIpyc47nEa2RIkTh5t6g93e2XLl8bfu9P6f7ETketnw/sg9U6dL78fx82f/P8KBHfxyy7uOJAE//Il4cEUeWCGhv9LVcPvKNQllULdu3sSZZGNX45c9+/8yb9pff+wUnYjX3nr7fY6fOfnPI6LF5l4IF1t1QNh5nya9X8Z9u3aGqccRkekzP8h37wgIMwd52gwZMxMhgmMdoqjz+61fD2snvSdzS7+ZB143r1u9PCLjcOcaxgqWG1YvW+xOfWsddo0JH5eRCAhX10Ia7Nj63xp3LEQq5MzjX5DjC2b9Pcl6nl2oJctXroZjZ83yxY8RNqWF7EIPxVGw3rThrbavX/vX/ny6t+ZTpE6Tbq2T/nuKtakv5AGO1NBnSAqEBamecEzj0CXVD05coilwwPIsgS/nuC6zGOQipAXpf9iJCFHI35SMi/Q/aJGssb9nh/11ad9pbn8lMiI6i0/sOjNvEFeQWqwJNIcg2/jOZt7Z6Z1OjLkmwgpiC2c/Dn3q49CHDGO9cB5NiUhHIXiCgHzN3EPYwt5fXtHawELEIGIgWOhbYTGiGyDgIC4YN+OCkODZgKCpaL+Otc+aXyHGmg8U47mCkOF+fL09ogXjbp/5ToV8JdKCyIDwIg9Nu0YPKHh7wBZ37xVX6uXOX6goYw0K3IwOidNCNJsrrSRX1+TJX7goehIhB/ft8TaW/JvE3wyz/57wu7fv5c32c+UrWPji+XNn3U1V6q2+8Lcvbe+SNKfeuoe32vUvWLQE32lhaYt5696xtV0wZWx7gra71FOLjrFLdLj/P/KwkDo3Ou6v91QEFAFFILoQ0JRQ0YW83lcRUAQUAQ8QQCDSkAVc1vaDz7sQ6XDm1MkTODKCAjZvrN3o9ZZrd/9zhZRNEAXUyyLvrbdBsLpTjx8GGRFvzr36Rqt3xs1atqFoqXI4YWwQGK3f6/glKRGCArY8kq4mniTNpU6SpE/j0LRxr4kL1mx7vfW7HzoOh3uTDsmdYR45dGAfKQK4t6mPk4aUAd36DRllbeOGiBHwmfPdfhwyCqHlQb27fcmxZ5I/R15xpxEW1H9KmBgJqQ7tOw72kZPnLuv6w+CRpj12YCZIkJCUJ5EupOWgEVc7XXFEkSt3+ootu4uVrlB56I89v2nbpGb58NL+eDK3oXMkuzEhmKxRKZEenEMDxaX/pJsKS4fB1T2ZBzB3JSbIubwFihRztXuVNFrkcoZwI62U9T44I2h/3colC28Ja2E9Z8TLRdR2m6tUVN5qGz2Nc/LwOj6fEHCt5Nl7q/3HpGN6WEhRgnMnqufNoT0cq0YsGQcuhAPPPyTUULHfxCCVFomNFSOlDs8rZAW70HFe45AmfVRnMfLE/yzWS4xIFnaMszMf4sOkBHqoieHlsWnzEUfApDnie9PMM8QFhBXrhdRDCGrzmwKyCg0bXo12BI4fohL43iZ9lFV0+4mSFnJv1jhEBIQbESJEB80SI/UT/ScSJIcY+husV0gXSAucREPsxvdIRjE0MBg/48Tp2UgMMXuwYY1TIjQ+Uvjx7yHkOv/O8x1uby/cFyLq+K63bioI96I4UiGPEBb8OyDBCU7TZfH3EXgfEP0oTyCh3eDArZvthJgnl3pcF0KFP2WCA7exZn225M5fsMiTikgJCyQTgeqLeBLZQySuiq9H3WNgoqViUoQaG9EkcC4n3zFRN1JtSRFQBBQB30BAIyx8Y560l4qAIhDHEdi8duWyCtVq12/9/qedcWSwG79ZjTKF2nz4eRdSA7wpDk5IjPG/Du7PZ0iM3Tu3b3vznQ8/OyUC1ewwL1e1Zt2aDZo0x1k646/xD0Un1yxbNO/Tb3r17zt07F/k1M/lX7AwP9x/7P7Fx+w+t0KPs5wf5c3bdvg4Q6Ys2YhokM3iV34fPuhHa72UadKmx+kSKLoS7kzdAtHaqF6v0euQB/Om//VnhsxZszd+o827pHiy9pW2+IFGCqgRk2YvJQ1Rt47tWxlnPJEh9E+GGLqD3VrAhFQPFarXri+kwNEqteo3JtXOO03rVKLegN8mzihXpUYdoi2a1SpX2JUT29V4cDYPHjd13uolC+Zs3bh2VeHipcqZlA0IqIIH98uR279AweKlyoLx5YsXzk8cM2LwmCED+rjrkA45KPH/bs4tfcXB4e48uDNXzuoUK1O+MkLnrC1P23g6eXLSyNhc7Rwj+oIUJ2iTTJi3euvwAd93WyUYm/uQ25f3c6dOHO94b+OMQL/D8dwr9hzFIQdc74r1ZtvzZ/49sXmbDh9DULBDsoCkd2jUvPU7rJMen7/f1tpfkTQ5zzO/ctG8WTwTPH9zJapo9C+PCox7ir21vpNIBxwU9X/kAAAgAElEQVSxJqXNBYmQwNlMWp9VYjhizXtSR0FEQI7i9K0uRpoco3WBs7W2GDvySeWG4QCGEMGZTWopnMgRTp8TmXHrtW4hQGQBUQbkzyZ6YoUYqZ5wzmM49Zlfs/uTaAuj+QBRQaql82IQBjzvfE88Er3nVi8iWYloBymMhfUGqUAECOsOvQ1IB/rGedJWsZ55b0iJNPYxQoqzziFeqEdUBlFHEIpgwHmjmRGhMZrovCnjfhsGmV1I/i1xdxd19lx588ckZ1skpyxKL0cLiX87Xf3bnjNfgULcUKSY3CYsEOfmb7LFc6dPidLOumjMRBPu2rHNZyNoIFz4O8jx78YngZ/jPcBTpED+PXJoPwS8zxQ2YvA3+AL5O8JnOu0DHZXv3sL8nvDmBh9PYUCrhMjy4O2+TVJ6Om6trwgoAoqAIqAIKAKKgCLgIwiQdmnmqoB9pFVZsSPknHGkTlqwJmBryMW7HEPLwTocxDrX7T11lWuwNRJ98cV3/Qazs9xx2ERnmLqTF63bXrlWfXaLOi0dv/m+n2kTBzLpCRwr0pcthy/cgbhwB2LyZgwcPWmmaZfXP+as2FRJxO8cryc6ZNvRy/e3Hrl0DwLHer7B62+25VqTGsrxWtrbePDsTeos3rrvHxNpwv3NcdqVoA121npUSD/0dZ9BI1bsPHLeOg7rezABX4iZspWr1+Yaj25ir+zu3EKigBVkUETu4841kAmbDp271e6jL75xp75jHXIGgxGpzZxdz45XMzdD/pi+AOLCWm/ExFlLFm7ec5x+OF7f/tOvemw+fP62s/kkPRj3bdjsrXau+u3NtunT7DXbD5j1wXP806iJM0SWJjS9lbXUf61lG86bunwXGDImIphH5Bq598NoCIf3/5PP8cSeEUst1kCsm9ivYrPFxokdtTwHx+X9abHLYpvtdb6W12xiScXii9HmI/eLSJ/1mogjQPYku+Hljy/2jFgWsYpiZcWGic0RGy02QuxbsVL28+3l9XuxfmK97McayWtlMX+xlGKJSZlk7hPxnnp+pf2+6Ewks/elsLxWFWssVlrsPbHJYgvF+osNFZshNl9svdhGMXbUrxHbInZEbJVYa7G2YnXF0oglFPM4mp3NB/w7RCrIIeOnze8/8s9p7o5y+fbDZ9/++Muu7taPK/XAku/Qjl179Xc15g+/7N6b7ykICHdxkZSD1bmGzQ7uXhOZet37Dx3Nv7fWaNTItBcd1xKZC2aOf7NGR1/mrNt5aNTf81dGx70jc08264BhszbtP4pMO3rt/yNANC/P1oDfJkyPSbjUqN+4GXPNnMekfmlfFAFFQBFQBBQBRUARUAQUgYcI8Md0zrz5CxmHbaUadRvijCWdE2LYzqBCTJAf1AWLlixD7uOw4KR96rsDOU5khOlc1YVgiciPUcbHdYgwh9UPzqdIlYZd3I8U+jRozOTZrpzfVGanEqQNu/ysF4NRS4lIgUhwBwNXdSA//CRCxDigIUVI/5QxS/acidzU6XDn/u7MLYQIDnn65E6bEamDGCBEDOm0InI94e6s0bCuJSVKluy58jirU7pi1Zrg7ewc69TsVnZ2nnXC/V3d25ttc0+eOX6ElihbsWp4JBnioKSoYldlRHD29jUOBMNT8jmRncR4yU5ijJXXIWI/iW0Tu2MhMSBVj4lRB7KjsVhyMdoJJS60PFkEDJGAw10sgdizYn5ilcQgLb4RGyNWx+6k/11ee4h1Fesk9pPYSLE/xN4Rqy6WUyyD2Ati0UZYgKTcH7IE0iKpWCqx3HaDlCkmBunQQay5fTw75BXSYp3YX2IQNifFEPS+LnZH7GexV+3XVrCPFVLEo+9fyPspSzaE7vJv1eGTL9iQ4M53OP8m8kzxvfVkV0vMv1uRkmUrgE3VOg2buOrtsAkzF7Gxwx2sTRuQ4rQb3vd3VCHEhgc2ikRVe9HRTv2mLVqD2YsvvZIiOu5v7kl0DP0Ii8SKzv6Fde8W7d7vSN/52zKm9tHX+sVmETB13AgV3eNgfUJgswEpuvui91cEFAFFQBFQBBQBRUARUATCRAAn5+fd+w40zr6wfoArlNGHwC+SHiqv5BiOvh48uTu7S3Q9uR7pnZ40Ao4REQ6fiZhIIva8WCGx9mIrxG44kBZBls+L5H0NMT8xyA/Ii8ciL5TM8M5Mi5PdRFgY5z7RAhnFiEQoI0a0BFEU5cS+FFspRkQCxEV3MSIuIDA+Eysill4MMiCH2PNitBctERZWxOx9gJB5WYzIj8xiWcWK2vu+TF4DxGaKzRb7U4woC4iLS2K3xcaK7RUjyuITMQiapmKI4hKZwjjdJi2I/jPaTegj8EyQ2i+8mWaX/5N0nofXn5h0Hick2BBZ56pfK4OOXhg1dQEp79wuQ/+csXDu+qDDbl8QiYpstmBzANpXkWgm2i8lEpWoyOjuSLEyFSqzJqrVbfRadPfF0/v3HDRyPBuWWBOeXqv1nSNAJCvrwej5xRSciACatmwzOlFaFAFFQBGIcwh4HKYc5xDSASsCioAiEIMQ4Mf26GkLV6NFMXH0cARtEXX26d12MQjeKO3K+y1frRkTRCWjdFAuGkOL40ncR+8RcxFAAyMMQ7sAsWJ0EPi++lWMSKbCYtXEEPX+QwxBb1MQ754ntkCMFHVGDBnNhEc02JS08Oq6wNGOuDq7oYnA47cDqf5IZ4cWBOLT6MigBUG0EvWZbxySzN1qMTQd0ITIJUZKN6s+ilc772bj6FFcF0suZrQ3WG+kmUOce70YueI3ihHNiCA3ZDSaF+BAdBm4EOnFuiVNIvoX4MBaBRO3CAuiJV96JWUqEVhF8N62a2fgVrSkCpcoXT68sWQXXYDTJ08cv3DuLKLnWiwIoF9x/tyZ0yePHzviDBgJCs2EftCu7QFua0MQiQGhFBSwJXSunBXIfKJhSUkV2QnJkSdfgXjx48f39Vz2RD2iJRIRPKISTxN9Gbzd98SMWQv7RTz+9q2bfAdHqhQqXrocOmuRaiQWXAymQiw/kOfrse+AqFx3nkBFJDjf60H2fw88uVbrKgKKgCIQGxBQwiI2zKKOQRFQBOIEAqRKmjh/zTb5vZqgWa2yha/+e/nylcuXLh4XIek4AYAOUhFQBGILAjhzEV4OFoOk+FDsbbHuYu3FTlsG6ifvSQfWTWyPGA7Hr8UKiLlM5xVbgIoB48DRjtM9iRik0w6xY2IJ7fjjHF8qRt7v7WKQGgixQ1hkFCMFTwMxdAEQpUacmnYgLXDoR2tBiNveAUgVBOARhWfM/EZCGJ71yfrrJPaZWDl7fc4zFgpEDGkM0T4qKmaExmmT1IkQG27pWRgnqnFQ3b937962jetWu7PrF4fbnqCIOYKjdRKewM3zSLRjUMB/JJCzYgS3PXFeZ5BUhGTHFMICIuuxArnw59yVm/v9+sfUOo2avxnZYYqeeqgouCGzIttedFxPRAAaFnuCAj0mLLyBJ5stIvo3NPpb0aElwpojxagzx7qnc0pUwW9T5q1AK8fTa71RP7owZSz+hYqVPHLowD4IYuvYonrdeYJbpqw5cpEKKiKbnyC+n1SqOk/GpHUVAUVAEfAEASUsPEFL6yoCioAiEE0IIKKJNsOaZYvmvdWgail2CbLrZrdGV0TTjOhtFQFFwBMEwonAgMDAiY2jgOiLImJ1xTqLkW4FQdsa9vuxAx7yAocXgqPsik+s6aI8mQ2P6zI3RFFBMkFeMD+1xJgLnPIbxHaLEU0RJEYkDREI+cWIQCBtCWQTaS1oh/l2O+rA4956eIGdtKBPRFn8KwYRQdQFuk9ElhAVAkEG8WAKzu/LYuxwZoym3LGPMZ28FrRfC7kTOt7wUkPl8i9QmF3T+/cEh2pYUDavW7WcXdBh6e1QL4f8TbA3eEegpS/6VhBImSZtevQSwnL058zjz1zZPIleILqCa1ztfkZDiqgNdm2HHNq/N7KTkdu/UJGbN25cP7h/j8+mh0EnAAdwRCIsvIFn8A73I2qs80dEzpTF63eEpZcW2fl2dT26Fey8l+hqt6OBXLVlHNqHD+7j+zlaS3RiSgRUNtFKc4ZpVK87T0DOK5Fh/33HbHZKirpqi+iv0ZLe7rW33n7fk/tpXUVAEVAEYhoCj4TUx7TOaX8UAUVAEVAEbDb0Kpq1af/RrwP7fDusfy8cdTb+GPWXHy3TJowdqRgpAoqAIhCLEGDnPTv42aHPrs/xYjiLcX6XErMKtPe3H6cuO/9x4HAtTmPaeSjYDWGixWMEDKlAJAtpofzETGooIi5w8gMsERU4Vsj/j6MdsoLjzAkRCjnFTtjrE3HA3BCFEO0RFhZErH2BmCEVFKQDqcuIGrEWIjFCndVSIDggZMACnC6JEUlCtAVYLRdjPYIl50PXpauSJ3/honuCdgTcu3sXwiS0CGGxrOM33/fDqe7KoY5jnJSRe4N3KmHhAC6Ofg4FBbpO3ZQ9j38BdtsfCznEvLtVaJd52u0iWuCWsAsNyhXKIbxFAlJ1udVoGJVCUynJvYi6iWxb0XW9IXkiEgkUlXjiqIfImj11wriIYFG17qtN4wnzsnfXTqLKnmgpUKREaW4oGAZE9sZjhgzos3LRvFlHDx/cH9m2Int9dGKar6CQQPHixXOGaVSuO08xQgeP+++T9F+eXAvRkc4vUxb998AT1LSuIqAIxEQElLCIibOifVIEFAFFwI5AozdavwNZMXbYwB8MWcEpwsHJqbp96yZya2tRBBQBRcCnEXBCKOBAxmmLo/uERFBAXqBfQVoUhHP7irHzvYXDwL+Qz+gNsJOfyICY5BT3tTkCOxztkBMmTRKOV0iJfGIpxfg3CAc9n0mdhDMVMgLnPNenFSMSA0IjROyk/ThR3jHJ8UpfIRMYyzl7/y/IK4QL50gVZfK8G/aLdFjsTC4rRpQJaxWSg7RRYIClFgM/1iMRGaxpl2uSXPJzp06CpHtY9olTVLI/XihaunwlV4RF9tz5IPRsGmFhRe6/9zj67bnpNz9+9r8jOXLn8zhPPO0eFE8iUQ+u2kU3w9U5T46TFoYUVGtGDR3oyXUxrS4kz8Xz585GlMCJKjwf6ldEUBugeJkKVQ4f2Ls7OvS7ChQtURrS6uDe3USzRarwXLCGI9VIFF0c3ZgyjH27g5wSUFG17jyFimgaopGsBLY7bRQvUxEtJdu2TeuIetSiCCgCioDPIqApoXx26rTjioAiENsR4Afqx116/kiI8uC+Pb6yjrdU+cqhu4y3b924LrbjoONTBBQBRUAQwLmNI3mhGJFl2cQ+doIMRAbC3s3E2ImKwzg+KaMUxQghAG5EEOCkh6CAeGgohtA2kS9txN4Tg0iCsECoGictUQVEJpQQIyUSx4nSgAQwQrExbU4gLAwxA7EAIUHUDuNPJQYBRnQF65D0ZWhcHBKjEP3DWMEHYoN1R/0XxPi9xZghKlySFekzZs5KpISjjsJ9KVvWr15RrFS5SvZ7PfaCw11Sr18+cewIKdSirJC+J1HiJBAuMbYQcUo/XXVQoCnMDnI0v5zVeTlFqtTsuPckTzz3y54rj39Y17Cx5PkXXyL6KNzCGMLSQ8DRTxqg4DB0OMK9ib0CKW7CqpsmXYaM7NBmLbrbprv1/osSiZjOiid4Mj9hpVBj5zp9DkvXJKwxZZHJjw4h5AQJEiYEw6MSCXT79i3I1cdKsqefcSuckLZMyiF358+b9aILU8aU3x61cmDPrsdIoPDWnbt4O2IX3veWTOOzaFjsDHSukRP2+syZ55/jR0MgB705Z9q2IqAIKALeRkAJC28jrO0rAoqAIhBBBMpXq10f0mLciMH9HVMAlK9euz67bi5dOI/jRIsioAgoAnEJAZy+/BAfIoaY86diiD6bgpPwDbFvxUiRw/k8QlqgSaDFcwSIliBKgggBnPrgCPnA7wjICBygOPeJIoDU4Dy7znGocQ0EBhoXvCfdEqRAjBDddgIF/YJsIdUTJAukAwQYmimkd0LHIr0YhAXrkPOmEFFBJAavRFuwRqkDPsZc6liYdDnOoig2rVm5lHz5rpzaRFgQieFkPLY32r33SaMWbd51ds4c428NZ+e/6fvzryMnz2XcoSVztpy5fxj2++S/Fq4N7PbjL79F1Fnnqi81GzRpPm7Wsg1rdv9zZd764JAvvus3uHTFqjWd1Rd/+gtdfxg8krrr9p682vaDz7s41sMpmMu/YOGwnMuIlXOdSRlVtU7DJsMmzFyEbhg7nJ3dG+FoBKRdtct9x89etgH8wsL9uRdefKl7/6Gj1+09dXXDgTM3vv/5tz+41vEaExGwM+D/c9lnlZz7nXr8MAiMmJew7oPzvtV7Hb9ctGXviY0Hz94c8NuE6TisrdfwGYHwOet2Hho3c+n6JQEHTqGfFla7npzDAUuamj07PRfcdhfPbLny+o+YOGvJpgNnb66XNeEqhz8EEFpw1p3zZStXr92t35BR73X6pifC1taxMU+s+8G//z33p1ETZ0BEMSf9Roz/+8fh46b0Gjzqz/JVa9XzBI/w6nLPDp91+XaUaBFMFr2MDp9//V3u/AWLQCAesGjcWNup3ej1lst3HD5rnkuekS++/fHnifNXbxs4+q9ZON9NfbBhnk10lmN/mr759nutOnxCxOLDwprr/cvoCZ927T0gSdKk4f57yvPDc7RiR8i5ZYGHzvQZMnpi4xZt29NgdGAKWdew2Vvthv45Y+GUJRt28rxBVuYtUKQYv6fOnz0NIf2whLfuIJmXbT90plSFKqEaWzxnLd/58DNwHT1t4epyVWqixfVIced7iwvyCWnI/Y+KEPjXfQaNWBl09MKMldv2Fi1VrqJjm9QjfTDi6axP6iROnCQp6xPrM3TMJMe5DG/96XlFQBFQBGICAkpYxIRZ0D4oAoqAIuAEgQyZsrCD2LZ/d9AjuUv9JC0AOWyXL5wzQ4FTBBQBRSAuIGBEux3Gyi54cs6TJqW5mL/Ya2KkjyK6orwY5EUfMb5HNwhp0VwsqUZcuLVqcJwS2YJzHkICJzwpkBCcJi0U6Z3QrSD/OaLCpJ8gZRSvS8WIKsChf9R+HuIC8oPd8DE1VZc1NRTrC8clZAtrinOM5YgYxAsaFezaZ21xfJkY/y4jisxxfmdB4Jjd/5A8riMBxIl6TcIkjoiDSuo9UjatXbEUR6UrB3p2cbo7y1eOg+7djl16CB/hctd1g9ffbLt614nLCM863pcUVeYYzrcJ81dtxbGb7Jnkyes1bdE6U9b/d4A6XuvJZxx9OA8x0uwM7tO985rlC+fhVHXm9HslZeo042cv31i9XuPX54gOwV7R/Wgvzl10PKz3xaGIozxM/Ypc/6XTgnz4rFufn/oOHfuXCPD6Q5QM/WPGQgS7HccSXkohUu2I7/Nk2gwZM7vCgb5OmLtqS9XaDZvMmTpx/IbVyxdD2JQoW7HqY/cTge8L586eYdc053AmT5y3autrrd75AIxG/T1/pauICNbAgJF/Tvvgi269AjatX7N47vQpFWRDTNW6DZta70M7lWrUbbhswezpaKb9e/nypfafftXD1ZrzZH6pK2upEI7ViIhFu4NnSYk8FpJoY/qMWbL+OXrYoH+OHQ356Kvv+jrDhfkz5A/RGD0H/joOx3q9Jm+0gvjqL3hZx4cgdMo06dLfk9w8L7z4Mvo0NtL0pE7nl5FUXX6Zs+VI9ox7kQ3u4EbkA6Ler7V694NTJ44fvXHt2tV2H3b6Gsc11+/aGQiJ+ljJna9gYbQ17ssuJ8ihSUIsNpV5Fd91Up7bclVq1DEXnTl9CnLVxtgcG2LNfNzlux9av/9pZ3MOQnXs9MVrq9dr9DokKOfDGkuTlu06jJm6cHWa9Bkyjvqlf++Jo4f/XLZyzTqkuTX3fZKY8hwjRP3V9wOGSnDKLaKuGMuvf81ZBvniDNPw1l0ocZkwUSLqyddz0mF/zlj0ydc9f3xeSBAiuxo7EMXufm+Bj3nuOnz29XepZO3NmDRu1EuvpEzVVYhiR1KTe+fMl78Q/eAcKYOvX792NVXa9Bn4Dswo6/PFl1Pwb5EWRUARUAQUAUVAEVAEFAFFIPIIsBtGnGoP2FVpbY2dcVsOX7iTIlUacoNrUQQUAUUgziMg35UIbP9PjPRP6cW+4fvThU2U45XEUlM/zoPnBADxe9jwfYjFE0sullusoVhzsTpircS6inURGyg2QOwLsS/FSopls9dvLK+ZxF4USyr2tBgOHtrmHqEW3cXaF3vf6OPzYnnFSoi9LTZRbKXYUrEDYmfFuon9InZBbL3YGLFhYuD0oVhbsexiL4i9LJaQ9p2Nl125IybNhuhxWhZu3nOc3d+OJ9npz98E9YVAcDznX7hYSZ4BdkY7axSn+Yb9p6/PWh34mOguTq+tRy7dw9GNA3Xz4fO3J8xbvTW1eDhpy910R+7MLZEC245evo+T09QvXKJMefqOU9HaBs5UyAoiK3KIWDbncBxSt2L1Og2sdSEAOG5SADnrCwTF7LU7DuKspi4Oa5x+b7770ed8tjptzfVEdhAVEVbaIXbFs7PZ2T1xMP69dGPQ8u2Hz5IKhzocYy5+mzJvheM1REawQ57jdRs3f4t+sdOdXeo4gPlsdq47XgsJw3mIKc4xNna8g7m17uRF67azg9s4Q/2yZMsx5I/pC8x8uzOPYdUxeEb0b9ew8CR1zvp9p68RnQNBRT/M+nm3Y+fu1n6xGQg8WrR7vyPHvx0wfCzrnP7xLBFlwnlrNIL1eogD1mpURxeZe7CmWVsT5q3aYp4x5oTd8+bfM8bmDGsin36fsWQdu/iJUGJ9mR35PM9WRzfkFO0xz45t0QfOQeJwjrHO37jr6PTlW3ZDeizYtPsY30eu5pu2wajnoJHjTSQP2G6UKCJDujxJTOk/fWfdW0lYnm2DqeM6Mf0La90R1bDp0LlbRKgNHD1p5taQi3ebt+3wMThDgljT6XnyvcW9h0+YuZi+WaOE+N7hWFjkAxvaqANBFdlnVq9XBBQBRSC6EdAIi+ieAb2/IqAIKAIuEFizbNE8cWw8aNa6/UfsEGNnTpfeA4ezM27GX+NHR1S0UAFXBBQBRSCWImCEutnt/r0YpG41sU5i1og0ojCWiJHqpo78uE8hFs9OekB8PLRYipOnw8LBTpQF6TIwRFpxcPOK04q83xwnmgXNBrQWSFtBmiF27Zu0SKRaIk0UkQsxqpCFx2JmHd2WThJFQkRFgNhcMdI9mRRYkF3sWuUzY0O3AgxWiqF9QTQJu5gxxky6KacFZ1b23HnzuxLV5iLSQhUrXaGyYwOS5SUPu8T37tpB+rNHSqHipctdl93ZB/c+npudijhfcapNmzAWXZhHSpGSZSugmxCwef2aPkPGTNy3K2h7uyY1yptd/lGVHx2HKpECo37p12vyuJFDTScQ4SUdJn8LWTvW8t0PP2O3d4/P32uzJ2g78xLq7OeVHfDWurlkx/ndu3fuyPCdpsuibubsOXP/czTk8Kfdeg/4Y+SQn34b/OP3/O21dcMa5tHmzGGP03N3UOA2x3Sd5t70J5NMTHDgNqdC3x91/rYPaZy6fNSuxQH73CDe3bPzx++O//WXAdYxpEyTNj06GxIRsAFyo0ufgcMXzPx74lcftGlOGpvtW/7TMnOMLuEYhBWEBrhOn/j7bxxjbPTvrgNWRAuc/uf4Mc5TL+TAvj3vvdGguplvx/Xh6eecef0Lnjtz6mRE/nYNC09Io16Df/vzzp3btz9p83p9tFzo27aNa1cNH9C7++I5M6ZY+2p0G3YInqQHqtO42Zu9v/70vd+HD/rx9q2bN3du27zBFZ4cZyc7UVBEQ3mKQXj1cepDoKFP8VGrpnXNM8aczJr859jQNS6RHc4ihiA3ICbXrVy6EFIgqTjR2zauWX7T2pVEftmIXDJzGzqOvPkLhUZ0HdxPdNwjRQiLghwwkdzvf9Hte+GBnv3gzUa1Vi6eP3vjmhVLXpId+87Sl5FiifuDf9eO777FvNBWwaIlyjC+lYvnhRJv1uJNTLlP5+8HDIGY4ZmxRvjMnDR+tOlH4OYNax37Fd5zXKxM+co8f7VfbdaybOUadXie//xtKAT+gxsS4nBLHmrTpiffW3yf5ytUrATaRZPG/vqLacMQII7fc45Y8jl4ewD/BmlRBBQBRcCnEdBdZT49fdp5RUARiM0I7JcctcP6fd+VvLVVajdobMa6N3hH4E89v/48No9dx6YIKAKKgCcIkDIKosFScA6TwgjD8bhYDMc6352k5qGQdq+RWEuxRWLoYJD66KFjmTZpO44WIxKNExjHC1gixMuGJ5zx5MA/KAbwOOo5RxoohKd5xREGYUFaKdKo4NQP1X4QR1f0h1WEPamsASNqi8ONtFB8RisAcoZUUYwx1BknhfV1TOySGGnKGDPH0PKgnlXoGALokfFnEwFnnHnBkpbIVbc2SlooIgbYQW6cstQlBz1OzIN790AgPVL8CxUribYFwt2O5xBXxlmLQ3/WlD/HOp6H7MCJXrJc5WqSLeqZ1g2rlbl29SraHlFW2IWMbgBO+19/6ovmzMNSsnyV6gg0W8fKzvHW733aee3yxfMXz5n+0BGd3R5psX93MKnKHhZS/+zfvWsnjmhnncbZTcoU7NC+PbsG9er6MGe/DDX0C8V6fz7jNIQ4mDBm+M+ugMiVt0AhnI6QDI51uLZJy7YdSL20bsWSBdbzc/6eOM6xPvn1OSZrY/O3Pw0fe+JIyCEha4jcCV1DIj0RqkXh2E+OffzVdz/g9LaOC8ctY3BMN3rl0sULpOiJssl1aChHnvwFt2/dtD4i7YeF56vNWr3NM/BDt04fWTUIWPMjfurd43E8CxdjzZNii5Rfs6dM+P3v8aOGm3omIsAZntSBLNuwajnPdpSXt9p/3Im12P/bzh3Pnj4ZmrLJlH8lRxfvcbjzXDrevGCxUmUhEBIlSpS4cq36jd5v+WrNg/t2P/adYK6DuAkK2J+2tVIAACAASURBVLLJSmKYc0bXheeM6BXWa+8uHTtIRrJD1AkVbneitcK5zj37DyEFVffP3mtjJfRKVqhSnc8QGY599yamfI/Vatj0DYgSyJxHMf2P3OL7c8f/sXce4FFUbRSe0DsqIgoiqCi9d5DemyggIFVAepEmVZqA9CZduvTem3SQ3nuH0HvvBLL/9y5780+G2WQDCSZw53ludnfmzi1nZje737nfObtevjcDuu/IboJ0hAxs3KbTH+OHD+wNkWh3UwT1cytpitTp+GycPmEUPl3ODempDFly5IIsC8i/MFW6TFmc/iwWP45gv1l1gxoBjYBG4A0goDMs3gDIuguNgEZAI/CqCIz6s3e3WuWK5eEL8ZK5Myb36vhrk2qlC2YPiZVdrzpGfZ5GQCOgEQgNCCifC5vHJ7KP1ecEr9CjrytFyVmgMf+dFFZ2e0tB1x0zUT9DWgsREhqm+qbHQKCeQDXEBbgklQIRAUmBJA+SIhAYEEH4L7Dim2AbvzPIuIjjOh7FdX5Y+P2hvCx4ZLxgABExQwpBaOZJJg8BwTFSlHfFTXnOPQY2+FhA8kAWQGCAnyKB5On/NxWUDsgcmgwLAuxkPpjPJbjofer4UVZl+2tUXmDcevyIfx8sVadOszYdCTxu3bB2JcFb67nIKN2XICnBShZJvMrKeGub1tescCeDoWvrJnXUSmzqoDfPvPBcMJ9TtkrNusivDOvbzc8MmuB7tTqNWxAINWcDgBXSNof27XK70lg4my8JUFO6t2tWn0C26k/5ftyRQL55DJBLkBGH9rpvF/152pKkl5e8Buo0be0c+4Cu7VsGhg/HCSwTfCcoTyCzQ7O61c0B6wQuDwI0+c3tMQYkRckcIMtGHSOrhu+Qa5cvnm+uv/XfNSsVeePJuIJSBxNr2t4j2TpBOU/VdYcn161W4xbtznmfOjHj79F+2TkB9ZE6fZZs+L0gr3bv7u3bfK8210+Q6IWngxVP9uFJQrbL3p0vslqCc+O+rlqnUXPu4enj/x+oVn2QZc3zHa7MH2vfvF8hBDDehviCbHA3Pt4bBLbtgvSck1R8Xbwl8wLSBKkk8DJnYZH1A8FlJTu4RyFL/hrUq+v5M6chs/22nOIxckw8+aykZ0hiSue833j/DPqjUxsrHmIJ4cQU/wrzeySw+47jkCw8kllx49rVKyP6/dHJHd5B+dyijQxZc+TiWm5et9KPYKndtFUHcOd3YUD3nZybOyTuz+C813VbGgGNgEbAUwTCwg8GT+ei62kENAIagbcSAX6E92jfomH7Jj9XmTZu5GB3KwXDyuTR0Q0rY9Xj1AgEBwJIurkzRA2O9nUbniEgpMUzKayoRBqFIDuyRRgmsxGwJeA+RQorQDEGTSLFvDLes47erloqcE8gl1Xq16WQqULGAXI8SN5ABhGcuiblcykE7FNLwfgcWS7kepBSIvuATA2C92FhY+6QABSeqyyTqPIcgoY5c994u3BgH3OH1CEDg4wTZLHIqFBZFb522SUEpQOTy7l6+eIFZHqQITGDR3BRMgvUfex3CCKAVcBkGFjBTixGwSXLVKzK/g2rliN15W9DCgqpKUxeT504etguA+N1LyCrwTGP3rVt0wYlw6PazJGvYFGOWwPc+DdQV8m6INnSd+TEWWi69/ytZSPzmL6UleEcD8jkWfkUsPLaOgawo70LrlXlqm1luB1QuwTYD+/fu8v6fY2gM/r+/0owWa1WDwzH1OkyZWUMBLNnTBwz3CobJgbhTn8SMmnMbYEV/SspKI7Vbda2E1k6fTq1birKSbwf/ba5YurLi3JCCgU2pqAeT5E2Qyau5z6X3FJQz3eHJ54leGLMlAwJVskH1i7kliyKTyMqRU8xO+/TuU1T6wIg8CRQb7eKnRXu9GEl0gLr15PjpeR6kT0FMWAm79S5KutBSZVZ2/w6Req0EBGs5h/S+/f2AfVJlk80SZva45ITM9flOtEWZAbZOBAQ/bu2a2HO0kr8xVdJIYmsffxYs14TAv8z/x493HwMuTIyNUR26SXCKiQxxdsGyTmRxVp1Wj7HrONVHjjuMHV339EOGPH4cfxPEw7u1aWdHWGs+gvK5xbnpBMfitMnjx1R5A6ybnjrTJ/w19DFs6dNdHdt+czn/RAS96cn97CuoxHQCGgEghsBTVgEN6K6PY2ARkAjoBFwiwA/9DG9y1Oo+LcaJo1AWEOAoNja/Wdu5JCVgkEZO+aonfsN89NKDsq5um7wIyCkha8UAuhrpbDKOa+UXlKUhjX63WWkIF/SV0psybKwNUoO/tGFuhZVRgDzR4bkihSICTIoDkkhaM9+yB7qQEYQGOI59dBPR0ZEtRMW5KCUn4UiayAslKQSpAWB3iNSdklh5fonUsg4UZJQSGFRn99ZZJXwqDIsbH0s0kqAe//uHVsDu/rbNq1bnS1X/kKqHsQCuvWsXLaeizcD++z8KwhcK8Nou9W4CRN/kUTppY8d0q+HnWxMYGMN7Pg3+QsXp58povlurZszX6Fi7DMHVAl6Ypi8eM70SRwjEDl9+aY9mXPkyteidqUyyGia20Gjn9cBEQsQN9SZL75g1jHQF/us2CITg1yQXcBWtUFmi/KWMLeLNA24z548dmRg+HCcTA68H5DvCi8vhvXp2sF6HtcfvXzrivbseQoUXr9y2SKICXDGtJnV8sP6dOswf8akcdZ29olcE+RRGZFYCm6CndXoBOGPCInjybytddzh+W15IWUks2jhrCkTPGkXLJ3+AJjIi7fDqiXzZ5vP4/305dfJUuLXYtceGSt4QdgFvz3pP6A6kC+8zxbPmea8v60bZsqsuneXpSJ8ACSxsVCyKwLLhiIQT19cc2s/ZDxAZuC/gjH5lg1rVuCloOqx6AifCohM87nsL1a63I8L5N6yymnlzFf4pfezOjckMc0nmNLPotlTbYP8YMpxt4SFm/cx50CG8EgmivU+MuMS1M8tzmVcyORxHTr1GTK6ZaeeA5A3s5Ky1msHluzbLe/j170f9fkaAY2ARiA0IKAJi9BwFfQYNAIaAY3AO4IAKetM1cdGuuIdgUBPMwwjQFCR1YsSMwh0JaeaJgEQVsvdv/tCK1lvoQcBIS0cUtCpJ6MCORFICmSjMFqGtGCFNXIhBDOzC2nxLhMXStYIYoKsE7IJyCBI58KKVd7IRoEdBAaSSQTw8Xtg/w0pKtMg9NwEgY/EKuHE3CBrMOKGYFDSV8zP21UgLyA1mLuS4oGweG6XXYFZLkFCjwgLkYUikI40CENXwUWrHwHH0FfnEbko8zRZNV24VJkKBLiRFrIjO1iBzTk3rl+9smKxf9PiwCHzrEbR0j/8yCr2Nf/4lyZCpip77gKFL5w7c9qsw45GPy0/kiXcY2YvWz9y2sJVmNpWLpE3M0FVa69CWGQgSH7iiL3hOPXBgkcxEV718vnpM9K+VRoomQS9Mft2R+Kwyhlye8+Ol018CaCyon+jxbvCHWJkA0AcQXIMF8kZa1YE51HnhJA15hXwrPpmHOjddx0wcsK8tTuPYBTe/OdK3wckKYOsDdJEZL54dhU9q5Upe668oky2O6BV6O5acoen2KrEyvJNngLbN65fHZCmv7ldslWcr+WN2LdL22bWPpGtAm9rtoqqRyYUJFpwE3hkAqXPkv0b8ZTYevnCeaTm/G1IpCli0s5Hhu8lZENx0nSTSbM7TNOkz5wNfws7nw6VsQPpUbJsxarDTfJrtKc+V6wYQbjgwzPHZe5u7jtX/iIleL1355aXpLRCClP6y5GnQBEyb9aIX4wdFtly5yvE+8aOXAzofezEQTLQXuA9ckhA90NQP7f4fIcQihIlWrSZK7fuZ4FMg8rfFcFAPrB3W+oMWbJxTSE7Aqurj2sENAIagbCAgCYswsJV0mPUCGgENAJvCQL84GIqVkmDt2R6ehpvOQJJU6YmOCsrlt0bWVoh4Mc9q+Q8CUa+5fCF2ulBXMjgkDtC3gfj38JSzKvdITLIvqAUE+LiAyl+36HfRo8L/FRNxWq+rTIHyB5A4o/XZKxQD3ICfxC8HSCDcCyH3GD/Sx4LofamcA3MhYGZtOA5pAVm2zwikQVJwxyRgcK3AnKSrBLmr8yebb0r6AZjbB4JVgaGx/ZN69cQYCOgT10043m0k4RiVT7Bcas/Rb1mbTqRdXD54vlz+DuYjXFV/0lcq4eXSDaDJ1I7gY3behzZGTTt169atsjaf06Rg2KFvzWImC7Ti9XDXfoPH4e0Uqfm9WtULJYrgztj4a/l8/rEkcMHzL4U1nEQoMaUmlXz1mOZsn+T96DgZB4fxrdfiFYWZuDu5pw204vrKfI3KmPLWRUigCzTHZv/XecppqnSvTDcJptj9pRxf1n7hOyCHDlqkYNK68KqVuOW7fIWKVF6zJC+f5TMmebLNcsX4bXiduP+QhqrQo06jZzGysGw0Q7Xziq55WnT7vBE5/+FB8ualZ62lcq1aAZZHWtGDm0omR+J976UYcH1Q9Zorw0R5Wn/7urRLnPZaWNIzTkFipcu65RI27HV3z1lfb8eFi8Gu3lZ+wVT6/2p6uDRwnNW68tU11m/u/yfsPCPEVlR+G9YyVMyL3LkLVAESTsrGROSmDIHPsd4r9r5U4A55dTxI4fsiEB39x3tcq0+F7ITQnTpvJnISLrdgvq5ld4lO5anULFSfDaVyZc5hR0ha9chmUNkzQQ3ofa697c+XyOgEdAIvCoCEV71RH2eRkAjoBHQCGgEgooAPwZZNWk1sQxqO+9KfYI2GbN9k0c8Hj91OAzH5Yvnzm5et/qfV1ml+K5gFpLzJDgo6hq30Jr3tJ+ULmPGA3u2BxqM9LRNXS9EESCTgNWJyH6xoru1FGQj+M7MinX0/vFtqCNExSEhOwhcv/UbgftLd54YH8eKhJeF73NfR2SJwF8J7+VF5kA4OQxxATkBcRFRPq+iyj6C9UgogRH1CNrbbhbSR/k9UFc9V5Jc6rVqy/kao/UQ3sxjZ04QFGzO+UtRhAz1wEAZbFPHea5ddgX7CYwRFD+4dyf3VYAbnz+sbM6eO39hvAkwYWafnQRMXAnqX7pwzt9qbRYNFC5VtkKjqmWK9Rw2ftrsyS8HwRmAImeXL5g9PbAxvcpxiAICmTsleG89n/ERcNu/axvm5n4b2uyspO/W5pe6BN7NGQXWNgjuCjZpJTtkVkDjYxW13ec531Xob86UCaPM53+ZNFlKJIWOHtyHb4vtliZj1uz4U5izQ6iYXKSkyLjbaZLXCQy7VOlfGPuSFWFHcqgAu2R8+CNQ+M7Aef3F2Bv5KbuArbu+J44a0r/38AkzchUoUiIwgiOw8XOcICoZBK/uX2GPp/IS2bHl/3JFgY1HCIssvNcwhbar+5Vkq7D/yIE9LxFSKcWkmut3YM/ObYH1E9TjBL85x53cU5lK1Wtz3J2BfFDer3iz8P5zhwFBft5nZFe0rv9TBetceA/w/iTLyHyMDFS+n1rrF/22XEUwtyOsQhJT3r8QIrvdGL2XrVyjzgtMd++wu17u3sfU/eLrFwTTv6v/WRLY75mgfG7RtvL0OH386GF+A1g9VtzdW2S3QDYh4RfU+0/X1whoBDQCoRUBTViE1iujx6UR0AhoBN4yBJA0QGN33YqlC9+yqQX7dPgh1KRt5x4VfqrTiBWd5g4mjRo6oN/vbZsHe6e6wUARwNwW6Y1AK5oqoN2NrIioL7ykMR+UdnTdkEVABbxNgXNWzy+TwopWdO6RjFFR8czynGDNQKmPuehxKW6D8SE78uBpPZAsEWc2yeW7TyJeu/80SqTwXs+EoYgghESsWFEiPI4ZJYJPhHBeUZ/5Op4/feYbTYCILPGsB1Ln0tPnvg8f+/hCKoQXksP39qNnXtKX8nGgXZ47j7uesy+66zX7zabXmHdzDHIA4oQV4Bz3cY3f1h+CsQcjoaF8LdT1JpuCcdI394xdJkWAvh0EqFgV7WlQefvmDWswceV/KgFrd59JceJ+FO/G1SvIUvltzX7r1ofMBWSOxN/3PXc+DMlSpk0PCRJS2ZAqg+O46ASZx4eUUfJUaTPYGTSL6k0ciIBVSxfMCeyuh4hAMiiwz2tp8kNkk6ztlSpXqTr7Vlv6+lpMENgvMlNu/w8QuN1rya7gHILEPLJoI7Dxq+NIGCHxsnz+7Gl254jdgjPALivr/QXYwYr9M/4ePYz/P572R721yxfPp8/cBYuWDA7CIrusrqfdfbu2vuSX4Mm43OOZ5AWeZz3DE5kd7otNIsdl9ftQ4/hKnK15H1plwDiO9JYd1p7MIbA6yuD9/BlvMrP8bVlz5SuoMqnceWvwfuWk1W6kj8wNQiDx2u4eZT/eDIxHeZpYx0OGBSbwZjkpyEckqazZFRA8+YuW/P75c9/ndoTVm8D0gg2mEAHfVaxWi7m5k/9yd99xjrztPMY7KJ9btA2BzaIkSMo/Bo+ZjGSWJ9lJ4oOenN8Oh/bt2RnY/aaPawQ0AhqBsIKAJizCypXS49QIaAQ0AmEcAWQU0AYOyAAzjE8xWIbPD7y+f02aTTo4Uhfzp08aJ6tkz4iqUEzkH1YsmjszWDrSjQQJAX7Aoxu/buWSIBFuBAcOi9GopxIgQRqUrvwmECA4TjAQA962Un4xddpUnlMKS8Cc1eD4FfgRF8EYJH8T86QPAu/8NqBABigjbcgBsiSSCOnwxWNfR3ipeV8Iifd9Hc9O3H387Krsh8yJKaRFDBGTihwhvNdRX4fD59lzx2cCSER5fl2yLiAlaBcZJba4rnbJRiDASh/IKOGNkdz1Gi8IMhYI8uIpkkIKJAE+EZAEBPhOSInkahv8nSSGFNo1Zzq4ug36Axkmps2PlLCR3lAVA8yqUG2x8jxF2vSZyJbwdFQ7RLYHM1zIUFZWr162yFafHSm6a1cu4bHh3Fgxny1XvkLVvyuY43MJbrHPLjODYB5GsUEZk6djV/Xii17Vi/4vIh/mtzVu07kHsjIJPkv0uTU4G0sif3hqeNIXK6CpF5B8H6QIq5IxrDa3yarsUj9Uqo68jlULnnbJ7Dh94him6y9tXE/xAEhrp+PP/29OuOZhhh6ECx4b/yycPd1dViUZM6xeP3nsCBJsfhtY8eJV/MKQuTm0d9cORSp5gndAdZAvI4vl0vlz+L4EaQsMT3Ahw8iTRnm/UC8gEgb/BkguO0kd5IOQNbLzffCk/4DqRIseMybHr1/zTzCSzdOiQ/d+HHv65PFjd/ez8CzpIR8DMoJX/SNBx/sI8s86JvBO8FniL9hPpo3dmCEs9u7c6s+LQnjGF+9n0Zkzn1O6QtWaPnJDRY0WLbqd5F1IYsp3ZjtM2dewVYdufD7y/NDelzMsArrvOCdZqhcEEeRXYNc+KJ9bKvtll5hm/7No7oyGrTp2q9+ifRc8LALrRwgL52ceEleB1dXHNQIaAY1AWEFAExZh5UrpcWoENAIagTCOAEaVzh8HbtKvw/j0gm34NRu2aAtZMWfK+FHd2zatF5DsRbB1qhsKFAFRXslIJXcrHO0a4AcxP+4njx0+KNAOdIVQgYAbkoHA+BUhJZCHGiEFLflcpgEjgwGR2FsKUjFOU3aVtRCaiQsZIwF2gv2QCWQvxJNy0/VIUPtzKcqXIZM8f08i8SeElrnw3OH45pHP8yfyvJjszygkxl4hJeRz3pHBx9eYIcTFQQn8FZP66vzEUo8V/xAMbEmkfCzFW0ps2payRArSWxWlQBQh14FPA6tGkerCu+FfKQlc50NoUIfzITogNg5LIbBN0JbHBzJPpJueuvxKXN2//oONzFOQMm3SiEkqq2LtTF/djW7X1k0bCFIX/758Zbwc7Ay3OZdgvMQ4navrCcK36dZvCJ4UrNatKNl77L9qIQzYp1Zz42fw+gjZtxAtxosA7TOJZqoaaSQzAUkTbyEDWCWsvCfIJGG+D0UbJYpEEj0ZUzyJoFLvjDAL7uoTlEZuJYo0aq5TrW6TlpgY9/ythRMj8xZPmBaJyZ4leGzXboo0GTIRZGZ1uvU4rjDsk5gwmUL+ttTirYBvgrldkTzKBKmyZf3LhuLqZCSMCDxbsyjAijpyC0S1EjLWvvkfBaFglrbxkoUT5mvjCeZ2dTCLFvPzjIHp/LtrP2A8DS/eO+BtXhDAPqS0rB4NirDYsn71Swbt9C/8UGyIus3rV70ka8RxsjNuCNukxsq1CcgLIiiYqevOvWH2U6lcq0FTiCOuryTmnLTzY4kYMVIkCMgFMyaP96RPVuzb3Z+cC4HAohnuBztiB9KNckreoua+FOFivmfI4KrdpNVvS+fNmJI1V96C+MFwjno/hzSmT1zvUcgH81h5r5WrUqueQPqQY6dOHOX/hb8toPuOihDFZOHYEb7WtoLyuaWyX3ZueeFzM+iPjq2RZytXpWbdWZPGjjS3zec70m+KpIr/aaLEHDdL0UGsnDl1/FhgnwGe3De6jkZAI6AR+C8Q0Kbb/wXquk+NgEZAI/AOIpBC9JsJEAhhodOV3Vx/5DBqN23VYdvGdavR6dZkReh5oyRPk95JWFh1mwMaYcq0GTPz49wTM93QM1M9EncISLD7iRRWVpeUUkIK2QBq+0GeIBvFSkhWUvstyQ+NptyYhkuBqCBrAckrgv2fSCkopYAUgrWtpNR3PW8sjx9JIXsBYgFt8zJCUFSRCH0JKd/K8wayLzvtyPM6klVRVvZ/L69rSuF8ntMeK4YpPGcfx6iDuTk41nONhbYYR2kpYF7VVYe+GQNjYUycTz3aY8w8Zw7MhTkxN+b4IXM2G6bLvv90Uwar7gxw7QbHCu9Dsvr/O1m9zHF3JruPRNuG4wQgO/UZOuZ90cQZ1KNTG/bFjPUe+NlmWCgdfzIMQgqcO7dvQooZ8RO+CLLFlchbzyHjpg7o9tuvEBes4EZmZvTMJWsJ2FEH6SZklcwyicytRJkKVTr1HTrGPFbhZ5zybZjWBjQH2vwyafKUBJ+pRzCzRsPmbVhYIf4dL8kwxYgRK1ZAbSLvRXDQmplB2yqwKGbReOP4bdXr/fLr3wtWb2GVvHl/ijTpIQiNHW48LwjUk/FhJ2+kZK6sWRLpM2f/puuAkRPIFlR9jZm9bH2/UZPnKAwy58idL2PWnLm3b359wqrCT7Ubco3+Xb0cIjLIW2B40jZzUg1DVvQeMWHGyKkLVnLMP54ZMmE0b5dZQD2yK3h0JxcF3lGjvViVz/Zbz0EjR89YspZMmCBPzHKCMo7PXbBYKXWIeTVq3bH75nWrljMvq2G1qgdZwXFP3q+QG6nTZ85qNdJWbfFe4Dnkh11WqDLcFj7jgnkKd2/fcr2fP0vMfsbTY8jYKcvmz5z6cYKEnx09uH8PmTutuvQetHr3Sb8sqZDElPcABE8eE6YQaD2GjpvKeCF6IS3MBJGaU0D3HXWcZt77PfstE5TPLeXLslPMzumHjOolc2dMbtO175Ai4gVixrxGg2atpy3b6OcjApYcjxothvMe5XNxypL1O/HBe937U5+vEdAIaAT+KwR0hsV/hbzuVyOgEdAIvGMIsMqOL+6eGsi9Y/A4p/tTg6at+ZHdtVXj2naSBO8iJqFlzvyQ5Ad8QNrl1rGykpF9+3drw+3Qch2DYxxCWtyVoDdSEATB/5RSXArZCQSuJkohQI6h5yQpQdKPD47xuWvDlU1BYBapJzIbWFmeWEoqKfgvIJlCNsMNKRAZZCgQ9GMOSDlxP/OaLAy1Kh1zciSa2JB1UsEojptlLAL6zWE+Zj6H1ff0xUaANbWrX/okCENfZL+QZcEYwR2yiHkga8J4yOzDJJdVtmRoeFNXsGClNIQHht1ByopwjSdYHjJkyZ4L2aag+BrQ8dp/Fs9nxTj/J07K0ny7wRAgRwJq5LSFqzJlz5W3U/P6NZREFCvonRkGrpX45vPxxSCIZ+ftECyTlkbEbHst/f/apdegVUvmz65au3FzVnTLyu2DZI0IJ3P77/mrNvP/sE/nNsiuGQQ/i5Yu92PH3oNHLZk7fXKiL79K+oOslCZgO2/6xLHmsUk8knvYqFb3l5a7tm5cTzZKnkLFvy2WLWUicxYDq79bdOzRv2OfIaPRupf/wa2e+Tzz+e2XOtXs/gfTbpZv8hTIV6Tkd7T/Q7Wf61OvYZXvuSclkJk8FWTMT/Wbtsor/VUrXQDSzbltWL1sMWbGHHtw795dSI3CpcqUR0ufFdVWnXoIC8gpdwH2ROLUDHmjiCnz/FcKpq279hksgc7BI/r/0RlZmpJlf6zK/YBm/z2TjNK6FUsW4InCfSL/4nyy5sxTAFmuSX/ZSwJ5eg+Q1VNFrqu6Dtly5y+E38QVIQ1uSqoCxA6ZM5FIcREmgIxE5Mjwmpg+ftRQZIsCwnPBrCkTylWtVa9L/+Hjhvb+/bcH9+/fq1avSUuCzaPEVNu64IPvoPt2vZz5ouajyB07PKnD+4HgL3JCZCLkL1rq+4HdO7QKju+0ZNGwMh6PGVGHihU5cuQo3LvcW/Qxbu6KjcIB8Bn80kZWEjs9ydJCag2wyX6YsmTDzhH9u3dav3LZItXo5yLdyjWZPXkcWYQvbYqw4D42H/Q+efwocllV6zRuQZZFIbmvuarD+/3Rac7aHYd3S1bYoLHTF2QQIux3+X6rzg1JTHnvrPtnyYJCJb//od2tG8OQcatSu1EzMmW6tm5SB3IoXPhw4SHqrO/1gO47yD7u0z3iBeTJeyEon1tJxYvkhUH5NiQmnVvnFg1qcr16Dh07FT8QiNSo8l4B67OnT+Cf5dzIpOCxZace/eXtdeXHGnUbYwq+cc2KpZ6MU9fRCGgENAIaAY2ARkAjoBHQCLyTCLDKfPOxKw+6DRpFMC/ENlYYEUggUyHEOgmhhtH4/ffwxbudJHASQl3oZl8DgaVbD52dunSDP2PTwJobOHba/JW7T/gzvQ3sHH08bCHgWrGfWR6XSnFYyhF5nfi/XtHvyqaILI/xpHwtJaOUilK+VhZsSAAAIABJREFUl1JayiQp66TskLJCygIpe6Xcl4Kh9Xkp+6U8c83vnjxe3SXzleIrz8+Z5v3Atd+Kxau8RspJnUcf9MXrq1IYA88ZE2NjjIyVMTN25sBcmBNzY47MlTkzdzAACzABm/8k63z9wXO3uv85GmIrSBsGtxuPXLo3c+UWt+bPOfMVKrbr7B3fnWduP6/ZqAX+K37b9z9W/xn8lDSU+djkxeu2s3o8SAN6hcrIxTA+xsF3A74n5C1cgmvk2Ol961nPYeOmmVevE1jkM9V0TzgmLVq7rUDx0mWt3RP8nrFi8z5Vd/vpG87V3dZ6BG+Zr6q3bNvhc8j8uJuOeG5nWLv/zA1Vn+vHSmZVv0nbLj05tu7A2ZuQK9Z2GOvWE1chzJz3NfPvNvCvv5Wevrk+45+3btdRd2NJkjRFKtpo32MgMnUvbQQ0zVjxP4xsDnOGCicRDB0zaynvEceGQ+dvk4EBb/AKl9TfKRBPfO/bdur6E/M4AnvO/0xlUB4YngT4ze3RHyvPrWNnPtQL6L7mvUAd60p21ZbEub9gbNTZcvzKw1qNW7Z7XYzM50OAmLFasvmgd/bc+ZHAM/4cP3MRr+36A4O5a3ceURkyAY0J2autJ689Zg5DJ81dxrU31/+1c6+Bv7T7vZe7NiBrOFddH3O9HHkLFuU7LMenL9+4B+KJ9tX7mX2JvkiCF5TfFtKYMs5/dhy9oO6RTUcv38f/hwEg/cZ+CAzrfAO67/AC2nH6po85SykgzIPyucV15PPI2h6ZMVwX82cH9wMEk6pLVst4IbbU5woEh1UOKzjvV92WRkAjoBF4Ewj4c5B7Ex3qPjQCGgGNgEbg3UOAH9YEVnp1/LXJtHEjB4cUAgQ9CB6sXDxv1q/1qiEtEmwbASJfWfp08/q1q8HWqKkhVoASuKpUPHemwFL7MebrO3LiLFaQNa9duQwrslRTYN1CVljNm/r3mOVi1hkSY33X2kSzefWeU1dZdYhUl6fzJ7hxYPfObU1rVvjW03N0vbCJgAQJWP36lRT0z/FXUBsBRySNTkpxeluoLaS8LUzBdySfyCxgPMjLJHO9JqOAfWQl4C/B6nA+1whSso+VmmRcJJGKBJiov0t+NGSRJ2RDsKozvDxPJEciyuNtORZbRLDwkfC3WX9ovOIPDzI4KATXyLrAvJfPPPAGUzIoyKSgecaORwbzZuxkeiBXgnQUWTFkYbAPSRPqM09kvtBXZx+vMf825PqQvRGiG/JHZ2R1stk/wNMOCZ7fuysr8EXb3t05CRN/kUR8iR9btdb5H9Kl3/Bx44b172mVo+J/EStzPTUz9nS8dvWQgmIsyLOwarnPiL9nZhJJoh7tmzewarar81kpL8ouH7OqOyCTYQJ4XyVPkZrHU8ePHna3Ep6FDkpWaJ/4e7jzp1D9Q6IgnYM/CCbIZl8BAoTpMmXLiaSVO9145sxKc0OWde/bvW2LOzNqVrNzDczG6VYM8RthlbW7vj5N9PmXYsabHAmfY4Kx+buCtS3+z9GfnRTQq15jtXodMiqqYBMlSrRoYBRFVmioR+pgnv1QMiSQ27olX7JUdoQneH4l8jxfi6fAfXkvkE1Ddo7deMl4JBtJlNLu2x3nPhC/9AwH9+7a7i7DlXl8ECfuR0gKuTNCf1WsOI/vmbyvJbnkstxbB1QfZD0lloyifxbOccqjmTeyp8h4sJMhsxsLRu0OAdjT+uY28E3AYJv3nl3bTqN4GSdeX8/lRiLwD0k2b9rfY3q0b9HQDrOQxpTFQLy/kX9CPk/dH5ApZDdNHj10gDUbJ6D7DoKD9/+GVcsXB+Vae/K5xbXEeB0fH3f4pkyXMbPcqhGRjbJ613AORBH7yTgKyvh0XY2ARkAjEBoReMXfDaFxKnpMGgGNgEZAIxBaEShdvkqNzv2GjUUewSp7EJxjHjZ53nJWpI36s3e3YX26dQiutvlBPX/97mOkdg/r271jcLVrbodADWTD9/ky+a2YctcPK8NYVcfxqqXyZT2wZycBO7H09PJiNRk/eoMaXA+JOb0tbebIU6AIqxGRMpg7dYJHGTCsvlu65dAZ7kPux7cFCz0PewSEJHC+BaVgUv27lMqWmqy2RpqBin4SRJ6SFq72rZ3Tn/ouzyOBeLUvijxHQulLKXymIPVEcB9SgUA8gXlIC2SR4kvB7wDta857KgPENHi/r8MoKer+scWTYr6cROA/gzy/Ed7LeBTOy4j53GHEfeprPBX24H4ELznP4WzjczkOscG+DHKeU8pEnjs3aXMNAEhKQz4Gwm5pC1B85M9W6S+GvISQ8KYNKZyPSTNjQ4oEDKNI/Q+l7JJ2IFqQ6IHUQN6EeSPFA2GDOTJtINl1UQpyWBATEBpkVXAOY8UsHfNVgv9kLXAew6RA4qhrpvbJrv9vnl5HfyfpF34IIG/Va/iE6QQDTwu5UCZ/5hQaHo2ARiBsIhAnbryP/xg8enKWnHnyM4MC6b+MF1KLfcImQnrUGgGNgEZAI+AJAtrDwhOUdB2NgEZAI6AReC0EUqZ7of+P8d5rNRTIyS1qVyoT75MEn7pb/fWqfbMyj5WqITV+Vpih7zxvmn8dbnfjVStFWRl75MC+/5vuyRJBVsCxio0Vba86X32efwSSpkrrNEMNink2htvOc/bscJJJensnECCYfUrKT1IgFFtKUXIxU+U5gXYMpRdIcRoiKyIisIC3Ou7K5KCf8FIgKPBp4DWrKfGiSCwFEoJgPEF8+ACC/4mkwA9wDvUPuh6pLxyCs94N+RNdKj0QIiLcE18Dw+KVsi+Oj8PYcPWpETlyOOM5BIXs2xI9vBFRiIaU8jqK7Ieo2RMlnBFBzrv10NfwEtIi1ocRjUcPnxv3IC2kzj0hNCJf9zG2P3MYXh9HMu4KOfFUOo8i5z2WtmJIW7sihRMyRDIhZAzHZd9zITogW7ZLGz7PfI1D0u4TGW8mGUMUaee01HHIc/xDIDMuy7lpZTbXmIsUcIbo4DcPc4W0IEvjUxc2yqeDueKTATbzXFhBbnhLwSMCwsSJkRQIDNoI8QwM6eOt336sWa8JBPw/C+fOEF/epxiKv/WT1hPUCLylCGDa3mPImCmSKHAJXxq8WDRZ8ZZebD0tjYBGQCMQwghowiKEAdbNawQ0AhoBjYBhELw9dvjgvsCkFl4XK2QRgpusYEzZcuUvxOOubZs2vO4Y7c5PKT/o0BbesXn9Gk/aJ9ND/BcjYTRqlqPgeflC2dOQzh6ShqmejPFtqpNMLhAyEiflJvZ0Xph0IyuBvISn5+h6YRcBCAVTFgSZDPukKC11RVoQVJ8ihSydJlL8DLndZFAoQFTWBMF1zKTJdCAQT0CdIDsZEhAWZFNgAE6AnuwCSIrzrnqYV1OHwDzZFSklMh9VCmNAQiWCkAm0ee+Rr3H/sa9x784z41pEL+OyROVvnX7kuH7mkRExWXTjguz/5NYzI5wQCk/TxfQ6e/6xI4kQEw8ieHn5CtNxJ2p4L++7zxyRpQ3fRFG8Tku6xo0zjxxRbvgYZ4RpeC79eAkJ8TxDLGNb/MhePlLvU2Ffwgn5cH/ffceJuJGMh/L643vPjfvJo3uleS+CM6PjttS7dtPHuCmERHghS8iEuCXjYOyRpL0ZQnrEFrLDESO8cSucw7hIBoic5yVzlAfjihQkpTDlJgtEZVnwGjKCLBSIHogMPJCQhSLLYonrOHUgOyB/IH3Ajfpc6+fohv+X5t0yhjC3Ycrcue+wsWj3D+j+268zJowetvHoxXsz/h41LMxNRg9YI/COI0CGL145DVq0/32ZGEOTkTps8tzlh/btRm5PbxoBjYBGQCOgEQgyApqwCDJk+gSNgEZAIxB6EOAHAqvz3WkOo8mLfrOdzqndLCJLpPurZClSE/gPSnDWuapfBJ3t2sTg8esUqdLiqfC6yDEfNJjt9IXRbY0lxorutF9fp2/xtUt18fxZb/SVX6cdd+ei2c2xw/v3emTqjDbttPF/DbFrz6pVbq6DvrA7He+QmNebajOcbF+KnBYkzokjh/YHt7Z0MsmwOLRv1w6rznFA84OEOnv65PE3oQP/pnDW/QQJAVbqE+Amo2K1lLGms3+W56zOby8F8iGglfpkUiBnBAlBNgWZDATVeZ1UCt4M7CN7g+/1eaUo7Wr8GtggPOgDnwokochQEN5ASAJf45gQBQcl0yGSZEbcu/fM2CXZFEhFPV10zXFMTnomZMBVqfv4/QhG5MMPjOhrbzmiyTmfIAElWRdHJSvCkOyJy/efO3yvPTWShvNyQCo8FvIgQrxIDu+EUYxr++8bz6Xtw2efOO5KP8hIRVp43bj2xNcRI1YE407CyF6Rrzx10NQDiA5p2/fjSF6xhAy5/lEk45qQKA+F8HD6B8n4fIU0OSeESRRSQ8joEALj/nsRjVifRDKepYnhFV9ehxcC43zMCEYGqf++tPdESko5PfUL9SlnhgoEEm2CLziyH2IHsocNkgIskZei7mlX/UPyCBFERgcZF2SzYGT7QEgLPz8hVxv6wQYBzHAHjZ2+AP+KepVKF9q+af0aNN75vqIDnPqW0QiELQQwjceDLVf+IiX6d2vfcvLoYQP5fZJUvDfGDxvYO2zNRo9WI6AR0AhoBEILApqwCC1XQo9DI6AR0AgEAQHxpvzgl3a/9yrybbmKESJGiDhqYO+uowf36W5tokOvP//6QhiIat/mz8YxTBzrNmvTKdEXSb4mKNC3S9vmKoCN90OPoeOm0jZ1MadrWadKWYKudkODPKhRv1nrijXqNEKv9siBvbvrV/6uMOZ/5vpJxQyRIMT+3Tu2qv1xxDHzh2q16iPftHrZwrmBmdfh7dC84x/9suTInV9i9XfbNqzx4+b1qzG39ds69h4yOq0YmBbM+NUnVgKHfhq16tgdLwE1H8ZfrU7jFgRJyFTYtHYlhqzOjR9aLTv1HIB5IMFvDPuEJ3mO0TXHn0kHR0WKadywAb2CcNn8qqbLnC1niTIVqwrUceiLDBRImFZdeg0ytwdB0rtT6198RCeD/aTaFy5VpkL3tk0Jgtpu/HCEcLKSOgSIMD5v/nOl7zeuWbEUoqvKzw2bFSxeuizzmTB8UJ91K5YgVfPKW5XaDZs9FiPSWRPHjHDXCKtq7cwAK1Sv05CxmzHFHLJmw+ZtMKAc1rdrBztjUbwihvw9ewn3Nn1y/3VsXu+nwO4pTyfJmJAD4z7lHOQNfqrftBUGpQtmTh6/cOaUCda2uKYp0mbItG7F0oWe9kO93AWLlixbuWZdCJg/e3Rqw3vQru3f+48YP33CX0OVd4ldH+5wDsp4dN2gIWCSbTKfSNYC98hyKXxG/+Q6SCZEYSmNpayUYiZ8IRgIqOOzQACdYDntsI/V/+WlkBnwoRRW+2PQCZlKlgDf7SEqyKIgeE4wHVLktkTjfaVhLwnyC09hLJGSQLIYDl54YuyMGd6ILSTA03W3HAcla+GskAER/73t+EDOgQjxEVLAIdkWkWX/V7IvATJM8hjt2EPHg2jhjd3CNNC3j5AEn8aLZNwQguGREAUXTksewrpbRmx5LRyH8bnIQ52TJ4wZAgWi5QPpN/y5xw4ncUBGhIzxnrTvc/GJ48Gee8bTiOGMB3JOROnjmbQfXogHh7SH2be8NO7JsYdCjvA8spwfKUdsY2+SaMa1D0SOKmV0L1/J8IglbV4XMuN2hHDGXYgM6QuZKfpiHBBLkBX87wMzMlfAni2HFLwtwLugFDIrLku5JGWUFCTfuF6QHneFtLgij07sdcaFC0HLw+eyAmDUjEWrH4kJblX5bqJMw9NmypqDBQl8l7A/U+/VCGgEQhsCfEcaOnHuMszCm9aqWPrf1f+QlWbwvZ1FMiz2CG1j1uPRCGgENAIagbCBgCYswsZ10qPUCGgENAJ+CHz0cfwEo2cuWYux8sJZkyckT5UuQ/2W7X9fPHfapEvnz50xQ0Vw9bEEBdiXp1Dxb3uPmDDDIcvEr1+7erl0hao150wZPwoiAQmhrgNHTiDQP3JAjy5fy6qofEVKftemW78hDSp/V8QKP1kTA8dNX5AtV75CBHLv3Lp5o0yln2pDAPzZs3Nbc/2UYqbJa0VYEKwfMHrqPFZWElT/Vgy561YsVWDH5g1r7S5zpuy58g6eMGsxwfspY4cPImDfrsfA4aVypkH+xG+7duXSRdqUeHisO7dvEaDz20qW+7Ea5cjBvbvVyq8//hw9Wdoi8GfkK1ryu+LZUiWmDV6DR/I06TI+FHaE4HNsIRYkweLUJ59+lohV/Iz7+pUrBKxeactdsFipNOKLIXLdT8CcoPs9WYqfLHW6DKTE0OdzYRGOHT6wD2LBqZYuG4Fyu+wSNQgyAbg32jaqWckasP8qWcrUXDfOZ36Dxs1YiCEi8/oo3sfxf6haq97rEBaQUvWat+8yOgCD6e9/rP4zJNo3yePHQmJJjZtzm7bv2htJK0VYYMI6ctqiVfwYpl6kyJEi92jfoqEV8DZd+w2BgJs2buRg5la+2s8Neg4dPy1v6kRxFNHzShfJdRLvBa4H5EDBEt+VQ5uZ9xT3AfcmBIkVa8ghJL489a9g/u17DBj+XcVqtdRYHwlArepXd96f5g1cuJchLNzNq9ugURM/T/J1ssol8jh9NPT2ZhGw8aPwlUA2ny1cX+Ru1kkhS4INUovsi0ZSICbJnKBATChPiqPynIB6bSkfS0njOhe/jE+kQFwgC6UyKpApIjOAz0GyKQ4KuxBHHj+TclnIh51CHOyXoP/p28+MRyLDdC5qOOO0yDrdkdcPJYPiUyEBogs5wXsUIsXplSEEhPrMjSDHkKKin6+kLQL6ECNP7z83wj94ZHwt/fD5eFci+dQjEYINiSqIAAgB5JR4b5PFQJAfsiCVtEt2xhV5hCy5IuzBhz7PnWPwlvKeZF8wf4yy+VT8gOQO9guZwfngdm/dbcfNLXeM8B9HNqIlj26clQwPXzwz8r7ndU7Ij9uxIxg3hbTwkbFlFWLkQ3nk/yZYpXWNC5Nvsiz4naQyLrg2FMaaxFWog9wXxAWkBRkvjBPPi3NyzRk3xVeTF4KCbFGjRYs+SL47sCqgXsVSBS+cO0PWinPLkCVHLv7nqe8sar9+1AhoBEIvAh17Dx6VRhYLNTORFYw2vbyf+U62b9f2LaF39HpkGgGNgEZAIxCaEdCERWi+OnpsGgGNgEbAggCBzX6jJs/5QDIUapYtkouViASiZ6zYvA/iwkxYEGRn1fl4yQLANLrvXxNnHT98SLImKpdF3ogV4kriKEeegkXIkmjXuFblpfNmorFuNBASxMfnmStU7n8g7XsOHAFZQf1l82dhJmsQNK78c4OmIwb07GKWh0qbMWt2SYq4433y2BHGykqsc94nT9QqVyyPTCfi9OUb90iwvL4dYRH/088SM1/q1y5fIh9EhIz9TOvf+/wZS1JBzHI7Eut+ekOW4lvJCsaWOn2mrDzu2vrCg4JxQlZAziBnVaNBs9bf5C9cfO7UCWjLi0vswwc1yxTJ5fzRJdkVkD19OrX6Zf3KZYuC46Zk9TyFtsj+WLbt8LmpY4f/ObzfH53ctc+15wfg4F6d29nVYVX+7wNGTIgaLXqM4+IXYq2TIWvO3ATw9+7YsrGnZNJkyvZNnr5d2jSbMmb4IAgMX1/HaxnIYqzOqv6NpkwV8xg++TRhota/9/6T1bRmsoI6SZKlSMUY1q9c58SXVXl9JJvl6qUL5wf+0aFV2+79h+UtXKK0lbAgGyhPoWKlIN56dfwVTwBj55Z/1xX7vnzl4CAraO+rZKmcweGH9+/dGzh22nxWD3Lfk7k0adHabT/WrN/ESljgX8E5B4XkCOx+4br2/WvSbOax7d+1q/r+3q455F8RIeYaturQbWjvrr+Z28jyTd4CEITuZFMKlfz+hxJlKlRR93Jg/evjbwYBF4kBccHqcTxxICm+dvVeUx7JZJgjhfdhMilkASDfxDGIib1SyLIgU00RFirDgsA5pAGBdkgG2oAjgDS46ONrrJBAP6RDgms+xtbDDxx3kUi6/tRwSPbBbcmquHDpqRFHIu73JbD/RAgN6pJpQEYHmQgE8wkssx+CgYwP5KkYI/0hpwSZwbFo0jHECX4R9+Q57ZA9AbFAFghjg1xRPhu8pi6EA+dfdX0QJZTxRJLzyVyADICAQaoK0gOCASKAfpgz/6cYw1kp14W8eC7MwvuPHhk3LjxxXJLsEfEAN6JdemLs/jKqEf79iEb4DyIYRz+K5LVW5KaySFbGefCQc5kvY6MwZkgY5XdBBgnHmbfaNsoTskSQjILswF+knxRIjoxS8LxBPuqJXHfIHXVdTE28eBqY6fpLJ4TRHdXr/fIrGWtNa1YsbSYrIOaz5spXcOm8Gc7vH3rTCGgEQj8CLNog03vSqKEDrN+Pc+QtWPTU8SOH+P4f+meiR6gR0AhoBDQCoREBTViExquix6QR0AhoBNwgUK1ek5assGbltZJNINBL9eeyVN98GvJBBLF3b9/8LwHqY4cO7K1ToUR+Jcdj9mNIkDARQRfj8oXzBHyc27C+3TvaDaNAsW/LfPtD5Z/GDe3fU5EV1COzQsiJHFYvC8gSVqcLLxCVwCxB6DoVSuZXZAOrKclcsOvrt15/jiSg26zWj98pIkKmaztfpJ0O7rE3OJbMgwyXL54/d3j/np1kMzRo2aErHhAj+vfoTCAdwiJuvE8IUr20kWnBTknOCJG0doge2seUPKAbP0Xa9JlYnbrfzWq1oqXL/QghhNwTc7W2lTVX3oJ7d2zdVLJspWpkeJjJJjuppaC+CTMKAeI0pj56iNXFL221m7T6DY8UyAXrQa4P+9YsXzSPx0atO3WXBIXYtX8onpcMkPxyz5UUCS0yHcwZJvETfpaY+ub7dtXSBXMoQR2/u/pfJk2W8sa1K5drN23d4ejB/Xta1ateHjIEwoB7F1LNem6KNBkykS0iUBBkDnBr063vEMiKWZPGjuzRvnkDfDLu37tzB0IRosxKWIAz7yc7Pw2Cfg1a/taVDu1wDmws+njIIyCB6WcSvN4sPUGiDpaiDLmbcutLmSyF7Iv1UgjWE8Qn24JAOQTFUtMoITkgMVj1/0iC+wT1ee/fk4yKC0I+XBZC4qQE6jdKFkSMB5LnIB4UF1bccES6+9x4/ui5EV2yJmIKG/CR1OVzFQKAQD0EANkdECGQJkiTQU5gcM17lX2QCBANZDxAGnAuAX1IDY4zFkgKPB4YP+1DMkCA8Jz/V8gsUZ9CfQpzhCQgI4SAP0QMmQspXO3TF+QG0oOMgbrINEEusJ8+weM9mVOcZ8+NSzL3ByJn9XDJdccD3LfFb+Pxx2LsnTKGcf7bD71OJ4jilJp6JIN/LhkXZE+QtcI1UNgzLjCAiLhF21LYuD6Qk/z/ZE7UJ6OEa/WNlBlSII4gKrgunAu27HMlnbhaekceSpT9sSo+U9ZsPgh0FiFsXrcK6TS9aQQ0AmEAgRJlK1blO9mEEYP6mIdLZmxWWVwxc5J7edAwMD09RI2ARkAjoBH4jxHQhMV/fAF09xoBjYBGwFMEWE1es2GLtgSkVyyaO1Odl1RkgHguq+r96d0T2CSgSvaE/HaIScaAnXcA5yoygGC+sd39iJAUatm550CMnf8a1MsZGFXbvp3bNlPM+zDChgxZMnf65EatOnUXTuDTSsXzZDJnRiCtY7cCiwwOfDUG/dGxtXklZtJUadKTIWKeC6QG+rmjBvXpZh09gV+yGGZPHvcXx5qK98fNG9euDuzeoRWvOTega5AqXaYsZK4QtPb0WgWlHvJBL67fgQAJC8gg9L3tiA0C1bV/ad2BdtQ8zWNAKotsmxl/jxrWuE2nP8YPH9jbTDYFZbzu6jK+Y4f277ULpHMPlPqhUnWC+Pg+WNuQJAbnPcy9TeYCsk4E7yEr/K6RkBXW8+7ceiH95bxvQ2hDbx0z92Qp06YvVyBLKpW5wY/0Bw/u3bO7d8mwIJvJnRG9Gmr5arUblK1co87i2dMm/tGuWX3axFul2HflK1HH7KvCawhIpMSmjhtBoPulrZiQVviucB0C8rcIIah0sx4gIGSFuo+RF2ophawiTEm5h/leXt3VTAFTcwTxnZtEufO5nuJHEU04CG95Z2yVx3gio3RRAvK7JFB/V7IMvEWe6f6JR46rm24bl84+NsLdeubwve5jRBPzawgFRSxAIDAWMjcIphOsJ8BOAJ7sCQgHxoxHDOOAICGbgSwL6igpKjIMeE1dZVatsiIYMn1ABrCRdUHwn3oQFwTy8eGgX3CgLn1DmEAOMEbGS1YGdSAnkDqEROE1xAFkBfOCVKFdSAwIEfadEWKGVb6YhceRDJJHku9wVrIvHm254zifOIqXj0hHPS/7kdca8b2AIGFuZEtwLp9N9AeRAwbMlzFzrbhGEBtK3kueGs7/K64N8oT/qHy2q+yMC/Kc+UHevFPEBf9r+V+wcvE8pxeUeUMuEOJ8y4a1+LnoTSOgEQgDCLDgBlnM61cv+5NI5TsMi6nWLnuxCEVvGgGNgEZAI6AReBUENGHxKqjpczQCGgGNwH+AQNkqNesiuTOsbze/zAdWrOMbsWvrxvUE8c3DQgaJldoEf7u2blIHksHdsLdtXLeKYGmuAkVLKEkou7po7H8c/9OEmBp7ojOtpJjwgqjZoHkbyAdSxFXbtEWA9uzpEy8Ze1er90tLfghNFW8CVT+x6PIXLFa67Jghff8wj4+AN9JO+3b5J0yogwcBj9s3bViDCWChkmXKt6hducwTmQD7P0mQ0BnsRmbHbs4ZsubIvXvbZqeUVEhsn8kPPgLbynjUXR8Yip85deKYXRAcCSAC1QTP7cymycqhXTIrhKu5MiIA6alXnSOB9BWL/0+kmdup06xNR4JVEBI3xUDF2kfSFGnSeZ88fhQPkV+FECOTwZwhACFxV+TArP4d3PPgljNfoWLW7ItXnYf1vC++SpoIRO8tAAAgAElEQVRcOLVIyHVZ32N2fimQR3iJLJ4zbVJAY0DzGZN1vF06t2xYS82t2Hc/VFIZT0hEmduAzEEuy07yi/dRnaZtnJ8NAb2HgwsX3U7QEXCRFQTdCYgTDCfITiD9VykQquwzbyfkxQPMreURs2vYgF1CTtyUx9gSqQ8v+7x8fY1wYlx9WAy0j4ovxU7xosh98YkRafVNx42tdx33rz41ogmZEV2C9QTQyXYgq8tbCkEmAueQFGRKkLVAtgBkANl2kA9IPXEO42Q/BC+FoDtkAp+fyCUxL0gFzqFQF0KR4D7PlScEJIIiHhRhwWvIEkpiKXwWIx+FyTVkBP3x/wvZJkgQ/EAgJmgTYgHCgEwLJT8FOUB2BvVVlgqkA0QL9Wjj6YPnxjUpoiHl8Nop5t6b7zgeNPzU60y6mF7JZQKPBa/lYuaNfwhEBVkTzIdzvV19Q2IrEob/YZA5zDeTFDYMu3NLIQjf3jVO5kw74EmGjCIuXKe8vQ9kgfL/i0wK8yxZbFC45Pfl54gko/q//PaioGemEXh7EHgkWbX8LuH7B35szIzvKD83/rX96eNHD5Ph/fbMVs9EI6AR0AhoBN40ApqweNOI6/40AhoBjcArIoAME3JASrue1Ut9RkycifcEAXhzs6zEloXhqSA0jh85uN9uVbu5PhJCWzasWZG/aMnvzd4W1qFW/KlOIwL7y+fPnubJNFIJaUIgFmmbk5IaMFlMs83nfZU8pVOLHbkq836MxSWdvOAEyQRQAQyCuEMnzll65vSJY2QImOsT/CX7wM7kOGmK1KzONfbt2rr5l7Zdeu7etmnD2n8Wz1fnJ5KINM/xybDOCbkfsjOEsAixH12fCdMgMffjdpkJ5vEgM7R/93ZWQfvbXphdt+vMzi3rV68gi8FaR5E2EES/1qv2g3h9E8gLtg2cyOIgq8DaKEQKck7styNTIBoY38ol82Y5CSkxtkYyzIxHYrlG57xPvXR9aHPutL/HNG7d6Y9cBYqUCC6PETUHjLMxtycDaZolq4H3H++vC2dPO7NA1PalkAocc+cxQT1+3P/Wc9DIx48fP2onBunqmkF21HFlyvC+UUb1qu0UadI7A6HWbCr2lRbzepWtY4dzsF1s3VCQEXARFQTM+d5NcJ4gOkHb1FKQw8sjxUpW0E8SISQeibzTEQme7xTS4Y6YMRyWhiJHD2+EE8LCS/bdluD6vctPjVM3fRwRDz0wIieNZuydcMnhc+qREVfqvC8EByQBGQ3K6wGihOA6hAWBf44hUQUxoMgCMheQYVKm0xAaSt6IgDtEBRkXBPMhVJQclAraQ14QkIfUYJ6QGATpIU0I/kNIKFkoZU4NsaGMuPGroD9ICY6z8ZyxM058PiBNqEcfSh6LOUFikBnBXCBhOMZYISwgqhkvpA3XJKJkX0SQnp4ef2g8bnPC8bDBp8aeoh96Xbr/zHj6XkTDRyZ2WKSiFH6MgblBOpE5wXjon7Yge5B+Ym58xnKt6RfihefrpOC/wXnMnfGDMzJhb72/BZ9peADlFgk8PJUO7du1A6Ptzv2GjSVzzSorI7joTSOgEQjFCGxYtWwxXhWVatb/ZebE0cMTJvriy7Z/9B/GIpO28t3GusgkFE9FD00joBHQCGgEQiECmrAIhRdFD0kjoBHQCFgRwGeB1Ouev7VE49zIkjNP/vY9Bo5AYgnzSkgJ8zmYWhJMZd/YIf16ePKjARIACaZKter/YtXNpx2yJT6X1eYT/xrcz9OAd+p0LwiLtJmy5vhZTLYhFczj/Cr5C0NjJGzM+/FbgHRZPGf6JIK731WoWrPZb936EDhuUPn7IlbPBQiLYyKpZDVzps2kKdOkU34dBYt/V65muaKsePXb8CjgxakTR5EC8bely5wtJzsgOULqruS6Wudv7Qs9YH4AEpy3HitdoUoN5aOwd+fWTXbjxNuC/WQxrFoyf3Zwz+XLpMmdGNr5V9Rt1rYTgXiO243v00Sff8n88B+pWrtRc4gzswE75vFIi21YvXyx3bhnTRwzombD5m1qSAZPcBMWkC30+c/C2dOt95wQXbbeI3ipcE5AhMWPNeo25pp0btGgppK94pyylWrU4b1L9tJ1kSCThBmCyaZ7NXlKAntn5UKa90NasaKRfZxjzmIK7mut2/McARdRQaCe+5+V9QS3KXwG5ZJSWAqBbOemTA3M2mfyPKoE1B/cembsFoknAtyJxY/BRwLoe0X+KbU8jyTPYwpZ8fTkI+PRmluOj+dcNRySOfChtEfQnOA8WRIE1PF2gCzhOf0TwHfKqrnGSLYAxymKnCDTAlIFMoFCYJ0x81kOOUHGAdkPEAeQERTIF/ogyK+8LuiDsUAgIAHFXCAwlHcQbdAn2RyQIxADKpuCeTg/w1znQGpAwkBOeEtBVo99TmNx1yNEAeNgjhAJjIf+yM5gP9eD/jjGXE4jpSUYxx1w1nFu8x3j8ieRjejF4njdihtJOEYvw1tIIi95VHPk/c/YMd4GD7JU+F2lDMSdn3mmDU8LCuTLP1L4n4JPCfirzA3G8ZJMlNxHb40pd5/ObZomS50uw5hZSyFvnBvkdBfJMgssy9CCp36pEdAIBIAAnmexYr//PlmtSsoyuAGbNWncyG/yFynevEP3vhTV/rzpE8cGt+xocI9dt6cR0AhoBDQCoR8BTViE/mukR6gR0AhoBAxWIwLDI4nIj5m9bD2rEvE8qFwib2YyF6wQIX3EvhvXr15ZsXien99FQFAiP4O0VIXqdRpiqG0N/ucrWup7zv9n4RyMRAPdWDmfMl3GzBAPeG7ssgn6i61CGoIVJyxGzcyXsSP1NGj8jIVkV9BGtza/1DX7X6hBpEmfJdu6lUsX2g2KLI6jh/bv+bFGvcYEw60+G8jsEOQ1GzerdlJnyJINmSXr+AKdvIcVCOR/mijxFysWBYwpYwTPM6eOI0/itxGortmoRVsCPQT+97kx5BZCwXk/TB8/cogn5JWHw/erhj8GL7wt4yNjonCpMhUYH5kKkErWtr92kVZIlrXo2L3fz2K0ba6j2nZH6nA/TB49dCBySOkzZ/8mOCUIGD9j2frvOn/STOxTxIR1XLI/A8GBE0fszcfJiKrXvH2Xw/v37jJnPpHNUb9Fuy68r1/IpPknJegTLM57nz6ppBcUTt+Wr/zTBx9++BE60qK4tj8krnFQ7wld34kAQWuC2QThCVYTjCaw3k4KQXiC98gZnZUDnzkZAlnpLxF+VuhjEO0kxUSW6Bsxjj4oEffTIvn0fqTwxmF5XCGNf+sV3kgg++Pc8DGe/n3J8VS8KxJJO6z+p32aZCU/QXYelbQR+yETnP4OUgiUE8AnAE/gHdk+shiQb2MOBP8hO8hYcBJyshFkx2eC86kHwQA5oPgWCALmCqkBOcGm/CZ4hHCAXIDAIYgPTmSdUBRhwpjJiCAjg/GRzaRIB+aU2HWM9sCYOTNO+mN+ZFrQP/upwyMyTjwyVjVH5k82CWP3EYIowYbbjiuC/32R1bqUObbX3RyxjXBxI3ndlOyVWAKerxh3l5AJ0gaeFIyX9hknpDFjRQ6K+YELG8QPWSlccyT6IIyYHxjSL1l8ZGeAhVNaJbRuECiujWvM5itm8h4Nl8/5ikVypsezgs9KMjYXzJw0ns9DjxrQlTQCGoEAEZCE1y+69B8+Tv1u4Ds233tnTR47coksAgrO7wdkhzapUb5U0W/LVsyaK19B2l6/YunC1csWztWXSSOgEdAIaAQ0Aq+LgCYsXhdBfb5GQCOgEXgDCKTL9GKlPz9CWJHdqXn9GovmTJtozVhQQ0niWlHPjxNrcDOg4Y4Z3PePoZPmListGQ1Tx47401xXJJoKENgPaOW4uX7iL79ORhCW/gf36kKA7qXtaxGvJjBr9cNgvnE+/Chet0GjJkJ0MN+dW/71W5FpbohAOBkoe7ZvYaWrvw3vgc8l6Lx3x9ZN+G80rFqmmLUOQWB3wXB8GfihF5w/8Mz9Q8RAOuBNEdB1SZAwMauADWsQ+7uKVWu+JxpeC2dNnlCm0k+1j9gEfWgfDAiih5S3AfN4IMyO1Z+iXrM2nbhfHkt6wtXLFy/Y3a9fp0jl9Bghm2XHlo3rrDJI/ycs/MuGmfGaMmb4oKp1mrSoUqdR8+AkLJTEElrM1uuTOUfufGQa4bdhPvZ1ytTpThw5fMBOmot61es1aYnm86AeHVub76v6Ldp3QY4Nv5m+f02ave6fJQusfYIzkmjm/dzjZFew0rF89Z8b7N+1bcsb+EjSXQSCgCu7gkA237XJLCCbjCwCSDCC8mQHsMq+tATA70h5JvJOEcQQe4Ks4jce+xqXY0UwikpgPL28jPBhJCPpmUfG9bOPHU9lpf9D8VyInjCy8fyjSEaMRFG8PhQj6fySbeEtkXhFHkB2sNofGSgC4DyHfFBBZh4JqENaQERAVvCc+mQqMG7IBCLRPKosEepAFhDsZ168JgjP+QTtCdBDiHA+RABZGZAEYME4OIfAPG1AaBCsZx9ECGQDBABts9EG2R20Sz0IAoL+kBGMX3lY0C7jo03qQfiQxcE+CAEemRfjYj6qLcgPCA3OYwzMm7FRJ6Zcj2NiUv5g6XVHeDEu94oR3uFb7ROvK+JxEVt8Qq5GEVkuGQTnMG4ICQgLzmfOtE1/DaUwPuUBwjXPK4V7gM8+zMYhrQjYMw7GCiOgEm7kaejZTGQF2HPtIVjIhPF4YxEAmZoen6AragQ0Ah4j0H/M1Hny1fs9vs+LZcyj+J8l+jyP+Jd1G/jX3z9UqVWvZd2q5awm2R43blOR73VL5s6YTHmddvS5GgGNgEZAI6ARsCKgCQt9T2gENAIagTCAAD4KGFCTYbBm+aJ5gfkdJJWgKdNavmD29KBMb9O6VcuRk0GCyUxYEPQmsLxxzcplgfWt+kuV/oXR8+K50yfZ+Q9EihQ5MnJI/yya+1LGBvM9uHfX9p6/tWh0YM/ObQHNAbkpju+VaLe1HivkGTuG1Yf379mFB4i5Dr4LyA3Z/dDCxJs5I6kVFAyDUlcFxJFqCug84WQILBqXLpwjKObcGF/tX1p1wFsBSSYC53ZSXV98nSwFGKAdjqRWUMbnad244jliHhvnIfdVuFTZCo2EJOo5bPy02ZPHYSr80ga5xr1dsmzFqq3r/1TBWgHJLgL7Rw7s3e1uPMxLkTYBebB4Oh9VL76kv/Dc+uOezJgceQoUgQgzm8SSBSOeKWklq2mWXV9IX5WtXLMuJNjWDWsw4nVurISsKDJRZC/dFFd0spIunDtz2toGOG/5d63feRwvW6VGXWSzkMyq/HODpu6ybII6d10/6AiYJKAIppMxwOcwMksE3AnI55eivCqU0fU5yap4LhWmCFnxnvdjx0EfX8Pr0lNnpsOKxFG87ieMYnwmZERSISvuLL7u2H3lqXHrmo/xfsaYXpdzv2+kk9SCaN+855VRgutnp11x3Jb2yBbgM4PAN9/1CY4TDCdorvwmlDk2j0p6iTpkNBCMZg4E0gnIE0RnH3PiM4TAPAF1MhUgFyAQyMKgHu1Rj0ckzVS2B4FtpJ44h7rKvJvxUAjqI9ekvC9ok7EzZsgdSBMIC47TN+MEVwgHzocQYWPMZDhQGDN9UhcsGAtjU3MEF64Hj7TLGCA2mIciMGjvgZiaP5PyWOSifL+K5rhSOq7XKsE8bozwRhzJxKA+RAtZEiqLZrM8BwP6B1/ICcgMXnNt2QpJ4f8kc4Sw4H7Bq2enFPBSvhb/OXlhyaoAR66fIqaY538+Rhem+kEj8M4ikCpdxizITbaqX708WckKCLI2q9Vt0pIszkmL1myrVbZobrvvGO8scHriGgGNgEZAIxAqEVCrrELl4PSgNAIaAY2ARuAFAu9JQJLMilVLF8zxhDBIljJteqQXCPoHFcNFs6b+jQkypIE6N37CzxIT9L5oE0R11z6eFxzDY8CuDoFoAr8QCebjEBlo727ftH5NYGQF50FGYBpOsfYjSkpO3XOC5+OHDehlPa5W7x854H8M1BOf5+TM+dC+PQSPQmSDsCEY733yGKts3W4fxP0oHpkqyGeoSlVqN2wWPUbMmH/LStWkKdKkc2dKnSxlGsxnjZBM0Y8j47tx9QqrqP02PEcI6JMVwmo/d+PjxzXE0cVzZ73tZMO4Rhfk3mdVbkAYcd9yvSASgutiydvuQ1YPWmXIcuUvUoIxr5b3o7kvvETkmsQ6YfGUUXXyF/u2DKQF0gxqH9j8PmDE+CsXL5yDkFR+I/Je8za3jScNmRlmnOkLk+4pY4cNEk4LSRwxj7c3Jw8uTHQ79gi4yAqC4QTayaJAfomAdAcpraRkl6KIBNVIRvFN2CEyThvFIHvrtruOTYcfGBFnXTWer7xpRJpxxRFx5AXfE8tvOI5efWpc/zyqVwwyLy4+MXzlnLi77jmuShD9uLQRQ7Iy4nwR1UggxAaf22Q2QBYQ6CcAjucJ95MKxBNcJojOfh4pW6UQrCfrgUA/72cC0byGZGAjsE+wmvM5Rj8E1cnqoA6/K3hEkom2yDSAdED+CWwgBZTsE+1AFhD4Vj4fEBLgxz6yNmhXGWsrkoJxcBwCA5KC/iAg6E/JKdEGxyFgVHCdvlVhH3Nk7IyZ7BP2MR/aoU2eQyzgYwORkFlKMsE/7v77xnv9zjjudzjpOCTXZa3sx4OJMUBY8P+CjCx8pcAVaZTVUsis4P+xktSSp05SiXuCe4N7hHuFe4Z7h3uIeSjyh/r/9QaJg18I44LcAScw12TFf31ldP8aAUGARTDXrly6uGntyuVmQPj+iNRrwyplisaIGTv2iKkLVshXDz6L9aYR0AhoBDQCGoFQi4AmLELtpdED0whoBDQC/0cgljAWnhpd8yMEiST5wbLsVTBU0kpJXMF+2mDVOo/XRCPf0zZTpcuUhZXp7kiHr8SggrbQ7De3yVx57SNyO570lTZj1hzuzKaVNBYeFJvXr8bo1N+mCAvx2z5gPSaEBYEkIyQNjD9PkjQ5xNKD+/cDlNQgyP3w4QOkTZwbMlg1G7ZoO/rPPt2fSs4/hty0Y4dXslRpnYTFq94PnlwD6/hyFShSIluufIX6d2vfEqN22rAbn8TgoyUQvWWOTxw1pL9dX1wjTzxEIOeQvVLX3JNxB1ZHkliiPhIDbGs9TLN5Py5fOMdfBhPZLNQ9efRlXxn2Q3RAOCq5Jwi7XsMnTIdsaNOoxo9IrqmsG1HQ8kfAgTFtPHx43+8+qNO0dQdfh6/v+GEDe6u+JVZhex8ENld9/NURELKC79MEw5FhKi7lWykEuitKQdKI4DPXhXuJwLZzE8mhmeJFcejmM+PODR9HQiEi3o8dwYgpq/bv3/ZxhHM4jJhCTBy//MQ4dOmpwydiOOOD2gm8PvTycrYRQ2Sgsl54bDySFf5e0cIb738dzSvLl1GdfWGyrTI4+DxVMk5kRhCQh/xjPyQXcnOYf+OxAaHBPKivyBUC+RADKmOBoStihvZoh8A7AX5FYiCRxH3K5xrPIQboExJESSUxB0gV9pGdADa0RfAbOSfOoU/uewgF/gcprwgC5+zjEfKCOVE4h/qcR/sQvDzSJuPxlsJ1YFz0TdCdc5SRNiQGeCA7pXBjrmRFUAjUO7Me5Lo92n7XYZTZ58ucGT/tKlkqNUfwUR4gyFRBYpgzChkb81ZSYdwr3DPcO9xD3EvcU1G5x8hycFekTohsrv6YI/cEixAUEQTGiiwKkb51oxoBjUDQECBbuHi2VImR6LQ7k4VArepV/SG+yEsiMRu01nVtjYBGQCOgEdAIvFkENGHxZvHWvWkENAIagVdCQGLV9yR2SiAp0C1pyjROOSh+mARWmWwGUsjN9bxEjobXsiCLAJBzQ+qGx6gSYLa2mfjLr5JiJGzeT7uYXW/dsHalO/8Hsh44x0oWPHxwzxm8Z0V5YONHvz9Z6rQZrEba6jxlPj7z7zHD7doiy4MAstgCvJThoOSAblz7f+YAwX+yPwIbl6fHyeI4G4h/BW0h/2SWHmrTre+Qm2JKPnn0sIHK38IdYYE8GFkO7o57OtaA6r0Y32NnIJYsgDbd+g3BPwUJLnwX2H/VJpCOmTjyRxBbSJ1Z+4Aoo5w6dgQTYH9bGsmsIeCvdoaTFzx35x3xKvMkqyOKvPHM5+JdgbnkwplTJty6cZ0gpN8WL/6nziwHq8+EqpAibYZMXAsyNnhPte3ad0j23PkL9+varoW6hyWzydmGNaMksmDMfoUz92LlWg2aDunZpR3BCXBGGst8n7zKnPU5QUPAlFnBdYMsIPBPYJsV+RAHaiPzgQA5cmGDpfQUwmKnyEBdjRLOOHb3mXHmwH0j8qUnxtMHz40kkjkR4dYz4fmeGCvnX3ccXHLdOLHnnsNn0x3j02jhnIF6CILP1912fH3ogVAbQiII2ZEs9/teGYTAgAQmsM54IAwTU1eK8qNgH4Fngv7qtwDZDTwneM/4CZ7zuU+Gg7N91zEC1UpCif2ssOc9wnkE3wli815UfhUQChwHH54rPwo+55E9oz3GAlmgPlshHZR0ltpHpobKNlAZHvRDnxDpkARgAjaMmf0qW4J5QeBAjnJNmKvqHyJE9QdG1FNG2SflOZkn/C/dIQXyhfni18F8wOGD7Nt9o0t5PPWyA+IC2T4IF+YEYYLMFe1QeE47PaVwD3AvgJNfNqNrfNw7XAPuJa4hfb3RTAtFjEi/XDPuF7BBygu8zObm8lJvGgGNQGhBILDvQEi/jh3ar0fewiVKFyzxXbnQMm49Do2ARkAjoBHQCFgR0ISFvic0AhoBjUAYQABTZlZeQwSo4RLoLVGmQpVOfYeOMU8BooDXIrUUqJQR+vd/L1i9JUvOPGirG7Rfs2HzNuKR/ODA7h1+3hHnvE8TbHFq7Zv74vW0Zf/uLl2hSg3zfrwfkOfZsXnDWnfwUofgKunr5joPHzy4TwDbulKeQHgNGdtP9ZsineHcUqbLkJkxW42a1XG8HehjydzptmaArN6/K0FeshSs40Tzl31Ro8VwrmwH6ylL1u/MmO2bPMF1y2BMjtRXYO09luuh6lT8qU6jAiIt1O/3di3IKEBSiGN2hAD7wfHw/t2B3guBjSGg44/konGce7JTn6Fj3hdjkEE9OrVhX8xY7znHZ0eYcH04tmDG5PF25vAqA0ZuBwKBfhtk14R5KzfVbdq6o9rJvQGBtX3ThkCJOk/nyvuO+wAvFM5BBqpjnyGjyYgZOaBnF2s7cosSEDasRIaqh8QUfh2QFb/1HDSyXNVa9ZBMM/vFyO3sfI8r4k6dqzDmtSRRfdBr2Pjpxw4f2Dt/xiTnKknug6uWLBuM6z92kSiezlnXCzICBMi5j1l9zvdqgvyppBBwtm4EvBdLmSQyTuduC0mx6Y7jxpyrjkhSop5+5Hi6+qbjiazcj3/Dx/hAyIx9Qlp8JlkWhWVflB13jWdb7zgSP3U4fQ/wRIgqRIex5qZxQqSJblx+atz9JJIROV4kZ1CZFbbKY4LAPoF/gs9kGuBDgXk7nj6QtdxziiCgDsFxAv7UI/iuDLKVoTZEgJKDol2IOwL13lJUxgRm9LTBOFRWA6/BSPle8NmqZKMYF6QnffOZAY7KqJo6fMYwHqSieOQY86M+fVCUYTV985nBnLg+jJs+GTN9UHhOBgSBeIgHRQLxua+IDpW1ASHP/1WuM7jzSFYK/iQQDk4ZrT/POYyfDvpChDBfPHeQO0R2C48ixgPm/C8Fq0lSuBe4J6wb9w73EBiAF/cWfb60YMDm3NfeZTHWpl8IC7JoGAtzQGbMLwMyfULnx57eNAIagTCCwKhBfbpdlC+fSHeq77phZOh6mBoBjYBGQCPwDiGgCYt36GLrqWoENAJhF4Fl82dOlVho7I69B49Co//HmvWazFq59UC3QaMmWmeF/wReBwRbA5sxRsxo9BP87D18wow5a3cczpmvULEhvbu0N6eUk2XAqiyC9azuZwy1GrdsN2zSnGUSu71LwNncV4o0GTLxWuKp/vwpzHXQ6hcu4SW5HeosnT9rKpJCBKFz5C1YtGGrDt0Wbdx/qtGvHbrdvH4NXXPnpjIoUqROn3H59iPnCeSqY8gNyWL1REvnzZzizv+AgDgBZDuczpw67sSvZace/Vt26jng9/4jxoPXxjUrlgaGqyfHCTBj+O0JYXHW++QJZKD6/jVpdqvf+/zJ6v51K5YsoB+VEcN1sPaLVBQSYXvES8KTMb1qHXwTuF4jpy1cVajk9z9glq6IKMZHlo3wUC/JXiGJxf3nzpBbERbWa3Ty2OGD9FmrUct2YDJ58brtDVq2/x2fjm3/rl31qvOwnse9wz7ed5hiQ5KITcUXPTv8f37mc4T7cnqMVKv7S8tM2XPl5bxVu09eIQOF/dcuX7qIt8uCDXuOl6n0U22ySnp0aNnI3IYyze45dPw0M0FJVgYZFOWr/dwAkjFuvE/id2hat7rKYAJn8z2QLnO2nEu2HPBevPmAd+FSZcoHFya6nRcIuCR6CCAj34PvAKvi60mpLoUAr5PwNG0Qs8j0QQDcu/fc2CjZEydE1umk92Pj/IUnxg0hMFafeWzEFZ+E6JJCEEFSEfis4zxv2XdFMilu3X9uRBVTbrIAWO2OrNG5C08cm0RG6lqiKMb7WWN7Jc8W2wtSlTqMj2A6GQm0xWcExACvWbWPxw9knJJYIjMB8oFHxu8kG2UjuA+pC2mgSHOC6SpjAvKAwDztKmNtAvS0BSF70NU3vzsUYUKbiuygDoF7iASOM2c+lyE/eKRdlU3BeHg/8XkCocAYlP8E5AHPIXQgIuiDzZkhKBv/b5gHbYELmRbgqMytqUdgHhkmsigySAHLElIgECCCzkjBswJ8IDyYAwVyJNLRh4ZDsi282p90MA+IC3BwXkPXc/6v4GfB+LkXuCf8kfautrmHuJe4p7i3uMe417hWIfL7zZRVIV0458N8wYb7gXsNbw6us1O10mQAACAASURBVMKVenrTCGgEwhgCLNKZ+Nfg/vhuFS75vf5+EMaunx6uRkAjoBF4VxAIkS+87wp4ep4aAY2ARuBNIbB+5bJFBKhLlK1Ydeikuctadek9CE+DlnWrluvSsmEt8zggAlYumT/bnRSTuS5B386/NqyF/BKB5of37937tV61H6aMGT7IOrfeHX9tclWE9StUr9OQMTRq1bH7sUMH9tYsUyQXGRHm+p/LinT6N5ML5uOsMGeT+K4tWYBBNgbfTdp07jF04pylNRs0b7Nnx5aNVUrlzbJg5uTxqi1ZIUbwyPi1c8+B+AkQ0FXHokePGZNV/aMG9e5md51YjY9fhjtSZeXi+bMwjS5autyPlWrV/2XF4rkzW9WvVt4TXD25L5DSop4nJsmMhbmRWUGQu3u7ZvVVH4oYKF+1lt8+dYx7gcyFtf8snu/JmF61zpwp40fFlvQBMm4G9+rSznyNGB/X+ocqNQm8+duQOcI0nJV+dn1/GC8eQVchvvybokNytKpfvTyZF2AixE+84f3+6MS9+6pzsDvvyIG9u2dOHD08febs37QWouijj+MnAHsMvu3q/7Nw9vTjYrhdv0W7LqNmLF5T6odK1ZcvmD1NZfCADdcRs+xxco+3qle9PHMxtzV17PA/8RvJkjN3/hixYqlV7wb3HThDSEJ0taxTuSzEzf/vg8sX06TPnE1JwkEuQpSQ9ZIhaw5/mVHBidG71paLqCBoz73JCntMiMEX4knJ67Gi3ynt5dr4XOoqBfNlgvCPb/oYlyOFMx7tumtc2XbHce2WjxFTSImIEplX7wUC09zPmMjHEfmoqFLHS6SiHkkdsiLwQ2CVe9wrT40sYsAdU7IskJPyFR+LGOG8nAFx5TEAGQBhoQL1ELtm02s+h/ksJQjP/Uh9gtQqKwE/FeagJJEgLpTUESSdygSADOA5JICSXuJzDj8MlU1BX2QZQHJAPCA9BZ5kReAzxOp96jAOcIRkoE1IC14zB8ZJX/QNCQOmkCM8coz3DVJTjBvigL7BkzknlgJRAQa0C+nBo/JpYExc27xSwB6ygAwM8FAEELgyHjDGIwhyA9KC9uk/kmTKhJfMA18pkChmEoZ2+H/J+Bkv9wT3ht//LnnOvaNkqbinuLe4x7jXuOcYH5gF2+84U1YF+IJNLtfcIXDYR1YInzd+n1dkVujsCkFEbxqBMIjAAsnOxDerfLXaDcLg8IN9yGSasDAs2BvWDWoENAIaAY3AKyOgVhy9cgP6RI2ARkAjoBF4cwgkT50uIyov3iePH3UX6C7+ffnKZAKwItvTkRG8F+WjmGRmBHQO/g1Zv8lXULiAWKckWHp4v30GBYFdvvgHZFiN5v5TcS62SkKp/hlT2kxZc0SUJ0cP7d/jjvxgJTvZJO7aCWg+ZCCIhzG/2dxiRXAYWanAjLE9xVrVK1elZt32PQaOKF8oexqC3IGdjxwREj/mILU6h5X8h/bt3jFr0tiR5nZYPYfs0oZVy5EeCdEtYeIvkogP9WOr9BPj7tJv+Lhxw/r3VIbung6EgLsoGiXifrc7ByLkgzhxP7ohfh6etvkq9fCLgBQBY3cZOapdpNC+Sp4iNY+njh897M78MrBx8OPZKpMF+YAc1vkzp09Z24VUqVq3cYvubZrWAw/ef+hTCycXZ+60v8cE9t4ObDz6+AsEJLBL0JqAMSvuecwnpaQUs1wPAWpWzqMPznt7oxSkyih3jjwwIuy+53AsueGIfOKh078go6sQxCfATVCawAnBc+5tZcBO8JggOXJ9BLCTiF/F7ZTRjQ9LfOiVRLIsjERRvaIdeeA4P/ic44CQG3hHEHzmkXaVQTRTUZkFEASQFaymJ2OAfiEJyFDgNefRJwQAwXZloA3pQCAfMoAAPkF4JRlFUJuxqz4gBVTQm33Kr4I2CbwzRzLXGGt2V12C8fw/AmPGoVb60xc4cR7tUDhfZX5AHHAOYyXIDplApgjnKwNuJfvEdVJzoh7jZK6MlevJc/ois4BzIRK4nhArZKfwnPlAgKyXAsGjjMUZ/9PHZd6jX79N7h/a5hiPHANv7iFKTle7eFsUleKUI3RtXJNFUriHwPqA69GZpfi6xIGLsABLpK+YG/elynzh85dsEUga5/a6/Znm9UpP8c2avXrbwXaNa1WG4H2lRvRJGoEwggB+E2Qa/1AwG+/NQLdi3/1QiQUrf/bs3DagykjKli5fpUbJHKm/cLdwJNDO3pIK1ev98iuZusWypUzk7vfGWzJVPQ2NgEZAIxBmENCERZi5VHqgGgGNgEZAI/A2IQBZgSxQ9q8/jm7nofE2zVXPRSMQ1hFwmWsrmSQIBQoEoT9TdtM8B8pzMhEIdG+XAslwl1X3UebcJmBNWwSkyTAgAwHCgKwE6hOoR0oIv4TPpJA9QCYB8k2R5Mv7XiEq4kcPbyQs/qHX+9U+8fpKyIpoQn6cjxnBiLb3nuPchEuOu2cfv1jtL4WV/wTSVbaCCpgTaKc/2lem1fgnQAoQ+Ie0IKjPeJTHA+0QaCeYD0mgDAyQDCKLg7qQFfQLccEcCeRDOnAugXo2sijoG6KAviGNec586RPygD4VkaJkiQiaMw/6oF3GyZhpl74VscBx2mSu9K18MGiXcfPI2DjOWCA1aIOxsEEk8FxlqnAt6QuiZq4UAocQB7QD4QSRoLx2IIHAHsKCcUN0uZp96YH+lYwV2RzcT/TT1M0JzK+uFPqggPszua/8yAR3HQW0X8ZHv8hfQYpBVnAPIDsINtdet/1XGVNA5+QvWur7fqMmz6lXqXShrRvWrAzu9nV7GoHQhEDXASMnZJasy6JZkpsz99wOccXOYxdZzJE96ScxAvp++U3+wsUHT5i1uOdvLRtNn/DX0NA05zc9lr4jJ87KV6TkdzmTx4/lTq72TY9J96cR0AhoBN51BKz6uu86Hnr+GgGNgEZAI6AReCMISLZMBrJkNFnxRuDWnWgEXhcBgtuJpbAKHp8GpI7syAqC2AS6yRhANkkRBY9U0JdV90JaEPSnEBhWwXiC6gTtCfyzup0gOiQFq95vCkkRTkiKCGljeMXLEttInC6G15dJov1feipBFCPCvnsO7z33necSzCeYTv8EucjS4JFgNJkMBL4VoaGkmdhHRgUbY+C4WtzklLKSQgCb4D37lewSQX36I2jOceZB5gH9gAX9ghVkBB4IEAgc3+d6hBxQRAn1wQW8nX4fUpQEE8F9xgcRQlYI7TMG2AD6BnslM8g1oj4YqHlBBDBuzmc89AXGEDfMSUk+0QbPqU/bXB/GTT3mmc3VX2JXe+AChkpqi/lT7st1fsb1NmckWMgLlbHyr9TH84lxcw+QYQEuTlk808a4i0sh6wFCi+wdbykveQRZzrN96SLiGPsXrn4hi5g/WSUQIk7CJbRtSVOmTseYTh79vyxeaBujHo9GILgQwKPq5vXrfv5tAbVLViueZ9SJEzduvEvnzzmlU+227Zs2rEGWEjLkXScsyF4lg1mTFcF11+p2NAIaAY3A6yOgCYvXx1C3oBHQCGgENAIagSAhgOF28lRpM6xaumBOkE7UlTUCGoEQRcBmJbzyZ1AG0yllAJgh+/PtkdcE3wkM4S/BKnxkipAkcppc26xQJ1DNMYLmkAEEYAmOkyXAsUQSbf9AwuuOqOGMiJ9ENqJniOn1XuoYxv2csb2+ixreiCOeF08uPzEufhTZiHPvmXF0213H7omXHBfE7+K8nJNQCI5Y8lx5LxCQJrhPcJqgPwQGQX4C9irYzZxY7c84kBxKLAUigY2APuezAp+ANsFsCAVkoVRwn8A9/ZBpwHMC/vQBaQB5QwCeLAZl6k12CfuYryIDlH8FmQNgCEa0Qz/gpOSrwIm6ZEtAbtAn+7hO+EGY+1YECH1T33wu15dsEEgRiAyO86jko8CC+VGHgCGBQIoib7h+HANHSBhw+h97ZwEgZdW98XdqE3aXXToE6e5UUVRs7MbCwO5AP7FRLMQWMVBUUBFEEFEasRCkU0JAumt7d2a+8xvmrsMw28Eue+7/f76Zeed9bzz33pE9zz3ngZghhZIvXVNwCZFOySvrjvaoE2zoJxE6RNxAWIETpJUpiIEjBD5cDAFvlz/VlBEPz7VNP1HBffT5IrH1YoyFyCGEwf/y9yXUEI76NbR6SOUYrJ911DumHVAEigGBDMm3abNlkcc5tgBhYW5wSG7JnG4m3em6tatWNhZnfTF0u8xUSbrb2nWPb/D96JH8pmpRBBQBRUARKCUIKGFRSiZCu6EIKAKKgCJQfhDo0v3UnnaHw7Fg7h+cqtWiCCgCRxmBHFL24ADHIY4T6Eaxu8RwchvNBNNzHD7GyYujGkLgYB5S6WQ6bVZqptfaFeWwwuKdVmq43apaPdzWtnUFq3ndCCu2QZStau3wrNRLgUjZJAVU/OKD1kpJAbXu7yRv+L5Mq448H1M/0tosuaP2ikI3DnSc0DjCIQBI84QDHuc75IQRs6bPpIbilVP8jHGBGJEkRsuhmbwnioDPOOSpAy0Pk44JogBnPfXj6OezIQggSYh4gMThGgQBEQK0Z0gVo5dhxLAhHXiGfq/318dnCAIiRbgOscFnI5bNZ4gU+gkxAeHBvdxD/bRLm4wBEoX3kCWGUGG+eY7nIRBog35CHKBZwZiIYKEfkAxgSEQEnxHQpg0IGvoA8cH1w3Qs5HOowjwYIW/WDusJXJiT84MeqCefGQ9rkfF84P/eaHJk04QvNZUhaBgnJBAEHMLepLWCbIN4+1ksJNmSbcUl/EWT5q3brsmD9lMJd0ubUwSKBQGRe0urGBsHKZprCQsLz/pvEwptuT2wfs2qlaSGyu2+Y/n7xs1btUEjbNnC+aRv1KIIKAKKgCJQShBQwqKUTIR2QxFQBBQBRaD8IHDy6Wcj0mvN+fXnaeVn1DpSRaDMIYDjBw0FnMdXi10bMAKc2TiNKTjhOen+uxhOXyIVEvNAVuDodzWOspxVwmyuTjHW6R1ibC2quKxoSf1E2qQciwh3r1940Nr8537vqrUpVqyQHjjH4zO8Vt09GZZLIixwoBMRgSMcxxXOaJzxjemfGI50HP28h2QgOgJHthHphlDlM4QH9+DshojAUc/YTRon4+QnAoK2+EyUCeSFT3xaDMc7Y4IcMGme6AtOOOrDuA5JwX280gZ1gif1Qp6YaAujkUG9fMd1/q7Bgc+4jAg4GHOPSdvEc0RmEL3AdSIzeB6igf4Q8cG99AfiwaTuom4wNKmjIH5YH8v89TBe+gqBwzhoh/tpC+zyWugL95PqCWIEooR2uouBJ8WsPebjITHm4Usx5pcxgcFhRYgK5sHokpzpv8+k9YKEoc0fxNaLmbRgvjqOtsB28Fg4QV69Vu3jfp468fvg7/SzInAsIpCRnpGOJkV+xkZqo317dpsUedk+KoFKe8IjIiNtUrxS8tPGsXIvEc+MZfni+Rw60KIIKAKKgCJQShBQwqKUTIR2QxFQBBQBRaB8IFApoXKVsy645MoN/6xZRb7c8jFqHaUiUOYQwIGPU/oEsWvEECSm4AzGgYxTGocpmgM4Ocj5v06MyAMc1zi7sy1+HQt324pWWr+69lbHR/oEvHMsaR4rddxO7/gwuxU9dY9lX5ro3SspnyBK5glZwSl8iIb1Hq/VSO6ZKQOwJ7p9zn/+vY8jnvdECRA1gCOeKAJO85NmyaSLwiFPRAIkA2PFCQ4OXIesIGoAMyrSkBM4u/lMVAEEAQ502jPi3tRFhAr9wyFGvURCkFaKz+CJ8xxM+YzmBc+AoUmRJW995BHfQ7JAKBgyZLn/GsSKSd1kIgl4ZS55JWoAcgkigagZcKnnf8akU+JesOBeQ6QwNvoCLuDAmCm0b4gcnjvZ3w7X6SNjtBBZZ779z+TlhbYgUsAZPCEQWFcdxVhbPcSI7DBrESINzEaIQZqtE5IhK0JCyAr6C+l2mr9/Zj7BhD6inUEaKJybWQ7L0kZUGOCat2pLNIi1avnSRXkBU+9RBMo6AokH9+8nbZHwClG5aSygScF41635m/8m5VpSkpOTSA1VXskKAGoqmnIZGenpq1cs4793WhQBRUARUARKCQJKWJSSidBuKAKKgCKgCJQPBC6/7pY7wsIjIr776rOPy8eIdZSKQJlDACcxDmhOsnNiHQ0BU0y6DSIXcFZ/Joaj3qQLShZH72En1HMYvWdAA3tMnNO6Prt7NqZa20Zt965PEb0KISGmSFTFgs2pVkeJouDkPY5tnPikJBothlN6g3ictyW7LXkkS4uBaAPSNxH9YYSsuZfrcwLq4Tuc85zkJ10Q73FoMzZO5+PkBxsc/vwNgSOcZ3Dwm5P9EA0QDyZKg3s5wY9zHbzq+fuyXl4hAOg/pAQkCk52sCMVFfWTgopXCADGSJ3UAZFACiefJoXd5htbBUmttddls8JFv8O7N9NXT0ys00oTomddkts3DvpA35hDE1HBWMGR9iEBmHMTjUG9OLCIAjFC44zvKzHIkS5iFOrm9DP9N7oeYEY9BTmxbEgdSAvqg2QBQ4gZCDTWHiUwLRlr1ESSRAlJQT+ZH4gicOwnZrQ1GBfYgTOkEfjj5Cz1ZAWDbta6nY+wWLl0Ef3Xoggc8wjs3b2bvW3FxsXHp6ZszjFdW2Zmho8sX7FkIURkrgUSBNIi1xuP4RsgQdesXLGU1FvH8DB1aIqAIqAIlDkElLAoc1OmHVYEFAFFQBEoqwgkVKlW/Zpb7rxf0grv+3bkpx+W1XFovxWBYxgBnMA4eXHOI65MKijjIA4cNo5kTqQTnYBzGse8Jw9poLLq4NS9Z+2BPRId8b6kb2olIto7d6RbeyUpx+7f9nsPLkm0nJtSvZu3pltOiaRYJfetllf6hEMK8oEoBpzsOOHpBxETONK9uzJ8DnQIB07m4+xmPJyoxym9WsxECfAsfw/gwKZAPvAeUgAsiFiAJMApT5QAz5koC65xH6QDbZnUU0bfAcca12ifdkjDZAS6iUCgLogDolQYB6SBEb2GIOFeSAra4ToEC5ofiYLXBiEnUutEWM0FtxrHR9qqN4u2qoqex36JVqm8IsnasTbFm9S2oi1TOpMoabP+Oej24Qb5ABZGg0Pe+saL476Rvx84+5lP5pi2iYSDfGglxlo4VcykimIOqIt6ec5EXXCNAua5FqIZQuioGE0PE91C+6TzMqRIYL30i7VKvzGc+j3F0KiY5++XifoYK59nixGtkZ6fNZvrQErghhZt2ndyZ2Zmrlm5nH2nRRE45hHYu2eXj7CIrlCR38kci10E0rhh5dLFeSL0oqIrVMiL1kVu7ZbV7zlAVL9R0+Zj9RBRWZ1C7bcioAgcwwgoYXEMT64OTRFQBBQBRaD0IOB0ulwD3/rwi5jYuEqvPfe/B4WzwOmkRRFQBEoHAjiWcaDjfMf5TFqji8RItWOc+6anw+QNDl9OvOPMRlzbl4Yjv6VqmLVv0m7v2KphtpXzDng961OtsBS3tVEiKZpLiMSFUh9OfJOaiCgD0jrhFOf0LJ+NDgUEBffiNMdhBbHBCX1IA07W46THAY7Tmu8hPIiiMKfq+Q5SAOLB5D2nXeOYx9kPcQGBgAOd8fIdjnyuQ2zwrNGRMMLkECDgCZlCH+gfz9E/sKY++sN9/CZCUtBv2sPxnh5htxxC1HgTXJY9zmXVPb+yraXLbjUVUmLTeZVtdbekee37MqxqTaJtTSs4vPPk3nUVRMB8dbK1VKIrRB5EOmcXbNy+8YIZjnpSYdE+4zZ9JoUKfeGULddwDjYXIyKBdF+sCaIV2olBcGAQBaRqAgOeI1rBR16JgVFGXtNBZZOCiflxC5lBnaRAor+QU13FbhIzhTVKlMXNYuBI/0kTBuZE0YwSIyrnO7HZ0hbzViZLMzkNvVoEt/NzGrpD15NOSUlOSlq+eIHmqC+Ts16wTtepV79hx27de6xcunD+iiWL8hRxULCWivepvbv9hEXF3AmL9l1OQO/G8khuqLz0qlqNmrW3bPqX35Ss4nA6nWitSZTGvG1bNvFbecyWpi1bt2O8yxap4PYxO8k6MEVAESizCChhUWanTjuuCCgCioAicLQRuOOhx5/tdOIppz3X756+69eswgEYssgBtoovvPXxiM4n9Tj9z19mTB358ZA3j3bftX1FQBE4DAEc7Jhx5PaS93f778ARvV4Mh/5CMXQCZonhfDdO/XzBKboGvvu7zRXFCV8dXqPDgMMcUoI2/xYj0oDIAkgKI0qNBgGn7Y24M3UYfQkc2zjXjSYFRAGkCmPDkQ1BQL9xZtF3kyaJ73B6Q0YYPQf6wnujo2A0FcCI/lCXIVOMroR5hs/ck+GyMsIdlnundGC927JHpVthfMffIBAsjJVnGAugeCV6Ik5IhmghGSJ6V7clnRhnq7kr3dsk3mVL2JDqXVc/0tYwymHFNImy6ko6KHftcJutWpgVJkTFFiE3FottkmiUapIOauPs/d4D4XYrUVJkQVJAOCAsDlkCkcPYSS0F8cAJZsgpiAec/CYtEyQG+CGmDSkEYcCzRFAgSg5JAG7gDGkDHjzL+CBd8poeTG7NsTAP1G0iQ4wGSVu5xnzWEyNFFcZnSBaiPxgP/UcUfCLPC1mRHz2N3PpVot+jAVW9Zu06v82Y8mNeG77oqutvfvrVdz5CgPjUNsdDUmkpJwgQ0XrF9X3vRFB66cJ5cx67s89Vmzdu4PexTJWd27fyOyUpoSrxO5Nj6XryaWdygyssLDBlXLbP1Kh1XN0/f5s5LfCGZ18b8sl5l1x57dQfvhv9yO3XX55bm2X5e6OJs0zWR1keh/ZdEVAEFIFjEQElLI7FWdUxKQKKgCKgCJQIAuuEpLjlnkf6fz3pt4WQEOO+/nzY+rWrcTL6StXqNWuddnavi2+868HHeL9k/tzZ/PHnkVIiHdRGFAFFIFcE5PQ6znyIAZyZ7cU4iX9JwIM4fki19I3YVDFOo+LgxoGMczjfOgVy6j6wXx4hMCABIAToB05uHFQ48XGS8x5nPiQEDisc/Tii+a3hXhzmOLLpD+9xnFMPhXuNQDbfUw9EAs9x3ZARgSLV5veJ/nCfcbozTpNWilcTfcF7kw7J1E3fM6JtSckRVqqzvn1d4t+eJs5IK9PrtPbv2++N8aU2SbPCE89z/dhgqbuFa4PnuDghKyxJ41TpmupW3QSXrZmkdzpZLtmi7LYVQkAcn+qxrZNOLBPdj6ZyPUWiUZLCHNZfezOsLUJORPyTYq3eleHdszXNihadjwxJG1VLyAr6SR/pE6esISZIU2UianDmgyvfQ0KwDoyeBjhyP0QHBAdOLXChPp5BrJrCPcwPdVJ3UREVvspJ2+TXpYB4gShC12KmGOQPDkpwN4X5p3849SeJTRfbW5aJCjOwZi3bsD+t/JyGjq9chT1krVub/aGCAOz07TGEwEtPPHz3kEEvPHXORZf3vu/xAS+//+X4KZef0bV1bsLVpQ0CE+UQn3BoLWdXiBToIgdj+N4uJbdxSIap2Bq169TdtGEdv4FZpTztmRZtOnRiPaxdvZJDA1oUAUVAEVAEShECSliUosnQrigCioAioAiULQR+Gjf6S/7Qe/Cpga/1ueP+flh6WmrqQRGpiIqqUCEyKsrnNOSPoWHvvPbi0NdfejY/aSzKFhraW0WgzCIAIYEANClzICo6i5FGiUJ0AyfUEVomDRT3krLogHEAh9AeKAgQONU5kQ+JgPOfdnBOk56Jk/I4n0jNwX1obEBEmKgI/j2Psx3SA2e10Y3AwW6c6zyPmVRF3GMiAAwRYe6l/1wzZkiK4HGZlCPme+6nDV8qpNr2zc6K1sHkKvadzkrWPlekPdX5UsTjjfd54/at9jSyWjqW1Uqw7Q2LspJazXO3m5dmi3YMdQ3dcmstW5OGUb50R3GiV9FAIidWRzisLRIp0bF+pNVSyIlZuzOsxcsSvYvnHbTs61O820VkO/1AphW2/5DYthmbN9rhwwx8/JEsWZEcRlidvoI5Rnon7lvvx5Hfb4gVnITkg4ckoH5euRcSiwgRCCUwgERivUAeMYeZeU0HFQxsqM8BpIUZD+sVEorT0aSpgkAxTkoTGcMaof9EzpTZNFAGjyYt2zBOa+mCv/7MC2bc88m7g1/6efLE8f+uW4t2i5ZyhoBk39zz1acfvJOWlpb61Ctvf9jrst7Xj/784/fLEgz8G5IIoSrVa5DSLtvStmPXEyEhuIGoktzG2KRFayK0rOWL5h+WKu2hvr0vqVajVu3AAzi51VVWv0cTZ4WkDJMMWnlKoVVWx6n9VgQUAUWgLCKghEVZnDXtsyKgCCgCikCpQYA0Azddclb3Zq3atD/p1LPObdC0WcuKMXFxqSnJyTu2bd28dOFfc2ZN+fF7hLZLTae1I4qAIuBDQMgG/i3MiXq0CdAFQLjYCFMjwoyjeowYjl/u40T9nmI6rW4iG3As4xjH+UyKJ6MvQb8gMYywsiE2AskHSArjqDJERCChYIkTPTAixPdeIjwCr9lC3ZPDkvHK86bvtJX5RPhLVjP7Ss90dw97N8efmVc4R3fz45vgtWxp3exzwp1W5nHS02SP136wp3NG/W3OFgvfqjH7xozobudJJYhLM27hK6zVkXZrpURMbJEPU+Yf9K6bsMubLqLkJrrEpLACt8BxeJLcWZoedN9En/Ac9xKdwJyCmYlggaiCpABbnPyQEczDP2JE1RBpYSIweMbUBeFBVAYaFpAI4FxkkXSyTiGwiKwgrdUVYk38Y2jjHxekGkQWItukvKknRtSHOTmdKHVslXVbpJEfjLMkS9MWrduJFEXi2lUrGG+eildKfu7PU6V6U5lD4IcxX33+0FMvDu4mKZPKGmEB2Fsll1XV6jUgSrMtJ556xjms97yQFVTSvsuJJ/MarO0i/3xNKg9kBela6zZo1OTXj997o8wtaO2wIqAIKALlAAElLMrBJOsQFQFFQBFQBIofLWBESwAAIABJREFUAQQdy7KoY/EjpC0oAqUHAX8aKKIRSP+EMx2iwjiDcLpDVlAQVCb3Pw5s9Ax2itOXyIQiLQEponxplvwEAI5y2sURTl+NyLXRzTA6C8Zhb/oUTEh4glJQHdH3oO8Lk+LKF5XRf6qPNLFd4vqOvuFEbyPEBKRQmN3miffY7GHiVou22bxum+XdG2mlVK8SHuf+N6Jpdz9ZAfMwRhQ+ZsozM/dlWuslesJ9VZOYDMEmMNUJp2JNJIgZl4+wMaRLAJnCvUZ3xOhxMJcYBAZOcKInOKFM5AT3GkPXAmLDCI4bcoJXnmdOfPUUlKgIEalDFAjrE82SE8QeEWONQpRAnDEGIkgQ4yZN2WN+ALjflB7yhrXM33yzpA2It3SiNQLuKTNvm0qExfLF8//Ka1pFlyTybyqHCUjHmN0ga9Wpe3x8larVNkg6RzlXAD5aSgCBuPiEyscd36DRjm1bNm/bvIl9V+hCfdlF0hDdul7SgjHfhW5IKiCCVgJqU/K6FgvbphAW/1aT/E051XPKGeecj1B289btOuaFtOh84smnbVz/zxqiUEy9pIOKEa2M7HTZSnrchcENDOwOh8OdmRmSqCUdFKmzli0omH4FmjpJElJd3JHTTqfLlZmZUeT/7igMtvqsIqAIKAIlgUCuuQ1LohPahiKgCCgCioAioAgoAoqAIlASCPjJCk7X1xPjxDwRC5yqD3QGrZfP88QgK3j9XmxNKLJCrhVHt3H0G/0IQ1TgPPeljhKnOOYW86UdwjmfgxVH/3Ks09bTRyIYXQxO/tcWoqKCmC9Vkt3yRDts7ih59chrhFhmRObapnZvOpEMviIPLxdNi98kLdTe6mFWhohsu5k7PyHAeBm3GTsEhTEfFqYeg4sfOzA1qbJ4j4MaEgJnEGm1SLXF3ENOQQqgE0KUAtEVpHuaK7bYf41oF64TVUE6KMgLyCbTdJ5f/WQFeEFSkIoKpypk2UCx8WIviEFW0B9yrZPe6E2x6/z34JD/QYy1uj6gYdY0C5Q1zlqvJxbh3wN57l9puDEqOrpCnXr1GxLVSH9wyr4yZPioD0f9MOP8y3vfEKqPV/W59e7Pxk37w6S+CbwHMmPQB1+MmfD7kn+4Z+qCNdtuvf+xp4pirGddcNlV1PnRNxNnDhk5bvK7X4z96Z3Pxkx885NR378x7Ktxgz8aOZa2H33u1bcC26ssR+jf+vSbCSadZKi+4LwMC4/g96vQpTDtdT7xlNOeeOnNoaLtnCXuDAnBmAa8PnQ45EF2HUTXa+q81VuHfzf19x9nL98AFhGRkVGFGRD9GTdrwSpIrezqgZCSaYf8PaKg/3DZdTffPvTL8VNHT/tz6cC3Px5RpVr2KZhGTZm9+O5Hn2Z/+kqPM8+7kLkeOXHWX2ibFWYsoZ7dumnjBsnSZFIVHnFL7ePq1a/fqGnzGT9N+I4vHTKgnPoQIwrebTt1PfH3n6eic5NVnnrlnY8+GTPpF/AI9XxJjLswa4s+I05O+q9fV2w58PvfWxOzmw/SQXH/kgVzs1LMNWrWsnW/Z19589EBg95u0LgZZHvIwj78ZursJdf0vesBcwPkx5U33HrXmOlzls1atnEvfeA+8z3jGvrV99PoV/+Brw/JaX4gWtgnk//6e/Ofa3em8pvBb1bwM7R3450PPBp4nTG8+M6wkUQU5fRbUtRrVOtTBBQBRaCoEdAIi6JGVOtTBBQBRUARUAQUAUVAESjtCOAUxvmPs/pSsdPEAk9hrpHPr4jhQMZRnVSS6XSCRblLO5jB/fNO9aVR4u8MHKu85wSv0XxAnBonuskZzjxEhmWs3xOT9NOi3bE3kPKI8qxYD7H1YjvExoqtFWf7IT2GjQeMJgei1LlCFEhi+EkF2g/W4TCEBgQEhc8QCUaEm/c4aM2zvgiP3CJYTOdCRFEYnIikgFxAS+Uc/7iJmuB6df/zv/lxQEz7dzHIHXPqFpy/Fhsp1k+snv8ZyCLW9kKxz8TAmrVf5vQsGjdv1YYT0xAWPc+76LIX3/l4JLn9XeLF69itew9y/P8ybRKkTVbZsX0bKb0snLl/L1sMBlkFMuP0cy64ZPpP349ds3LZksuuvfn2Ox56/NnZv0yfsnjenD8C783ve7cc6cbhKHICcZxeP7h/3y4cwFGSg0YO5leoWqNm7eo1a9eZ8+tM9EeyyvmXXX09aXrS5ch2qDajRaBg+Lipv/82Y8qPrz//BBE3hSqFaQ9natfup57xzecfDwFbnMQ4uus1bIy2itW8TbuOl57W+QiHL+kz7xFH/8qlixfMmDThu9PO7nUx80BaIrS+CjogE+lQS+Z65dJFpPI7ogjnVZF1EvwFRMvbw0f/0LJth87okiFyfWavi6+AdLnu/FO7kGYp8BnGypoy1+597JkXwWPPrp07cFr3ufP+fp8OeeOVojwVv3Xzvxuq16qTLWFx6lm9LqI/U38cN+aufk8+z/rLCUvux5n++8ypPwXet3P71i3gIdmSYgIjL7inpMZd0LVFH6tWr1kLohAy7vvRI4Y3a9m2/R0P93/uh7FffQHpEzjWFjLfzNmWTf+u5zrO/0eeeekNsOO35pwLL7v6gu5tG4WKvKpZ57h6CZWrVsuQyB2eZd4Hym/SWedfeiVRK4kHDuy/+Oobbvl72ZKF33z+0RDIg6tvuv3eP36eNolIH8ixH8Z+/cXCubP5XT+sMC+DPvh89Mk9zzl/yoSx33gtr5d6z7zgkitJbWZu5r77+w/wrbNP3nv9Za6zhod+NWEaBC+fw8LDwl/s/9BdBd1X+pwioAgoAkcTASUsjib62rYioAgoAoqAIqAIKAKKQEkjgNMZIWJ0ADix2NzfgcB/FyOc/KtYnJhJwVTS/Swz7QlBEVgCxV6Ns5/vIR3AEyc6mg+EIqDLAAGx0+bN3B13YMz43bHXSySB7Wl/hafKKyeAmZtbxYjQwOkEoYDTHcfydiECcBoxTyFTfwQTGkEaHWh40JwhJwLHgqPSl6Yr4KKJdAlORZXtfAURFSaSAodSezEICtJlcdqXdWkKOh4mVQ5RHhAOk8UQfc80aZ2kbqN1QmooBtI7oA6zplnjOJLpO1EaEEhlKi1Uo6YtWzOu5MSDB4lS+HX65ImP33PzNZwq/2LCzDlX33THvcGERWZGOuO11q5eSVTKYYWojA3/rFn18K3XXopD+sdxo7985JmX39i1fRsEZaHK1B++G42FqoToiOHfTYFwsvrdkUXO+W7tfFKP0//8dcbU7FLY3Pu/Z17k1HdhHPuBfSpoezhzcYyizbXm7+VLqfOZ194bVlVCAJ64r+91515y1bUnnHL6WUTE4LwNbPP8y665gefvu/GK83GOf/Hh24OfGfTeMEijwoC+6d91vugs8VdnmzYpoWq16iuXLJwf2A5E0lsS+dKsZZv2Ax9/8M7RX3z8PuvhulvveejBJ18Y1KxV2w7BGg9G+2Hubz9Pv67v3Q/iYMeR/MLj99+BuDfO/qIkK+gvznaiIiCtkhIP8vt5WOlxdq+LVq9YupjUZnzhzCXCAtIvXXJazf191ozAisT3nb57147twWQF95TEuAuztnDgv/bhiG/jhUi46dKzukNcNWraotWoKX8shrgIJixat+/UdcmCv3zRFRdcfk2fx54f9M5P8jvw8lOP3HvuxVdcw+8B0VIQDsF4N2zSvCXXIDx4ve2Bx56GVEDg/dWn+93XVbRS3v382x87SdqtNh27nMB+uOvai8/+Y9b0yd1PP+s8IqkgPEKteUiIU84494Ln+t3Td+yXwz8Ck64nndqzRev2HQMJi4ZNm7ckMmnW1J8nUA9r49Whn4/esXXzpjcGPtnvfy8Mfo/IHyUsCvPLos8qAorA0URACYujib62rQgoAoqAIqAIKAKKgCJQYggEpIOqK422FcPpHSqHz7dyndPrpPvJs2O6xAZSyhqSFFCBxesnMIxmBGmK2skZ5SjRrQDvbW6Pfb+g6rHbvW673RNps/lSHP1bMXnmLqd772uZjniICp8grJSzxIgcIFIglOgsJ0shniAcPqJ+MQgM5i9PwtcBBEZIJ36QKLmJysiPwx9SgcgG1l0NMdJPNRDjlDzC2aHKerk4GFzEiA7YJCSFaTvwfvoB6eNLSSXG2u0TVCFrnBPhRGIwB+tlL6SUJS2LBk2atti9c/u2vvc/+iSnlvvdfsMV4ltNx5lMpEVNOfIeDCLOZpy7xokb+H3NOvWOX7bwrznm9Dw5+3EoZjMXRXb58YGD32ssKVtuufzcHoFOYRznbTt2PXHo6y8SWXREYXyX9O7Tl9PeUyeOH1PYDhWmPaIYxDca+8O3X38BuXL6uRdeimP04duuu2zaxHFjOKGOg5aUSsGERU3RkOAZyArGgMDzo3f2ubKw49mxdcsmSIJqErkSqi6cuWD443ej+C3JKnc+1P+5VuK4fvrBO24c/82IT80Xf/3xy0zeH9JNWfBX4DNduvfoibM/UdbWfY8/9zIi3i88/sAd5p7i0EJBw4L6Bb96EBOB/SGa4NDaeelZ1jN9E14MMjhkwVHe9eRTz5j+4/djwT/wJvbMsoXzSX13RCmJcRdmbV1/+70PQ6RBBJooG5NqjKinwAFVl/RarM8lCz58F/Kh/0tvvA9ZAQkKhov++tNHKopsCL/ZR5QGfsKC6AxSMN1898OPz5z8w7hXhOzgeYn88qWCOrnn2b2Sk5IS+8p+X+0n5apLeAbf7ZLfs+CKITd633zHfaM++/A9yAq+pz7GkRk0BlmbEN4WkUq8SoqyF2RbxtKWdOuf0yRyqdclV10H4REcJZTd2tDrioAioAiUJgSUsChNs6F9UQQUAUVAEVAEFAFFQBEoTgQ43U6udJzHOBRwMq0MavAe+Yw2ASk1fCe0y5JjtzjBy2fdYO1dt6GKY8XqGjNTUly7a1Tbn5GSGlZp2/bYK0RGND4yImN/q+abfqhebf9mp8Pzu9Pp9rZcUy9xYZMDveTZj8Uu97dJ1ACn5EMRFqT0It0UxaTJ+VDeEyGDDsU6cc6bNEg47nHYe/MzpwEpn0KSFCFSPfE3FuuMaJJ4MUS8XxVrlQOGnNQdJ8bpaaJIOPkLUWGExT3B7RA5wjjkunHGQdywdlnDbwe0BW6ni+EAAwv65sMhh/6Uqq+Ob9ikGWLATVu0aXfZ6Z1bQlbQQRxxSaJ8K75jdDoOKziily74j5QI/PKApGrKKcVOcQz+oquuv/nCK6698d1XBjyxYO4frM+sIiRGG5ySK5YuOiwCwNzQ975+T3CCfMLoLz/DIV3Y/hWmPaMT8ev0SRPJq//QkwNfmzR+9FeQFfQrMG9/cD/BHbIEZ7EhLQo7Fp4nJZTod2+sXiN0hEWrdh274LhdMOc/3InO6SP5/yd//+2oQLKC+pKF6eKVNEjB/evQ9aRTFopDG60DTui/9NQj7LdiLZKm6hBhIaRLMGHR87wLLyMl0U/jvvmSe5KESRGChtR7IctFV19/M3M0UVISBd7ANVJ2ffjmq8+HerAkxl3QtcU83XTXQ/8jXRpplEz/m/g1TVavODyCp1W7Tl24Z9nCeXOfe/39TzdvWP/Ps4/cdYtx7Butk1C/KzwnP0ctuXfV8iWL3hj29XhIqmcevutm83zd+o2I4PTtBUgQQ1ZwrX7jpr6ozk3SZjDO9z8+4JW9u3ftfHPgU1m6FKRZC5cfh+B5l6Azn14LY2YtX3H9LXe+2P/BOyErTNuWrPliXZhauSKgCCgCxYiAEhbFCK5WrQgoAoqAIqAIKAKKgCJQOhDwR1dAQkBUIGrcVwyHcpWAHpJPmhQmJg1UmXHolg6UD+uF9+811cOXrajVOjkl7PyMTMd5Bw5GZkqUhS+vfVq600pMirBm/Nr0OLvN+12luOQ5F5yzABHsDHHCH5T5ulHeI4J9t79WnDzDxMjhTfTEY2IQG+g+mMJ15pe5xSjMJ+lmcNiT/oQ8+S6pn7RIOPdxSBrh7MCIDBw91GcibIiSMGLi1Mv35m8pvoMs4HsiQxDMhkSBKGCthTylK9dJ9QSB8InYKDFICxzvPnFyf3150egw65T+s3YZM2v5RDoqpbv/FUzQZuE7h2CQL+LGX8dReRH/XzOc40NeG/i0yTlvOhIq3z6n/Fu27dh5xEfvvB6qw6RegkBAp+DfdWuJ8CnWggbH/yTlzOxfZkwZ9u6RWg1tOnTuRgeCnZJcI7XS+ZcdEhYPjhAoaKcL016TFq2ITrPm/v7LDPL0o3nw2nP9HzJ9MeLQ+/fuYV8dVsCddFykxfl25KcQi0VWtmzcsB5tkFAVih5AL0gNc3Kee/rccX8/j8ftJn1O8DNGA0AyPB1GDnGdtFxEmCRUqVrtijO6tc4uhVeRDUwqQntDpE3SQp34P/eiK3qvWLJwnlnHRBVFyaYI1T7ExqW9b7yV+n6bcbh+BQ5wUpYtnn+khktJjbuga+vSa2+6TSRiKr436PmnzLhx8l8vqb3m//nbrODfDMhM1kOTFq3bNmnequ31F57ejUgt8yyRHrzP7rehQZNmLfiuVfvOXTudcPKpROgErnfIHZ4nUiJYJ6TTCd1PhVQgYixwjlrLbwBC6OjTEJVhvut7b78nmNOZk36A0M4qTZq3brteUoBB/KG9QeRZ4J4iigSCUKMrinInal2KgCJQkgjwj2stioAioAgoAoqAIqAIKAKKwLGOAM5lnNk4j3GGQ1YEF07x4/DlhGJIPYRjHaSiGJ+kiPIuWFzXvXZ9VdeBxMhbhKwQnQBbEz9ZcViaJrlWX1JEPbhnX/SLv85ulKWeLaQFqUqeExse0Keb5P0tYjj2rxHjhClpMc4QIy3GrBD9hzg4V4y6LxRD6PgXsWVinAj/WWyKGHVjV4kRtfGE2G3+91xHuBRh24fFSEOF8x/yBDFwHK+cjN8o9r0YGhz0r4cY6w3iA/LFl+9cCo5cHOmQKB3EBoiR5sUn8O6/vyBkGWuWtcsaPkK3Qa6x5ln79Im9UCYOr+EcJu0NKZS++uT9wMgRi6gEHJOb/RoGfnzlBHTzljhZOQlvrgW+jv3qMyJ4rMvE0Rnq+6K8RjqiQZJbnv73v/eWa41AdGAbzSU/PfnwTU78wO/ueKj/s0QlcPJ62aLQ6Xry29/CtIejFAfwPunQjXc98NhnQ98cFBgtwelynKQbRcA6uF/Tfhz/LdoXxYE7UQjVQmhYEFlByqq/RK/B6D8gznzOxZf3njT+26+DtQ3oM9/zGky6NBRNBOqDGME5jMM4v9gX5H7wFP/2FlJCBT5fu+7xDXC+/zj2v1RXwhPtQu8iVDsQRZAepBsK1tnAYS78jXuppEoLfrakxl3QtYUGxZL5c2eb9F38LrDnEqpUq/7SEw8b0jtrWK3aduyyWUiD6269+8FRIhwfvK9I28bNRFAEY0HURN36DRsvnjfnj1vuebg/ovMTxnyJxpCv0HaXk045neiM9159/snA51lXEF6QKMH1Mgaip0wqKL6/7YH/PY2exqtPP3o/+8Y8wxqEBIVcIgIDTZLBAx5/KPC3pZ7sw+CUbAVZe/qMIqAIKAJHC4Ey8Y/UowWOtqsIKAKKgCKgCCgCioAiUPYR8AsTc+IUJxROa5NCyAyO1Dvk958thgOKk5YFcRiXfbCKYAQf39jdtmSFp4rbbX9PtCsuCagyRXQrRjocnpWSAiouM9NeWcgMvifKxb5hY+W2J3VdDaHgK0Ja7JS5u0/e4qjhlQIRgPH5BzGc/KR+ImogVoxIDCIcOBmNc57T4OEBfSCiwRQTeYD46bsB17N7GxhhkYfbfbdAICAczrri1Cy5+yETiO6AWCDKIa915XYf/WPt0hZrmfGBg+9EvL+w9tkDECObBd990n6etD5ya7y4vq/X4FB6lcnfj/k6OOe+OMcRJ7dWrVh2WF5/nK84eXEqhuoX1+fP+f2XS+S0+UdvvfpCcegOmHafFUHqWqLd0PfKXqeFIiS4jxPbRsA6sL84I8+64FJINAvnZFGdli5Me5yCJ1LhzF4XXyG+2ajPP3j7tcA+UzeERqjUVZxi/+rToe9warxL91N7/vnLjKlFtW62ic4DxBaROCZlGHV3OalHT5z07776HCSkr4ApjudQgsp8j4Oe13+CBNsRceY6URWfvvcGxGWJlR2S86qG5IQKbPCCK67pQ18mfvdNljbHHhHNxlEfqmM3SFQJ9389/MMjfu/YM6tEHyPwdL+po6TGXZC1xdxCIBhiovOJp5zW/8U33pesY7Xvv+mqCwPTMTEeyD9SX7FO2PfvvTrgMFKBe9Cl4LdmUwjSjZROrJ00Wcwdu3XvgYB8IFFw6lm9LoJE/fKToW8H/66cfu4FkOHWrCk/QmwfVrqdcvqZs6b+NAFigqiqxwYMevuEHj3PhvQYN+oLovCyCkQVhCx6Iwi/E7lldFe4KbZSfEJ85SpVf5k+if9GalEEFAFFoEwioBEWZXLatNOKgCKgCCgCioAioAgoAsEIkOM/hJG6B4c1DpzOYmeK+QQxAwrOTgSOl4rhyC3VDtwyMPPhQka8YMgKkfycJiTFB9FRaQ9Vq7J/aJOGW8ddfuHcty46b/6jNarvO8nldL8qaaH+FvKi8bAR3UnblVXEmU6KJFK2nB807jfl8yCxy8QaiZGSaZfcP11ecaC+L4ZQN6k9yFeOsO+9YkRFFDR6Jqd84Cuk3sDT1qSfgow5SQwhZRxORIv8JH3cIJaM/kQRkhUGHtYua5i1zJo+zJEvn1n77AH2AnsinHRpofZOEN5H7SNOexr/89efs8gs0xlEgnkffBK6dbtOXdcKi5FdDnqeeV/SS5FG5sobbiV6pljK1Tfdfi+i1O+88lz/UKeqaZTT0mh0bPjnyNP6t9736JOS6mgd9y2WE+RF0cnCtIdWAKfE/16+ZOF1t97z4KdD3ngFzQTTL5zBpNkKdTLd3PP50LdfI9LhpjsfIK1bkRXJjLOJlEekwgms9NJrbryVPhLdYa6fdNqZ5xIVkh2h1bX7qWdAuKxZuYJ9lFWI3OEDAssS0UFEVYkVyK5qkm8rEOuLrrzupplTJo4PTC+0c9vWLVWEuAnuWPsuJ57crlO3k8Bh+9bNm4K/b92uc1eJSIL4PaKUxLgLurYYFx1OEabl4zE/zRr61ffTIBOuOa9HJxz5wYORAIfWEAqkjSPFXGDkgrmXe9aISHaoaKjWEtHCfc3btO9IZAYkQ2Ab519+jS99W2CkhPn+jF4XX866+v3nqZDYWYWIHfRJNvyzZtWA14cO/27mvJXNW7fr+OAtvS/+8K1XjtAUMREgzGOvS6+6bkhAKiwqJYqD15z2YYktXG1IEVAEFIECIqARFgUETh9TBBQBRUARUAQUAUVAESgTCOBkJnqC6Io2YqQQCi6kZyDKgpQ9hRa0LROoFG8n46R630lSf1kaFZk+LCE+cf+OnTEt9uytUE3Ii1lxsSnuvXuja2e67Y1EGnSl12Pjb5MaEqGB051IgX03f/ILUQNoOnBSlDz/14tBRHDqnqgZBKTT/PcgQM18I1TtFjKA59DFQHh7rrxyWAuHPYKmvqgOMerHCUifqStSrKoYJBen83FQ9hCDSKFuTvRzKhwihXQhODTRwSBqgvXDGtsshkYGawlNjmKN1oH0CBLkpl0iT8ABLMEssLAH6CdCvtwHfsXax6D28/URBzgPrFv9N6TQYYX88eT2J3974BdtOnY5Yc5vP0NeZVvmSoog0shceeOtd3/y3usvB6fIyVcnQ9yM0PODT74w6Jdpk37AsZ9dffEihiCBCtHB+fIhMYgEGP7+m6/eKOLQ9LWwfeL5wrRHGhrqIM0VDtavh39w2En94yQchpPrOTlKcRCPGv7hezfe9eBjnGQPpdtRkHEaAoG0SSYVjnSx/mlnn38xp92NRgGkBvomP4ujP1TECmNj/aA9EBipQZ8aNm3ui7AIFukuSH/z+wzpqVq27QDR6Cunn3PBJYiXfzvikw8C6yK6RQIsagZHmtx8z8OPc9+nQ14/IjKEyBQiFRbOnR2asCiBcRd0bbXt2NWn1fPs4CGfoA2BnsSEb7/6nPRWoTBu2faQ4DZrZMzIw7HjeqWEylWIUJkRpBlh6mrd/pDejAiEt3/wlqtJE5hVIB6I6CFNVPB+huijr6y74EixNv4xMEeQrB+/M2jg8PffGmRSmAWPo3Hzlr59iObFX7N/+xnx98B7/iMslh6R0iq/607vVwQUAUXgaCGghMXRQl7bVQQUAUVAEVAEFAFFQBEoCQRwNHPaFCfFddk0iCgzApikHkJvQEsBERCygSdxfgcQP7YVGRmOxG3bY48TciJWUkW1nDOvQUO5iXkh3c1xEo0xXSIx3rK8tpryGbJgg9gBMeN0ok6cMvPEENtGe2Cif95oi+/52waS4ojiJw18RIYYTnoMRz8kBFEIJnqCV0NOcAupOxDqNkQIkRwmQgPCw4hjG3Hu34ohaiLUkLK7Rj9YwxAmkBWs7VCFvQDBArlCqqpSG1VUs/ahvP27dmzzzZkpnJA+4ZTTzyI9ESeqzXVEoCE5PnjzZbRBciyff/jO4FeGDB9Fbv8Zkyagg1IkhdPirwz5bNSu7du3Pnn/rdfnlMqpao0aPr0EOSwNgZRV7ur35PNLxRFJih9Oei9bNA/SrdClMO0Zh/1Jp55xzoiPh7wZ7HglHRQdXLFkEZou2ZaRw95/64bb73uECIFXn3n0/kIPSirYvmWzL+KB9FumvttF/wMiKpAwqiqpgkins3LpogWh2u116dXX4eyf8sN3o4O/x6kO4fL7zGmHnZAviv7nVgeERWVxpBMhw3q6/rZ7HyZl0R+zpk8OfJZT+kS6kCbJpBkjEom9whoPNTcQNNSxSLzfofpREuMu6Noi6gQR8ecfu+82xhcqKiJwTC3bHSJ9iFwIJZhuiBNZHyHXMJohPE+6sCOiKy7rfQOE2LSJ49FHOqyc0es+zRe+AAAgAElEQVSiy5m7qRPHHfEd6au4efCA/g+PGTFsaKi0XIGVkbKMMRNd8egdfYgePKw0aNK0BWskuzWe21rT7xUBRUARKA0IKGFRGmZB+6AIKAKKgCKgCCgCioAiUCgEgk6Ym7pwKHMKH7FhnBScog8uOCVw1uJ4PsLZfZSdz4XC5Cg+TBRDVg51ISPeT01zrZZrzEeDEP0ihVGyCHCDP3OEEz1Uai7jjB8v3xPlYKIvAkmDfA07IPohMMIg5Mlcf8VZjvF8NVTyN4MluLC2WePBkUXgzJ4gusiQdYeRFuyp0rD+JR17ZU5LB+eD737aWedBTkwPSPUDzCZly6JsTosHTsVMOUXNieaTe57dq6gIC5ySA9744DNOud902dknI7Zt2iS3PI7jHwM0B+IrV0VDxQpM64OeACfob+994Rm9LrnqOr7LzYmZ1yVWmPaMlkHtuvUbfC1aFMFtmpPd2Tl7zf2QT6TrAfeiIixMhAWRArSDTsE5F13eW6I53g0ku0y6pGACzPTt0mv63Ao5MGXCd98Ejo+IEsSsJ44dNaKoo3HyMneIaUNExAgZ1qBR0+Yt2rTvNPDxB+8MJsOM7kYDSV9lCIt7HntmIPe9P/jFZ0K11UbWG/iFSnNVUuMu6NoSOBKIrAhM+ZUTnghus+cnjRvzVaj7Gjdt4RPcXrFk4RGEBUQkRBDff/HBO4ODsT9PCAS+mzzh21HBdfc896LLWDeh9CsYA/eP+uyj9wLJ1+zGAVb89hktnlD7EFHxnFLi5WXN6T2KgCKgCBxNBFTD4miir20rAoqAIqAIKAKKgCKgCBQnAvxbF+PE/Cn+hhA7NoWT6OTFx7nLaf6CahsU5xjKYt2kS1oW1HHS+oQiK4hqGSeG5sQaMU6Rr5BUULv86aB8TvMgI93TQbFE0j4hGm30IALvK4vAFWGfWcusadY2azwwcsjsAfYEe8PskyJsvuiqCo+IiEwRsebgGq++8bZ7SAc16ftvvw78rk2HLifslqgEnJi59YKUP8sXzf/LiCzndn9evu8j6ZuI2HjrpWf+F6yRgJ7CwLc/HsH3pq4oEdLgvSEkOKH9yDMvv/HbjCk/IkqNyC/6DHlpOy/3FKY9g9P4b774NJRQeQPx9uIkDaWRENw30g8hHoyeQF76nds9pM8h+qFGzTrHQRr1e/bVt0TXIPHjd14jQiqrmPaCo0O4Ab0R0lSN/mLY0GDRcEkB1I57fpsx+cfc+lIc38sWgMS1EoTgQjx77+5dO4PFmPmeVESsJZGkQD/HQhi628mnnYlofXaputgzi+b9+XuofpfUuAu6tiBw+B3IC+ak+0IThznM7hnmH4J07aqVwf8Ns1pKmjfWFpooP40/nPCoLyQSZAYi30S5BPaHNFOQkAvm/PFrKM0MxsD9GXkYh2yXqFqS6oz7iRALNW6IQ0NW5QUXvUcRUAQUgdKIgBIWpXFWtE+KgCKgCCgCioAioAgoAoVFgBQ+OMKai10jFuOvEO0CU8h7T154TpibtEKFbVefPxQdMVAskBwCF5zmOJ5xomOcPOeEP3nwpwlBsVpsj1hOEQ6Kb94QMGm5WNus8UCNB7MH2BPsDfYIeyUnUfG8tVoMd+EAjxDSIrBqtCu6dD+15/ffjByO4zbwO1K2ZCemjCOPU9KB99uEIJCDz0WSCg7n8N2PPPn8r9MnT/z8g7cRfz+sTB4/xkeudO1+2hnmi7DwcDR2LHOy+oob+t7VtGXrdoOefewBrpPiKC8EQF6hL2h7OGpNBMWo4R+9F6o9UkL9s2olei6HFTQBzMl08wW4k74nO62BvI4n8D4RKF+P6PaFkmqK/P7vvPxs/+BIit07d2znmfjKVdCqySoQGQ89OfA1ImLQDQluv0mLVm25Nvf3X2YUpG+FfSYzPd0XAci4ILy+lLRawaQK3wPpkvlzZnc56dSefL73f8++xNp644Wn+oXqA+mvmko0SnZ7piTGXZi1JZzUQfl5yBPpJVEpHWlr9qwjxbgNNo1EcBuyM1SkQwe/wPdMST0V/P0pZ5xzPnVM/WHcEanETujR82yISHRRQs0BY+A65Gxu6wRihLpY16GiwiBHsFD7MLe69XtFQBFQBEoTAkpYlKbZ0L4oAoqAIqAIKAKKgCKgCBQVAqQ+5RQi4sy+nNNSgtP5/CXX1orhLDhMdNic1C+qzpSzekgtNEEMIgLNCSIuwJ5XTsIihkxap9fFnhdbKCSFip0XYpFks15Z06xt1jhrPbCYvcDeYI+wV45IF5xNqrVC9DT/j5qc/JyM5mlSoTz16jsfccp56OsvPRtYI87XVu06dQkWoTX3fDzmp1mvfTjiW5yWXIP4wAk5949ZhXZC45R/6d1hX+4Rj/iTD9x2QyjdCunyAa6nyvF+06fU5EMn5ymk+Xmg/4BXvvrkg3fWr139N9cqSh6iHUUYYVHQ9iAC0H7AsW3SDgVi73S6XGiH7Ni2hZRuh5XHBw5+79OxU34zJAEiz5f0vqEvp/qDha3zv0L+ewJHM2Ll9wuGaJuQYie4PpMq55Qzzr0g8Lv+A18fQjqpl5546O5Qp+A5eU9qrp0S7pJdH3EkQ+qwDgszjlDPGpz63tfvSfo3ctiQt7Jr4zdxjIv+eZM7H3liAOLvaHiESvfkW3Nt23cKExYruz2Tl3EXdqyFWVv8PrDuGIPpB/Nw3iVXXvv0oHc/Duxb89btOvL5rz9+mRmqz6TcIqIJbZBQ30NIcv3Hcd98Gfx9u84n+AScQpEIbSWChe+yw9hEZARHerXr1O2kAa8PHQ4+pj2jEzN+1IhPQ2lwGFJR+Iwj9mFh50mfVwQUAUWgJBFQwqIk0da2FAFFQBFQBBQBRUARUARKCgEcRpXEfhVDw4ISeHoRDQRSESHunKd0EiXV8bLcjhAPlt9IR/SCGKLaV4vhECZyAqzXiT0lhsNtntx/RLqfsoxBKes7eLPGWeuseVPMXmBvsEfYK0XuZC0KLIzew1OvvP3hVZIGavh3U38XOYH6Lz350N3BzuNax9U9npQpOPlHTvxlHhoJgX34ecrE8R26nnTK0K++n/beiO8mvT9y3JQt4uUmH31h+ooA+MvvffIVpAX2+fjps0nrdKKIU9epV78hp6JJN/T28NE/QFhMnjA2K8e9+NhJhWY9OmDQ29KvqRvFWfreoAFPZvVHyJXExAPspyIpBW0PIoAOjPrsw5DRFURQQFogBhzc0ZmTfxgH0fTRqIkzB380cuy3M+Yuj42Lj3/9+SceKZJB+SuBjIAUkelwPH7PzdeEEmAmFdAP3371BVEKDz418DXm6NX3P/vm/Mt730BkxU/jRh/hjKZ6xJgXCgmSU38Hf/Tld6On/bn0iwkz5uD8LsqxSRCQL8Kies3adegnKbCyq3/qxO9GM/a+9/Z7YuumjRsCRceDn2koWhdca96qXYdJc1duCo5Aysu4CzvOwqytn4Q8kExPsfw+oA9z9U233zt66p9Ln3/zw8+D+wVhQcRWduni6h7fsDHEh2TfyiIRTR1cb9a6bQdIK/RXgusmKgpSaPWKpYuDv6tSvWYtrq1fs2plKKwQ4oaQekx+A1iXaGEMGTlu8rBvJ/3SuHnLNgcl7Mc8B1ZEJY0Z8ckHoeoyhEWofVjYedLnFQFFQBEoSQSK9D+iJdlxbUsRUAQUAUVAEVAEFAFFQBEAgRCnwDk9TW5+Ut6Q9sMnahtQOPWP8xbHWqLYEdEViux/CHx8Y3cOOeHMRkwbB7hJ2UQkhReCIlSR6+gorJHn/5VXHDaI4YI1uK8LFVUh99IO85aoURf5X4VEWgTtB/BmjYM5ax5iokNAzeyNVmJEuLBn2DuH7Yf896JonxAB5wXffP7RkMuvu+UOThxLdpvkFx5/4I4Jo7/8LLglka7YhkP6RtGR+P3naZPIGR94z6BnHnsAsoPIChyXCCiTeimUHkN+RtG1+6ln0DdSVM2a9tMEnPdnXXDpVb1vvuO+wHo4Gf/EfX2v+3vZ4qwUXTg4l8yfOxudASIX7utzxfmB+gqkfrlIUhx99Oarz+c1V39OfS9oe8IDRS2Y+8evwbn7TVuVq1WvwfsVSxcdIVbMXOEQv7LPrXfXOb5+w/mzf5s16Nn/PUC+//zgnNu9nGCHEHqu3z19IaKyu3/IawOfbi8n4q/re/eDGNE6rzzd7z7SLIV6RmRGKiI+TYqp7OokaqfbKaedyfeclMfxv2fXzh259Tmv34vTGr0fC8xyI9ggKWb89P3YU84894KnHry9D3smu3YEJwhN65FnXnpj5CfvvxUoEp+Xcee1/zndV5i1NWvqTxMgInHyG9HrZYvmz334tusumyZEQGC7RGmZlGCh+kNkBtcROA/+nugnCLlh7w5+KTiygYia+IQqVUNF9FDPPslbR+QR0Veh2kXk/e2Xnn38wSdfGPTWp98QnWhBfrzxwpP9fKm/ArQtJINcxGeSbi679V25WjX/PjxSNLwo5krrUAQUAUWgpBAolXlKS2rw2o4ioAgoAoqAIqAIKAKKQNlHIARhgeMVouIssUFiCUGjxOlEihxSe6wUJ6+KbeewDIRE4JBTrBii2aTdwNBBQCwYkWxOiOMQg8DIKobIkOchOs4VA3cc5q+IfSzf++6X7/mbhDobi6GnEC2GY2ey3OOLfvGTJvSDuiA1IE04BevOjjAJ7Et5fi/7A9xIp1RTjJQoRL4Elt3y4WGxSX7cD9MQgQQpDQXxXzk9X2354gV/5XR6mBQ2XjldnpPoLDneISlCpVQpyFg5TR8nlXL6OvB5HKRNmrVq4woPCyet0yJJpxQqNz76CfUbNW62esXyJZkiqBFYx5U33HpXgyZNW7zY/6G7QqWZKkh/i6M9HPZ1JQ3R5g3r/8kuzRMOcMZgBMYL0vfcniFtVV7qJyqmTfvO3YjIWbpw3pxQaaBMWziqL7jimj5jvxz+UU5zAAmCMPN6UWzGkZ5bX/PzPf28/Nqbb/9+zJef5eX0PFFGVarVqBkqfVdwu6Q6Ii1RcMRSXsedn3EU5N68rK1mrdp2ED3y6qRS2+iPWgpui+gD9n1Oab2atGjd9t91a1YHi7ITuQMxScRXqDUAoQGGEKHB7RJ1VTEmJtakecsOA0To6zdq0ox0TquEyCyIvkuYEBoShFM3t7YKMg/6jCKgCCgCJYmAEhYliba2pQgoAoqAIqAIKAKKgCJQ5AiEICxwfpOT/1ax28SChSwhMUingFP8oDhkD3O0F3kHy3iFQhYwAjCtI0YubURr7xRD+wBsOcGPsxsSCG0EnLaksIDE4LQ+Hu++YqSHop4BYmMQ1/ZHVDSUzyeKdRaDoOA5SCd0LhaJMT84202B0EBomX6kKWERgEyIt7I/ODVcUQwSjz0BORFYmLOhYuyJf/xzkPV9aSEsch6lfqsIKAKKgCKgCCgCioAicKwgoCmhjpWZ1HEoAoqAIqAIKAKKgCKgCIAAB3JIiXCJGKKqONQ5sczJfArpoP4Qg6xIUrIi90XjJwQgEkjvtMmPKSQFmNYWwxneXmyVGCLPG8UgGtCtAP84McSdo8TQryCiJVrqglRCjNREVxDFwVxRH/eifQFZQSoU0hbhWCdVB4RGclTNhp6mt79ptz5RwimnWWSNC2lBNAprnrXPHjBpocCbOWKvgO0IMVLElKq0UDmNT79TBBQBRUARUAQUAUVAETi2EFDC4tiaTx2NIqAIKAKKgCKgCCgC5RkByAqcr8eLISSKQ5xiyArSF30qRgocHLIaWZHP1eLXlUgVsuFVeRRBY4iIbmKkiCIVBlEPp4q1E+sthhMcpzjppCAhiNAg7ROvrf1zgJgshASvpJciOoN0U8wl0RSkkWK+qJsIgD3SD7n3F2vB7W86/BEEIedSowOyJtinNyLG2h/mx72TvJq9wV5hz7B3IDYgh5S0yIJP3ygCioAioAgoAoqAIqAIlBQCPlEhLYqAIqAIKAKKgCKgCCgCisAxgIAR2+aEuE+gVArOcuN4jZf3RAAgAq3RFYWYcCEMICK+EBss9o0Y4rkHxCqLQV6Q5omUUaeIoZtA1Av4Y+eIQVbgFCf1EwQGURYQEogkUxfkBxojzOUCsbFis8VIN5XuT1NlCSGB3gLzq6luBYTsij+SiCgL1j57gHmggJ3RTGDPgLcR386hRv1KEVAEFAFFQBFQBBQBRUARKB4E9B/2xYOr1qoIKAKKgCKgCCgCioAiUEIIBGhYREiTOMI58f9GiOZXyLXnxcaJAxfnrZYiQEDIAxzcRE9wWh+i4lExdCtwjqNNQaQE+gmIZUNSkBaKV+YA5/l8McgOIix+Ftvj7xbXkow4dxF0tdxXIXuFiJULxZ4QaxYCkPvlGmmjFoul8r1GqZT7ZaMAKAKKgCKgCCgCioAiUKIIaEqoEoVbG1MEFAFFQBFQBBQBRUARKCYEOIjDKX2Em6/Jpo3v5PpWMU7layk6BMAT4oFC2i1SQUFQkPaJ9EKodqNPQXQ3J/o53c8zy8Rmin0lxul+tC0yhKDQVERFNzfBNYE7e4C9EIqwYO9wz99i6JboXBTfXGjNioAioAgoAoqAIqAIKAIhEFDCQpeFIqAIKAKKgCKgCCgCisCxgADOcE71Q1yQiz+4EF2BExaNBNWuKMIZ94tymxpxcOPoRnh7o0RfkN6JCAzIC+YIQ1SblE8QFAhoc+p/9yFdCi3FjABrnz3AfLAngkkL9g57iL2EsLqSe8U8IVq9IqAIKAKKgCKgCCgCisDhCKiGha4IRUARUAQUAUVAEVAEFIFjAQHSESHUjIOVFETBZbVciBPjwI46YUtgxoWsYB4Qdj5ZjHRdpITi7w9SPqFJwSl/IjOqMTdyvx6mKv55Ye2DM3uBPRFcmDPuYS8ZQe7i75W2oAgoAoqAIqAIKAKKgCKgCPgR0D8KdCkoAoqAIqAIKAKKgCKgCJR1BDgRjkO8ixgiz4gIBztb0UaYJkbqIU1zU8wz7icrKkkzF4shxM3JfiIqiL4YKfah2CYx0ngxH6kSYaFEUjHPix9r9gB7gciXC4KaZO+wh4h8IXWUpoUq/jnRFhQBRUARUAQUAUVAEVAEAhBQwkKXgyKgCCgCioAioAgoAopAWUeAU/voIrQR4xQ/2ghNxSAxTMHxitBzoogIa0qoYppxISogjzil317MRFcY8ghH+XaxlWIbhaDwaVYUU1e02hAIsPZFeJtUT+wF9kRgQWSbuWEPsZdmiREBo0SSriZFQBFQBBQBRUARUAQUgRJDQFNClRjU2pAioAgoAoqAIqAIKAKKQDEhgJMcB+wWsbZi5OE3ZMW/8p7T/Dhhd4vDVh3kxTQJ/mrBuZvYRWJniuHsRq/iD7GpYugnXCZWu3i7obVnh4B/D+z27wn2BnuEwp5h77CH2EvsKfaWFkVAEVAEFAFFQBFQBBQBRaDEENAIixKDWhtSBBQBRUARUAQUAUVAESgsAnI6PLgKDuBEiTUQO1WsXtANCDrjkEX8Oamw7evz2SMg0RWIaV8p1kOMiUIngSiKSWKfiPUUu07M7vbazr3jwl6fzdkdx6l+ijlIRXoojCgY3/t5v36hsBc9AuwF9gT7AzOFvw/ribGXIJmS/BEZh0UlCelR9D3SGhUBRUARUAQUAUVAEVAEFAFBQAkLXQaKgCKgCCgCioAioAgoAmUCgRBkBf3m37OQFZwMPyfEQEhr86vYfDGc51qKAQEhKxBpvkUMUoKUUAeFbZgvxMTmHanhX87eFbetY8L+sdUj0lp6vFZ9p917c52o1MgFe72TMjw2TvtXFUM3gQiYWDFSR5GOKL3DSdcyb9nqjiihUaAJBdM5/j1B+i60RgILe2m8GMQGKdbSA79kLyppUSDc9SFFQBFQBBQBRUARUAQUgVwQUMJCl4gioAgoAoqAIqAIKAKKQFlGAOFgnOWrQgwCp/fdYnv4ThysKrZdgJkWwgANCswj5ICJiPDVNOCqM5xVwtPivJb3XskddKEADFmR4vHaqv19IPr9Zfsr7t6d7qoon8N/3FLF06BC8uQuCfsedNndkXFhGWe3r7R/7Z+743bKM0RjdBRrJYb+COmjIJpwlJOeCL0F3tO+77S/9MUrfSNlkc5rPueVvSCkA3jO9u+dE+S1WlA17Cn2FntMiyKgCCgCioAioAgoAoqAIlAiCChhUSIwayOKgCKgCCgCioAioAgoAsWEAM5UBILJux9c/pELOFxxaO8WB61NSYu8z4KfDKgkT4AxJIFHroHnXv9nK8W9MyHDa3/Yabmv9HotT7rXnp6c6TiwLjFq7dw9sZ0lwgKnOGLbXnm/ZvXBaG/ViLS19aJT6ie7HXUruNztK7rc2w9mOI6XewJF0klJ9K1YI7HPxRCDph6Ii01iSdIXBmOXV0gMiAsjDn0YgaERGEfOOXvBP4cJ/j3CXgkmLHrLtYViC/K+avRORUARUAQUAUVAEVAEFAFFoHAIKGFROPz0aUVAEVAEFAFFQBFQBBSBo4cAugec6G8ndlOIbhAVQLqb38XcSlbke6JwYBs9Cf5ugLgAc5zcCDLz+WxJ8XSxRFBEprrtO7elhm9bvr9CyqbkyGbyYLh8j5YFERR2y2ZrIXbaH3srt7Js+6yaEclWjMsT1TohLX72rljL4/HJVqz0ejxEWCDefZW/xy3k9UcxyAranCe2Toz0UXyGsIDMWC+2SwyS5DDNhXyP/Bh/wB9hAcFj9givweVmuTBM7Gsx0nUppsf4utDhKQKKgCKgCCgCioAiUBoQUMKiNMyC9kERUAQUAUVAEVAEFAFFIL8IcEKcf8vWETOCzcF1jJILa8R2iYPWnL7Pbzvl8n6JWoAIgKwAN15RWQZrBM7RlqgQ4fDE70oLuyDc7omxh2dkJrmd0Qv3x+3amRLW2GuzHHa7wy2poiJtlq2Nze6ob3c4ZM7ki7Aw62+riuSN2mPFutKsOGeqVTXKY+1IoUmbCwrC68kU81gStUHzRF4Eaix0lc9ok0BqcAfOdqIuPvX3jwgQCIxM0kaVywnMw6DZExJpAcHDHmGvkJIruLC3mPf9YhBEimcesNVbFAFFQBFQBBQBRUARUAQKjoASFgXHTp9UBBQBRUARUAQUAUVAETh6CEBY4Kj+V2x9iG7ggB0hhmgw0QBa8ocAJAGRCghgS2CEjUiWzpbNXkPe/yFsQqcIh7tGmN1r7U4Pk1RQzqR/0uJ/OeCotF7IizpOm72tMzwiQh60hLg4aHc4IT6cmelpVlh0RUn+FG1tteKFvthiRXq3W5Wj7VZKVA2Jl3A2cGekW+6MNMvjzrTc6anyPl2iL+TxQ+wFBQc6otCkiZopVlcM0e4TxRL9/V4hr5uFeEHQ263ERbaTz95YLYZOCITFFUF3rpfP7DH2Wo7i59m2oF8oAoqAIqAIKAKKgCKgCCgC+UBACYt8gKW3KgKKgCKgCCgCioAioAgcHQTkJHhww/w7VjzfvtP+6CwEFx7g+l5NBZX3ORMHPyfqiaI4TixNCIfGNrvlFNJB3jvOdjjDjpNoicqejLSz0pyRkZlOz9wMj+VZkxrnTnMlOBxWxjWO8KiGdqfL5nC4hGOQLEI2W0X5bNltDiu8gvBMdschwQl7hLU3M8aqZDtgRYa7rDBvuGULi/KlhvIKQQFhkXpwr2V3ZViZaSkigmGiLiAuvPHyPwhFQ0jQV9bCyWIQFTjWiQiYKzZJbDU6F0paHLkOAsS3a8u3R2wy/x6C1ABfIiwgsXyFPSnP531x6Z2KgCKgCCgCioAioAgoAopAHhBQwiIPIOktioAioAgoAoqAIqAIKAKlCgH83aQDqi6Gs/q8EL0jvxBCzhtKVc9LYWf8JAVEBVEVcWJNJDCisTPctk9ez5TAhk52hzfGGemqY3nkNo+3missooLHHm5tzrROSs/wulJsETVsmRmNJZJCeA2n5QwLF6IhTIgJskDJ/wrr4csmJO99JIbkihLiw5YUVs3aKERFtDPJipXv8IxnOpha0kK5fcSGVzrA+4y0NCstaa8v6sKnd3Eo4oK5h5xAX4FG1ovheEdno7JYtBhaGjjaNS1Y6PVn9gqvwQV8R/rxI3pF00KVwj1c3F1yucLCatc9vkFYeHj4xvVr1yQnJbEWtJQSBJifhCpVq23bsmljUXYpJjbOdxjgwP59pNkr9hJbKT5h/949kNDlrkRFR1fISJf/y0jPIoXLHQg6YEVAEVAEAhDILt+vgqQIKAKKgCKgCCgCioAioAiUZgTwVtcUQ2y7YYiOzpdrnLZHqFlLEAJCUtj8hjMfpxRpltqINRLeoLkwBRc6w2yDKlS293GG2Vs4wmx1qtT1WtWbeDLjalhRLpdbIibcVpKtoistPN5yRsaINkWE5aoQa7kioy27M0xSQQl5YbdLQMWhV/kfrxAXXq7LNbgIX9lni7N22ipLWIRTWIf//jwRQsNyRVX0iqWERVV0R8ZUssIjK1rh0dKWRGyghyEFMW/SVjEGjvufLtZWjIgACCvSRLUUi5Lx6mGt0DuBPcJeYc8EF/YWe4y9doR+RYjIp9At6NXDEOj/4hvvP/TUi4NLOyyS/s3W995+T0xf9M+Ob2fMXf7VT78umLV0496X3h32ZUKVahDGWkoBAtf2veuBUVP+WJxdV5irmUs27D6hR8+z89PdF98ZNvKZ194blp9nCnpvizbtO81cvH7XKWece0FB6yjLz7383vCvPxs/bXZZHoP2XRFQBBSBokRACYuiRFPrUgQUAUVAEVAEFAFFQBEoCQTwVGOc9s7uNCZObA7s66n6oBnxR1QQSVFNDP0H0gHxuanYaQ6X/a2KVWxnVW3grZlQ177zuHYZ7vqdUhMT6qbui4z1Ol2RNntyaobl9kjkhKRwCo+OlVRPYkIkSOSF5SCyQsgGXySFZSM9k69IlATpu7KIisBupUsQRKoEeHiP/FpIDptkk3JmiGi3BHVI2ihJNWUXy7rV6+VvGiCNztsAACAASURBVIwIAcZDqqjGYpAxRAi8INZXrJOMPRaipiQWaRlqgz3CXvHplYQo7DH2mtl3ZWhopbOrPc+98NIq1atDApXq0ve+R5+885EnBnz/zcjh1/bq0fmKM09oM/j5/g93Pfn0Mz8dO/lXcwK/VA+iHHSuQ9eTTkk8cIBIs5ClTYfO3SRYIt7tlrx6eSx2KW07dTspp3rzWFWebmvVrmMXbsxIl1C6clgYvwRXlMuxl8Pp1iErAopAHhDQU0Z5AElvUQQUAUVAEVAEFAFFQBEoNQgYsW3S/Vwrdn2InqFdkCyG4PYRp8JLzUhKsCN+Jz3Y8e9/ohGIREgTMiBDUi5VkPc3ivWULE1WTPUwq1pDtxVTLcPrybQqCTngiK6UUiEtOdUKi8y0HBIx4RGOIHmfzcpIzRRLtiIqxvlICo9bIi9EyULkKkzJ+ntDoixydMaEICuoAyIC4kHe2S2H3eX12NOFJ6ngI0QyJT1UgBj3oTZttjC5BmFBWiic7c3F0LeYLsZp4XFimtLmv/XHHmGvsGfYO52Clubj8hlSC3HurWKkLNF9FQRSXj/Wa9i4aVx8QuV1q1cR1VJqS+Wq1WvcfM9Dj3/z+UdDXnm6332mo6tXLF0897dZ07+YMGPO/f0HvPJcv3sgA7UcRQRatu3Q+c9fZ07LrgtNWrQi6sxa+/eKZXntZoPGzVqQpmjJgr/+zOszhbmvUbOWrXl+2aL5/AaVq1KlWo2apMNaOnbUiHI1cB2sIqAIKAI5IKARFro8FAFFQBFQBBQBRUARUARKNQIh0s4gclBLjLQ/weUTuTBcbIkYp8bLvWPVT1aQQ6mqWA2xBuLUbyjEwhkSufCkvI6wO+09JVOTFVfDY1Wp5xYNCnQjPDZnmEeuOqyoOC+WJFISO9LErR1R0WbFVk20XBGpkgrKeYgz8GlV2AirOLJ4vYtlJgp1ehQdjLDoihkS0ZHhDI/yRMTE+6I7SDkFScIrRQTC6QcfILUgLkwhZRQRFz0FE1JEaaTFIWSYPfYKe4a9wx4KLuw19twhgREtBUagTfvO3Xh45dJFCwpcSQk8eEaviy4PE9GKT957/eXg5lavXLZk+NC3BvW67OrrcbSWQHe0iWwQQFvE5+zOgVho0qJ1W3Qodu3YBuGYp9JCSBBuXLpwbokQFo2bt2qzeeOGddLNPXnq4DF0U+PmLUnHaC1fsmDeMTQsHYoioAgoAoVCQCMsCgWfPqwIKAKKgCKgCCgCioAiUMII4GTGQYYDNZSjbJtc5x5EQkM7z0u4wyXRnDjfs2uGA0rGed9D3q/lRnH+VxWnfzeHK7y1EBNyIXGD3e6uW6tlmlWpdrKVmeYQMsBrRcenShSDM13SQGWEV/AetNncBzYvi0yKqpRSp1LtVEkP5bX2bo0WwkJCKyT2QpI3kV7o0KEor/dnaQhR9OPltbWQCL6r/vkpECwSxZHkCA//y2tlxogAeANbRFikzRYZnZmeKdEdZDvxcxC05fUS5yGBG7Z0eS+hGD5ti45i9Ilc4emCm2fer1+Um3WSA+hgwJ4BQPZQcAnccxq5VKDVe+ihlv7UN8sXL/irENUU+6Mt2nTolHjwwP6tmzZuCNXYlAnffYO+RdOWbdr9+cuMqcXeIW0gJAJEV/DFkoXZR0I0ad667RohmfIDIfWmpaakrFqxLFttjPzUl9O9Qjg7GjVt3urnKT9+X1R1lqV62EP0d9nC8hddUpbmSfuqCCgCJYuAEhYli7e2pggoAoqAIqAIKAKKgCJQeARwnpLCiDQ/wWWGXCBlzTqx8q5fAXFA+iciDZqJnSukwVKJqugur+e6IqIsZ3ik5c6QVE8RjrqVRaI6vIJDNCgyJfWTJy26ksdWsUqm0+vJcNgcXqdwABGRMZkJUZUyDybutJKc4V5ndHxmpsPlXXdwV1jNjDRXZYnA2GOzvDuEJKgpru/fhSioLO8PEQJeb6bEbaQcin7wRUDIJe8G+cyp/Xq5LAvqYDwbHU7nAYczOs0R57HbpGN2Z3Kb/duiwjPTXFZa4gEiQ4SlkP8TDkXSRtnkM/UHRga0kT6d5SNUDjnnITPKe2GvsGdID/a32P+CAGGvgdUrYv+Wd7AKM34RF+64c/vWLVhh6inuZ+XQfmWPlOzaITXU9Ree3m3J/LkqFFzck5FD/a3bd+7qzszMXLFk0fxQt5F+rHqt2sf9PHVivsiA1u07daVO6i7u4dVv2KRZeERkZGkn8YoLh2Yt27RPSkw8uOGf1fz2alEEFAFFQBEQBJSw0GWgCCgCioAioAgoAoqAIlCWEMBpzSn9/1QS/us9jpVVYtxTbtJBhYiu4JS80X5AWLuDWB0hBq6xO8MsV2S0LxoB4WqJshByQoSzKzityLhd1sGdCV6HMykptnry/oiK7lib3RsmmZiyirx3RMZ4Mlzh1lohLDIj9tucRFdEx+/buXuDfU/SvuhouRndiAghJS4U0oKUTIdqgJjweNOERNjrzszAMSNZnFzJInhBmqbcii9Aw+5wN3OGu6tYNu+2Cgket81yJ0dUyJgUFes6effG8DiHM8FKPbjfp23BA15vyKxPLrn6P7kB/Y7vBD/WEo7Zw9KHSeRFbn06lr43aaEgI8CCvRT8t+KhiJVD86lRKQWYfZcrLKyhnCT/dfrkiQV4vEQfIYVQRVHVxpHMSftQjStZUaJTErIxInaIgshujpq3asvvv7Vq+dJFee0t2hVoWIwYNuTNvD5TmPuatmrTnufLK2HRtFXb9n8vW7QgJ4KwMPjqs4qAIqAIlEUElLAoi7OmfVYEFAFFQBFQBBQBRaB8IoCjNEoM51moU/Hb5XpDsc1ixX4qtJROgSEr0KyIE+Nk/NXCFpx8iKCIFH2KcIlCEF1qn+9ZMiY5wsV3H2elJ7kOuDPDdkfGZURUSEgWbQrB0CtYi9/fjztDTrHbvbtEnPtrkYpoGBnrcUXut3Yk73PWiYxN25WWHH6WpJBCoLmyEBOp/uclEsIOkSHC3PZod0b6TmEqGkkakHi5kiddC588hsOTapd4D5vNm+IMczujYtOdNsuzPTrBvkBok7Dw6ANd9m5xVtq9IcInyG0JWeFNT7HsLhmrHBQ/lDLKV8KFqGgiNb5jd7ogNiZKnw4IQVHe9U4ACIFztCrYS7wGFvYce489iGi5khb5/BFo2LRZS0iLpQvnzcnnoyV+OwLNsjds4rduXVLCyyU+yDLeIBojTVu2bvfdV599nN1QmrVu5yMs8qOZQjow0jTlpItRlNA1b9Wug/wme4WwKHcaDrFxleJr1al7/PSfvh9blJhqXYqAIqAIlHUEVHS7rM+g9l8RUAQUAUVAEVAEFIHygwDOeBzcu8SuCBr2XPn8hxjOVIRFyyNhAT6GqCBtFpELXcW62x12y+50Wp7MDHHcuyXtU7hPsJpXcUx5M9PDrfSUyAqRMWkJmWlhLneGK0MqOyB0xnp/nebUfaSIc1cLi/JeIIRFVUkHFRlXM6leREyqJzUxvK7d4SX1FKSRkCW2Sh4JdRCygEgGQzC5JaqithAW1aEv5D6JxMheGJ2oConyOGB3ug+ERWRMdbjcfzrDMxMTjtuTWiE+KUPYhiiv13W83LYg/rjUPU0kzqJWs/0HKlbxWM4IhLilCWkGogZy4rDi9Vbyetyvyw1nyfd6kOvQnmHvsIfYS+ypwMKeY++xB1WwvAC/u01aHMpVX1KO4AJ0MeuROb//PJ0PXU8+/czC1KPPFh8CRCZAgOVEKEkKsk6kdVqzcnmeNSxaSTooer1kQckIbjeTKJAN/6xZlSSiKcWHVumsmegKeqb6FaVzfrRXioAicPQQUMLi6GGvLSsCioAioAgoAoqAIqAI5B+BGHnkdLFA7zO54DmZSWQFeg3liqzwpy7i3/WRYghKnyRWR+xEsRskusEWFhVjRcTEW2HRMT7HPeSFMywiU8gKFLdtpE5K3hdpP7AjxnlgR8Wk/dtj3PLZmZHiwkG9X2yTGPog6BjsE8NpvUO81uiF1AuPSju5QkLSBWHR6RAMvlmVw9nhQogkCDlBpIfMiZd5IaSBuYPAmCwWqC2RtRqow+70LIyISVkRW+3gqgrxyb9UqJy4TIiKpIS6e9NdERkuZ0RGTYn2qCwki7t+5+0tK9fdvyu+dtKuxj32r42rkeiJrZZmhUWJ793rtdyZ0i9fnw7/80fIlKoed8a1gkPVE8+5J1Sasfyv0LL9BHPEHmIvsacCdRaYN/Yee1BLARDgNDwnyZctmn+E4LZoszhPPavXRdVr1mbvHvVCFMieXTt3nH7O+Zcc9c5oB0IigM4EXyxdkH3EDmTAahHcTk9Py1M0G/VR7+5dO7ZnJ7helGuVSA5Ep2VPBBOkR3XWiXqoL0rgxd0JCCXaWLZoXqkaf3GPW+tXBBQBRSA3BJSwyA0h/V4RUAQUAUVAEVAEFAFFoDQgwL9bq4hdKfZ+UIdqyuezxXB+bxTD6Vpu0vuIBoNJlRUr424ido5Yf7EbxEPvIyiEnLBcEdFWVKUqVlRcFd4fEEJB0voQw3CoQFqkJ7ui9m6Oq7tjbWV7ekrY9rRkV6w7075DvoaYyBAjJdBBsTSP235AhLYz0pLCtqYnh9ncGY50r9uWnFWfx50oaZggNyAvRMzZJ7R9KA/VodRDncVwgmf14ZBOhZAVdm+i2HoiJ8Ki0jdUa7hzW7WGu1aFR6eviIhO2yf37EtLCt/mDM/4V1JQhclztcIiM3eKrsYi0bY4eHyn9OkNTziwpmqDJCu2mtOKjo8QsiZaCIwKh6ItHIcFVJwiRMal0otIwbI8Rw4wL+wd9hB7iT3F3gos7D32IHtR/5YMAie3j206dDkhu5Pkz7425JPBH40c+9BTAwfnVk9JfC+RWO7JE8aOatKidVuctyXRpraRPwTQryAqYf3aVStDPVkpoXIVCLD8kgHUmxMJUpRrFcFtkUmJWrrwr1KVJm3g2x+PGD3tz6VPv/rOR2HhEUQCFktBY2T/3j27N21Yt7ZYGtBKFQFFQBEoowho6HMZnTjttiKgCCgCioAioAgoAuUMARzbnDzGYY5jPrjwx/5IsWViONaPuRJCXJsx4jRGH6KBGGmg0B0gxYSc2hThB8nb5HC5LI8nE/0IE2GQ5M5IWyXf2eX/JX2TLevEPKRFRqrT2rc1Nl1Iiw9iaxy4SogIl0RPSDSGN0NiMZZK9MNeUZJIT94fWXf/torVE3dVyBSiIyxpT1RkaqLoR3gO+fyl/gq0b4ocLMcZnizkBZEgRjzdLe+zbpKUT0IoZFrRlZJ3h0eneSMqpm2Nr7M3LSo2paO012nbqio7XRGZadHxyfWcdndiSmJEgtvtiKxUY79Hnq0r/YsQfqZS1YbuNEn3tDH+uMxdG+aFd01LirQS94RZIgwuabGsw9qUPoaLhkULT5q7i/RlgdieY27x5H1A7B0iK4iAQTC9XtCj7D32IHtxr1ieT23nvQvH5p0IGTdu1rL1T+PHfBVqhPGVq1Tl+rpsnM9HA5WJY78ecVWfW+8+//LeN7w/+MVnjkYftM3sEWjZtmPnZQvnzSVqJ9RdzVoeErPOD2FRvVbt4xIqV60m9WZLIBTlWv0vwqB0RVg89eDtfQa88cFnF111/c216x7f4LarL+gJiVfU6xG9kGWLFxwRcVXU7Wh9ioAioAiUNQSUsChrM6b9VQQUAUVAEVAEFAFFoHwiwIl8nC8tsxn+UrmO4xtn6jEnBpwNWQEzAC4QFecLRXCORBp0E6ZAiAVUqsWcYSKeHSmRBRV95IWURIkm2OKKjK4g3xJhwWl60khVDMTV47bV2ry8epPdGyutC4vMiKvVYutSScO0LuVARBWnyz1PUj+lbF1Z7UaJrqiavC+qYma6I8LrETLAnX2AgnRHnOE25ofT+xBQOH+YK0NYZEgbHiEnHJL+KVVIi7j42vuqy7Xq8mw8cRnxdfa1Sj0YXlfSVVWQCIy41ORwyA0EondIxEcFh92N0zfF4bDC3V5rh8PptVesnBERVzOjQaUUW8WIKJe1aWm4w+N1WDYR5valiBIFcnemu6+EmKC98YlgPR6cJNVWkTunSuPWbVcnxlqwMSt1PPPBHDEn7ClSQAWXtnKBvyP/FlPCIo+T2rp9526kv8lO/Pihvr0vqVajVu31a1eDa6koS+bPnb16xdLFl/Tu0/fDt159Hi2EUtEx7YQVWyk+gciXSeNGhyTAgKiJpFriNT+aKTjQfc/kEPFQlGu1RdtDGht/L1uysDRNK5FQfS4+48SHn3px8NU33X7vDbff98gn7w5+qSj7CPEDQfT9mJGfFWW9WpcioAgoAscCAhrGeyzMoo5BEVAEFAFFQBFQBBSBYxsBI84sQs0+EelQBedykthhZAXO2GO0wAzg+OcV8WkPZAXpn8KjY1wRFStZrsiKkgoq3HKKsLZoSWy1O1z7xEG/RyItJIWSPVaegeioK0aERnCpIATAVSn7IxpKFEXCyp8bRi2Z1KzjP3Pqnblm9vEnrpjRqMn+bTEO0bsIS09xxUsURqXsyQpvspABkhrKR2bQFuk1cIhDlEBc+NJESXREpuhWMNfrpb7NolvhkGiNmikHIiMl6kMSP7mPq1g58fjImNQYIUqSDu6K3pWeGPZPWmLYzH1bY/7P3nUARlW02+0tvQdIIBB6BwEFUcECKnaw4Y9df7s+sfde8Vfs2LGhIliwgGIFRRTpvQYCCaSX7fWds+TiZnNTEERYvnlv3u7eMnfm3Bkf+c6c7yxEPzZBIcKAqhmP0uuNmr625FB+6+4Bb3peoDCtbWB5WjtfcWKmDymhdvpZcGNyeHMy/zcUnltHo3KexYG4OFg9LbiGuJYaI2yIEzHie5S/J1v4H5h+gwbTW0azdtXyJWq3uJxOx/5EVih9/Oid11/KyGrVmv4aLRyqXLYPEFCUCfQaaexxXXv07ud0OOwb1q6i8rBFhe3W+aw06qmwN+cqCRJ0b6nX46aqa78qVFRMeOD2G+kBMhakBQnHvdnBXeqSJt7h3nyetCUICAKCwIGEgPwD80B6W9JXQUAQEAQEAUFAEBAEDk4EuJubu765k5T+CdGFqaAmoa5HPVh2ABOTLNQkKCkGoB5rtMbDoyJTY45PDvtWGJF2m94VepPJpzeYEhBsScZ1xEcJNJfjO1QWjabQqgABsBE1HQTCYNQBIA5yPU7TsUj9dIWr1nIojuWDVICzdVMFzMBOo20+l5+RpBKD4jT25q5yP0QPPqSh0oGc0MObwuu2m2n8neWotLXG91xUm99jsMEzwwKPje0+j96F9FUj3LWWEeiHDqQHO0LTaBp9p4LEiTNaQxqTNbQSGbFecZRr77Im+4pDQQ/SZOHRdYTFzowqIapVetfdS8VJ/EFKWnCOcC1xTXFtRReuQa5FrklR7Dc9+Xed7TtwJ2GxfvVKKlfqFe60zuvYuWtLmjIYkONtH5avpn/wrsNurz1z3CVX7sPH7tNH4b+LWhpJ79OHtuBhTb3rHr37D2ATyxYtmN9YUzSzXrl04YIgSgseF74EHMeALZs2rKuprmLKtwZld+Yqb27K/8FkMps7d+/ZZ8V+5l8ROWiSFh9NfvWF9MzsVsSmpTi25Lpe8ArhdU35hTTVTlx8QszuyGgJfnKNICAIxDYCQljE9vuV0QkCgoAgIAgIAoKAIBArCDCwTfNnqgKiC42duXOfOzRjzmxbJR0U/w3P4Hof1HZI9XQByIph1qR0BOYToKyI01BhoTdaoLZICuCYDwQGTK9RtFqa5zLIwZ2irDRrpWdD2Bw7qlASwdzaPE+ygTURCPdBzUFlCqWWFAbAq+suZN8ZPOO7ol8Cnx8OkIMYKfC5TdVQStiR5mkDUj95XNXWfs5qSz78K3KRnirOYzfXet1GP65J87kMh/vdpqN8bmOKVh90mGw+tqsoT0iicMwgMTRF8NgOmeND7ryB/pzOQ/0rWnfxL0C6KPAVuGUnWcHusW9MO/Yb6m2oR6EmkLTgO4iuLRn4AXoNweD74ZpSmxdcg1yLB0XKrN19hwwyM4XSi+99Omvq7N+WPfzsa+8yyNur38BDqyrKy8pLd2yPbvOeJ55/7c1ps+Y0FTQ/+viTT//o23lL/9hU7p32/e8rmEpmd/v2d67nDv2Zn02dMnDIkcPbts/v1JI2OI4x4y65YtKUz2fTuJgGxlRpqN3LNFgPPj1pcmTbvP+iq/7v1idemvzRkGHH0vxdtQw6/Kij73ps4iQGvpULklPT0m994Mlno9tUayApOSX1nieee3XuqqKaX9cU2y+99uY7WzK+3b2m9yGDBk9886MZPy4tKPt+8caSx154Y8qZ4y5VJYC4i/+iq2+87ZsFa7bN31DqphG70Wiimq5eYSqlHcXbtpaVbC9W6w89U3LzOnRUFBjdEWwnnq9+9OUP9CRRu4fETfc+/Qc0pdpoyVzl+yOWsxeuK56/vsQ15es5C/leop/ZpUevvlwvkaQL/TOuuPH2+2h2fcQxI0ftLtZq13PucR0m4oWrnW8P4+83p38zt7HzSxbM/5X3ZbfJbXbNHXns8SfxXT83+eMvO3Xt0aup/lNdUry1cHN5WQnTGoYL7793wguvX33L3Q8loEON3X/SmHPP/2HpplKFtOBc5rwn1s+88eHnHNPewE7aEAQEAUHg30Jgv9tF8G8BIc8VBAQBQUAQEAQEAUFAENhvEWBgnbuPT0LlDnilOPGFgWkGBXjNrsgzL4iVdFDwUtg1YATNGVTnDmsG+TuBgBiPdE9HkaCgqoKVXhWhEM2rLQsgVcjX63VIGRXGibF5BvQZ2CdZwM9NqDTq5neaYRNDEhQMLrZC7YBagEr8GTxhwIfXKmqJXX1r5AuD2iQrmJ+c7eahUtWxte65PMbAyomoOnhhaEo3pbWqLY3vCiWFPim7BkoLvQZpoTQBfJrjPduotPC5TBwL+1Gh9+k3IU3UIr0hwDGSjFE8GBhw5zGkv9LozXGhU6G0qAn4tJv7nOL7w+3QvlGyQc+goVpQ6Zq6PjM1kkKyxBwZpryzKB8LZR1xTSnYKGuNt3ANXov6Beqq5ibAwXSewdanX5/yKYPDc3/49mvuVD/+1DHnMjBrtdniFv0xb64aHqU7iosY0I3HjmlsbG9g+n7hlTfccv0dDzy+9M/f533w5qTnzjjvwsv/+3+333v/TVdfsi/wnfbem6+MPu+iy1mffuium5t6JsfBYG3PvocM2rp504btRVsLR5x0+lkkJMadPPzQaINoBl5ZV69Ysui91158hkHzR5597b0RJ59xFp8z/PiTTjvxsJ55xCj6uQzsH3bE8OOmIm3VmhVLFzNoS+JHUat079NvwOijB/VQ629mdus2r0396kfunJ/x8XuTu/Xs2//Km+584MtPPniXQeS9hetZ51921a0PPPEszdRff/6pRy0Wq5X97tKjT7+p77z2UuRzGLyf8Mo7Hx957Aknf/vFJ1NJqY48efTZI0454+wvp33wTuS1TCe0BPOhsX527t6rD7Ek+XDsqNPGPPr86++7XS6nEezHgMFHDCN5Nue7WV9G3s93hCmY1JR/RXNzleTRM29++Dnfy/czZ3xSXVlRTgLv/MuvHf/sY/fdXm8MmCP8rRAWfQcedvjTr035lHOI8+SUs/5z0X/POfmYBfPm/Lgn74Nz8cTTzzpv4fxffuZcjm5r2IgTT+Gzu/bq2//3uT9+F32+FnITHmtK0cB3d+ejT79Ek27lfhfYvluuvCA8j9UK3+H8uueR5Ll/wotvjBp9zjiOne+uzyGHDrn87JOYprBBocJGj5ugFAyQmHrlwy++J/lH7w2SHovx35pN69fIf5/3ZOLIvYKAIPCvIiAKi38Vfnm4ICAICAKCgCAgCAgCgkAkAjT/jaoMsDNwmoF6fxRaDEZ/iroFlQFVBuFjvSiEBc2laY56FNM+GWCsbbTYgnqjCf4Meg1SQPFYV51e6zLFe+baUpzlBjOtLiiyCHH3PNP6EFviShyJnxeVRISyE5oEBXeUbkCluTJ3+ZIoIVGgulNVBXz2lzvyqcYgIcLnMPhD0oUKCI6B14T/LkFaJ43XYdbYy+MCUFG4oaqoKd+SqgGBoYHKQlO5LXkzVBdukBUkJb7EWH4DUVEMvw22qygsSJAw6Mv5QNKChAifbUNyKrPeFCpJygrqDr/A47Qmhe7daa2hWo7D0RxUpt5iX+tdqSguGr37wD5B7Igp1xbXWHTaL65Fzh091mvjCB7YGOxW7xnMZACcQd/zTz1m8A0Xn33K+MvOO+OFJx+8K79zt3DQfNnC36neaVD8Pp+Xu6zVyIphI0adSrLii4+nvH3RGSOGPn7Pzdcx0Ly309M0NdhVyxb/uXblsiUnjxl7QVMqEJ57FrvLu/Xs0/+RO2686pQj+na67KxRwyc+eu9tDM5269X3kOjnKGlxFs7/dQ7PnXfpVTeQrJj09KP3v/ni048zEDz06BEkNOsVBnQZiGYwef2anWm27nvqxTcyEbS96/rLxv3603ezOnTq2p3B3Oh72eZTr743PRUE08WjRx7x6J3jr37w1usu16GQuNitF9/ExceccMoZtz004fmvP/t4yrnHH9H/nVeee2rypGcngETW//nb3J+ib73hzgefOOq4E09hX2696sKzb7/64nMZ8FfSPynXk2wh0bKiCe+DTl17hsl9p7229uGJr7wz9/tvvhoxoHObS8acQOWY5tyLr7wu+vkt8VRoaq6yvTsfe+ZlkhV3XHvJeTdd/p/RHAvHyvcanR4KAfnBdrzAApA5VCO88M4nM6kaIcl0zvFD+/F97I1UZCTD2DcSh2qv67Ajjx7B4xmZWSTpGxSFqHA67GopKTU7iaZ3p5GsIOFx1oghfT5465XnSQxRKaHWZrsOHTvTOF0xRL8XKqsTQKo88/DdtxzWKcv23defT6eqqTGlRP9Dwo8X7AAAIABJREFUhxzJe0kQTZoyYzaJsCvOPeXY04cd0nV4n/YZk1+e+OTemsfSjiAgCAgC/wYCQlj8G6jLMwUBQUAQEAQEAUFAEBAEWooA/73KwPmpjdzAHfU0HeWO/Rbn6W7pw/en6xAgZ2A4CZV5ry8E83AO4jlQVRhIVoR0ekO9f9vD0SHeZAmUJGY4Kwwmvz0h3RFC6iQoMELxOn3QpjcEjfCKKMHnGhyjKWuDnd04xkA1/RxYGLym70UznhVhBQUDO6WoCgnSBd9JspBoIIHBnftslwRJvUJbCXhjfIVUT6uQAmoOvvOZSqHSg7/Xoc9zkAZqW5sexUtSc6pc+E1SgqlhSKzwGfykopzP4Y5ppvUwg7TJBXHREYbcQ7sf40tIzAxOBL8TJnMiSgG+56FOQL0FlQHnvWq4Gj3u/ew31xLXFNdWY3nSuSa5NuVvSoBw+8P/e4E7+xmoXbl0EVOphctnH7zzhvJ98R+//aL2nhnIX7F4YQOTY6aEufvxZ1+heuCBW669TPEisEKu4fcH9opfz5j/XPzfo4474eTm5t+sGdM/TElLz2AwurFrrxp/5wO9+g88jH2lekBRUyg75OmpEH0vjvWnCoOkCNNcXXXT3Q8y2Pvy/x69T1EgqKWTatM2rwPVAD/PnvlFwO/3H3PiqaNJ7txz4xUXfjn9w3eZxorPUrv3/Cuuu4lkx/03X33J6uU7g9mI94b/uxZAY81h0ZLzTAPGdFXc1c8+gZPifws1/QcNPoKB+5++/erzyHb6DDh0yNhLrrz+o7dfffGTKZNf4znix37hVdfrExU8PL9iScM5o7SZ36VrD6Yfu+yGW+9es2LZ4luuuOAsmmVzblJp0TqnbV70OLpj174fjAT4H1VjeF7f2FzlORI0p5x53oVvgWiaCZJGaZ/KiuefePCuaGNtzhUqQACHlQH/EpAVVBRsXLd6JQky9rNVTtt2LcG7qWuomAHXUKMW/OcaQ/D/iMbmCo+TXOAn56nac0hKcQ19/O4bk64877QR61YtX2qvra7meiEBpXYPx87jSxf98RsVKEzT9ehd468m0UCcli38I0xutsrJbTB+ttupW8/eJOU4x2yQZl165onDfv/lp+95D0muaCXTnmIo9wsCgoAgsK8RkH9c7mvE5XmCgCAgCAgCgoAgIAgIAruDAAPQ3VEb2/X6A87NRmWQfFeJlXRQyoDqyAoG3xn4Z8qJs3VI/WSyJYKsiAMJoWu4yx0G1MGQzqM3BkK5vYp25B+2qaDHMWt+TW5d/XNSVu303N7bfut0+MZNrbtv/y0u2bkZxIUdQf9wmiVUEgssDNQMR2X+cQauSQIwzVNjQT0GdH5EZaoS+hxQTcGc/SQvGMSlZ4WizqASIpKMeA+/P0KlAfewuvt4bTiQCDUF+7cUOoev0deZCel2c+ehGwrb9t1mNlp8JEP4PAbaGGRfikrShMoQBgqZ5ohzhGoJYhgH+Gwdh/hNg8d6S/IG+L+xJISqQGQohe1xN/gZqON4fV2/Y1ZNoLJmiBfXFteYWuGa5Nrc5R/QyHUxf/iQw4YeNeqMs//DIDSDiJEDrsUOcv5mUH3pwoYpfLg7u1uvPv2VAGXkvRdccf3NDHw/fPsNVygBb6oYOnbt3mvd6uWc43tUuPv7jkeefomB/+YaYooiXkMvDbVrqWa4EL4T38yY/tHnU997K/IaZWc6UzZFHmfglWlsfkH6LB6/AUqSivLSEu4y5++mTKcV8mPu97O+osfD+LsfeWrW5x9/8N1Xn01r6l724eKrx9/OZypj4vVd6siUdatWLGsOi5acv/2hp16wgFi6D2m7aNys3DNk+HHH8zeJjMh2brjjwScqy8tKJz5yz63KcRJgZjAWDIBHXkv/CgakQT782VhfGJxPxFi7IvXUbVdfdK4yf3ifw1FbS2VD9L1UWKxbtXJZNLGgXNfUXOVO/5vue+wZKiRemfj4g5FtM5UZ1SWRxziv2+S2a79s0R/zr7nl3odhM5EzHoqMSLNvpq9S62dL8I++pmDDujXtVYztj0I6KGWeNeazQnKBuG1a1zDFElN+MVUaU3Y9csf/XUlSkWv0hNPOGss+/Prj7Jlq/aWyiORQRVlpyfh7Hv3fjKnvT/74nddfVq5VfEvUxt//0MOPpMLIbDZbmO7rzusu/c+Gtau46UCKICAICAIxg4B4WMTMq5SBCAKCgCAgCAgCgoAgEHMIMDjMf68yHQ+9BNQKPRgYeIlZf4GoQXOcDMQb4U9RZjBb040WK9JAhZUT4ZRKrExehCC+xoSad0hhanyqozWzYidm1XaKT3MsRFqlxUmtqoch8H9oMKh1umssWzf+0a60tiyuh8duSQ0GdsXl8/Askg0kAxjAVjwwVFNn4DyVDdtQqXagioIKCpIcJEH4yVRQJBB4nkQG0w4pRurn4fubqG0xFptOF+qHcbkNZn8hVBdlOn2oPC7VuSDo1xWl5lQmtepakmCyes24lsHWbFQal5Ig4Y5UfucOX6aSYZ+Z5qpn3XW8nuf/MFlC8entA7lIDeVMyw3+sHau4YSqIp0Fz4tUkVBFMB71A1SmRyIOMa3mwfhYONe4trjG1ArXJNemgWmhQHgcLGuwARaX33DrPQxUTnzkXpq11yvI3EOPGM1KKAhoYB19Hpl7+nHHfTSZwUD1WRdcdhXTP0WaEnMHO1MCMUVUI++lRYe5q5vGyEzdREVCczcVFmxcv3VLwcZBQ4cdo3YtfTaYT/+ZR3aSDZGFBtD87cHO8cjj9Fng7z9+nfNDxy7dex530hlnMY2WB1vrebxVnckxd4xHt6mk9+G9p597waX0PXjqgTu5TsMFPEjYIDn63tFQlMRhR/qLEx66R7mWWNNjgSRCEQbZHBbNne/So3dfBpKpLKCPR+T1h8NEfC0ICIf9r/RCNOUO+zfAHyRyjlx23S13URnw46wvP4tsg0oI+qM0Fczv0KlLNwa9X3rqkXujx6TmlUKzb5JAX07/oNG50NhcZd+YDim7dU4u1SRURjSHkZIKzAkcLr7qxttI1FBZodzHthj437Jp/brm2mrJ+a2bN24gIcN3H4n98aeMOYfvKKdd+/zGjOz5ztavXrFM8bJQnsf3dsv9j0/k+iQxpagaTjjtzLEkY3idmicGj/fqN+gwKl9IGtbWVFUx1VvkONq0y6N/lIbvOXp8xI6kF71f+N8BhfBrCQ5yjSAgCAgCBwoCorA4UN6U9FMQEAQEAUFAEBAEBIGDDwHF/Hc9hs7d99y9r/hUMPD3DCqDqeFUG7Fa6tQVTEfEXbrcRcn0Rk6kMEoP+r0avUmnscR7NCmtqzXmOK/GaPVpkltVa9LaVm5p3WO7GwTFAAT1cxD8RwapUDJ+D07PKx8KMiMN6ouuRrN/II6d0q5fYU52p1K7Oc7joZqhDk/+vUDSiAFDBh0ZqK8XdIzCnYF+5glnsJCqDJIDJCdIcFClsBaV5AVJBCodqODgmNgm320n9KnUluQqTMmpWp8/eNPnWR1Lf2jTY/va7kev3dG297Y0KEUqoarAWD0cFxUTJFO4c5sECXf8M0DMvvKTCotKVKZ0opcFSZIaVOJZjF70hdIiMz4tWJuRH9jcc4TvdYMppLZr+QRcPwqVxEfMqiwwtujCtcU1xrWmzAm+J65FrkmuzdDBTFYw9/6gw486GulYvlMzuVWUAGqeBQSbQU8GH6ONjoePHHUa09V88ObLzykvZQgCp0w/w93Yf/z6c2PKF5XXWP8Q0wHdfN/jzzCFTbTxc1M3L4LPBG4Np2KKvI4Eygmnnzl21ufTP1QzrOZ5Xh9NHnTpvtNTYOnC+fMuve6mOxf9/uucH7/5KzjfDlF3ni8s2MB5Vq906d67LwPxVZAlXHT1/9329qSJEyKNuXkvA8iFUYQBCR+qWZS0XUy5NGHSOx+nZWRlP3bXTdc0C14LLjj34iuuI/Ew9e36ptpM70MlClKD1TNfZ5+oalBSQfERNFWnUfST9956Q3SgnP4lkWnHorvE90OPC3qiRM4fXsfxkqDZtmXTxsj78tEvnmuq3cbmKts558LLr+H7nfXZNBK7zZaeCLrz/TBlEtUB773x0sTImzp16xH24FjbRHqqZh8ScYEyD+gxoxxWUpy9++oLTxOrVm0app+iUoXpl+gBEvk8kilMx+R2u113XHPxWKoleJ7Ez+XX33o3v3N8kWSjcj/xh61Nb2QJ844ASffkfbfdQGIqsv3OeCbnM83Ro8dJoo/PoVro+SceuHN3cJBrBQFBQBA4UBAQhcWB8qakn4KAICAICAKCgCAgCBx8CDAwzCD3UNQzUXMjIGBAmilpuHuVaYZ2lVhLB4WBkTRg0J9eDMThLv4OhQIao02nScioAWGhQ3BEi++1Gng/aFp13VGbkOZYak1yrwX5MLgOHEUVYUSg/yQco+kr1RNx+J2ZmGH3wDOiCObWrWFiHfI6TWgzfCcVEMNQSVaQXODOeh5rzNuAASG+E6aNoqKChWNgcDLa9JTphEhWcGdtLvoal9yqZkpSdk0CUj5lJmXXdoOiQg8SJgVEBjFgkK0E13FukBRhyijm+uYng+usJCgU5QYD6yQ02Ff2h+oP/g3EuUQvEO7kZioof0JGcLvXofWZEzQBnyecDiq6UJVBlQhJGQbvY05RwLVD0/uIQpKM64w1vEsehe+U+DFVFhU0JbjHfrCSFsPrUiR9MW3KOypzRtNv4GD+90vTFGHBHffR6ovBRx0zgkbcv839cTaJC3oRnHfJVTfMQ8opekSoPaulxy648vqbmW5n0tOP0Ty9xUXZAc+gb2Rge+Qpo89hWp3GyI+OIHX4kMgd9PxNJQLTIPH7sSeeNubiMccfGdkZ+jCE71vfMBUPFRZLFsz/dcRJp59FT4/olEP5Xbr1IKERmd6IhAH9CBRigkTTnY8+8zLTEd1w8TmnrsMu+haD0ciFNFI+4dQx505/f/Kr0QqIw4ePIPGpWYx+R97Od00vDhITNAm/7cEJz5GcevHJh+7+7KN3qTrbVUg28Rkrly7c5ZMS3ZW8/J1Ezzczpn1I34rI82BMwn4M4AjqpZlSDNGbIyzU5ip3/LeHooPvwOv1kCRutvTqu5OwoHfHpTACj0ybxZtJEoT7CS+LZhtrwQXbtmwOK8Vy2nXIX7VsyUJ+H3nyGWcH8OCvP/3o/VGjzxkHLq6BQfvpYy+4lNdGq5DOvei/15KsvG/8VRdTeaR0YfTYiy7nO6TKpAweItFkE69jCjgSHr2RauoP+E4oacyUNmg2nt+5a48F8+b+qDY0cEvh9TQD6gqm4GrB8OUSQUAQEAQOOAREYXHAvTLpsCAgCAgCgoAgIAgIAgcNAvy3KgPRNBgdpjLqb3CMRrXNpp84wBEjDkx5dDzq/6Fa6bVgNHs1cSlOKCm2a6xJDpfXYdJYEjxBmGtX47PaZPN2gKqCgSsG7KNLJgiO3n6v/iukkKKiwKMzBJNhXm3LaF/ug1ojQW9sYFNBMoAKCZIRi5vAlMQGyZXm/tYowDUMpjFIlAXdwnIQJ3+m5lauzO5cUpTUqsaOlE+5lkR3psHoLwJJUYBqQCWZQF8NPoMkDE1NqXwgmUAigfOBu1KLUUlI8BxJDAbSaK7Ke6jyIHHB9FokM/AMTSdrcqg8o31gHfpCFUt0uRYHGKQn0XGw+DYQS64xrrXoMgwHuDa5Rpt71yq3x8ahIUcdM5L+FD/MnPGJ2ogOO3L4cUwXxeC62vneSA2DAHYDM27mqV++6M/fmRbo6/krNzNASoLhuovOOlnZzf13EGTu++NGnX7mXHg4lJVs5xppcWEAlheDP1F8aML3Dj16xIncDU6vAlUMYNRN4mD96lXLI89zF/0a5Mo696Irrv1tzg/fRt9PNQIDvtu3bd0SeR93llO1wXvHXX7tjW+99MwTkWl+GAwmqRId7CambMcFduj1aTN/nvTBjO+Yfuq8UcMG8vktBqKJC+nxwRRf0+uMsyMvPeLokVRpaZb8+duuucDURyQhNm9cv/bBpydN/vTHP1fTVPvGS8ee/uqzTzwU/SgQC2E/JyXortYVel/w+Py5P32ncn+YjI3Ghu3S52L96pX13lHk/Y3NVYW0o39JSzDkHOzR95CBDMzP/vLTjxdCWRN9HxUIXDfr4QDekjabu0ZJzUUyQbn2pDFjz/9h1hef0jdjMzwuSATFQZ6inAcPFnfa2eMuppop0iOCapwrbrzzfr6DSL8WKluuHH/H/fQcKdq6uYBppNT6RbImfBw4TLj/dv7/9HqFc5cqDDWyhnOf6hne8CHM6Zsbt5wXBAQBQeBARUAUFgfqm5N+CwKCgCAgCAgCgoAgEPsIMAjKYDOD9WqFwXgarDIVQ8zsdkcKqMixUknA9CtUEzDgnoZUUBor7ALS80go1GrMVm2lLaXSjtiHO6V1jd5g8YXMNq/OaPEboUpgcIr4MKVKODBf13gIREU6SIuxPo8hCV4WAZ0hUKszBouBpFZv8uclZDjM1dsTzDhDIoCFW++peDmurq3GZiD7zHRQzQX189gASJVac7xnii3RvcGa7DJm5JX7rEmuSoxzA8gJqjWoiqACgztu2X/m9iYRQXPtVcQElc/k83ieZAXzh1MJwTGzzyQmGHwnhvRlKKq7l5854Wu1mgLguqjT4f7ckg36ux0VWjWPAO62JcFDlUFTqbE4tAO9cE1x7hCv8I5tlcK1yTXK+bXLWPhAH/ju9J/qgVXLlyxU86dgwJ2VQVe1ndYMPHLXP1IE1SMsGBBl6iXWocOPO2Hm59M+ePmph++N3Mm9O32MvJa59ZkKp6md9I21TRNpnvMhsq1cw6Bzz74DBtFwXMnhH3k/A8DcRU/zYcX4mefpr0ATZBI59D+4etwZYfVBZMlH1FotaKt4X7BtBvs/nPzKC5H3tYXEgO1H39t3wGGH87r7//fSm8Ty3huvvOiL6R+8E727/+9iy/sOx/uisiPaKJvB8CHDjhlZsr1oWyQB06euT5dce9MdVGS8/vyERya//OyE6BRBSp+oLCHOq5cvWdRYP5W0R2om0QOHHDmcKgj6J0Te3xntklBqjAxrbK6yjUPha8L53dI5lQf5AIP7JPqee/z+O9TG0RkyBPo3tMQPoyXva2tdCiyFsOC6pKeF4mUSqR5aBb8ZtklDbaqb3nj+qUcjn3HBFdfdRC+MiY/ec2vknL9y/J33c209eOt1l0945d1pP33z1edqfWM6LB6nUbeaqkeZ3/jPRgN1iaJWYh/3hiKoJdjJNYKAICAI/BsICGHxb6AuzxQEBAFBQBAQBAQBQUAQaAkCisEzA8pqhcfpRRAzZIXKIEnakDBQdmrGMzRvsoU0ae2CGhANoaRWQZ8t2a1NyHRswalEgymQBaWCFcF+BpqpYKAJNVUPDPo7/F5DqQsaDLQT73MbMnGtHh4YIUt80KLTBR2Z+WWW5NbV2uodCb6APzdUWxJvYropFJIBJBAaSwWldJ+BfLXgNVUO9XZmw0hbA/+MYEqb6iFQd7jwXK9WF/TotCEd+sfnsP80vR6DSkNtqkWYmojpPX5GzUAdihnQFjwLsmRpF3vdxlkmq+9iHLegLROIDz6XBAMxDO/WxXi+BWGzABh1xvhJZnBcGcadJtx5h53rKfxhkmVHMADlR/3Zxb7kox4sf0dx9FxjTa1Bzq2DyddDmeeaLDg7M3C56I959TwJlAtGn3fR5fzeWCCXgXyeX7KgPmHBFEU8zoDm808+cFe0wmBXB/7Gl5T0jDBpWYF0U7t7u5IyJzINTSb6SlPtxgLoJ40+dxzJg2+xkz7yeVQBMI1UH3h4IPi6kL4Skedpop2Kvn71yUf0SqlXOtalxCGZ897rL02MTnvEdFC8IVqFwPdFT4CHbrv+v9xZzx38u4tBc9dzPPN++r6BIonmziRGosepvOv/PXjnTdPee2OSGvEV+czO8O7YBkOGxggNXts6p10eP6MVNPQ9oCKIJJFibM7rqHiAn0if6HcU+dzG5irfYefuPfv88sPsmS3Fs2e/QwaF5/cnH75LM/doTE0ms5mpu7754pMWKTaaeyc8X1JctJWEGfg6/vdbc/KZYy8gPoqy5i/ComMnkgGc0+f/97qb+D1SfcPjo8+7+L9UA82f88Ns5dlU75wDFRRVJhXlpSUk8vie1PoGwmIQ58IrEx9/UO284t+xevnicOqqyKKYzc/6fNqHLRm3XCMICAKCwIGKwMHyD+0D9f1IvwUBQUAQEAQEAUFAEDiYEVDIiMaCSkxNtNcDTv8m4FHqCnaFZAWVA6zn8QDTQZnjQpqE9BC8K0LFloRgBQLtCMIEOiK4TswYPiZhQEUEU7gw8M+d0d8Eg9rqquJEtjXK5zJ20OqDZq/DrKktjXciDVNQbwwmIjVUIsy7Q0gt5QZ5oXNVW+GLsevPhnCwp5nC4PXOftQv9cgKEAUapHzyWBPdeihBcp1VlhDSQVlBmlj8PgOIhVArEDIlIBbcGI8f5ALVEb+RjKnDg79JNLQFAeEN+PUJ9vI4y+aFORmtu29fa4nzdsdYfEaLbzkqU0CVgKjZ7HGa80s2pieUb0npmturqG1Wp5IcEBxUCpAQwTM1fTLzg92TWwUfq9yqezqKDSOBohiIkxCKqfnXyHvlGLnWmIYruvCcQmo0Ny9i7jyD6hzUts1/5bBXBsm0SVQO8HdjefgZ3N5etLWQNRIcZH2hakjz9WdTp+xNsoJtKjvWU9J2Ehe7Uw478ugRFWWlJUp6Hd6bUZeeprH0UqPPu/BymjF/+8WnUyOfpeThp1fBVeedNjK6H1RX8Jha0JbeATxHP4IP35rUIC3OX/fu9CpQCnGlsuK7rz+fvjvjbum1VFFQiRCtrmDw+ujjTzo9AMOEpdHETN27/ujt116MJBEaeyaJhdUrGldX8D52gwFxpjqKbIcpqThnv48aP1UqVKs0lsKIbTQ2V1vnts0jaVHUSHBebRz0vODxj995/WW18/QuIblCIqul2Dd3HcmUrQWbNlB9wrZHnXH2f74AIaioazasWUV/Jo3i/3HBFdffTMLs7v/77wWRbR99wilnkLT4GOSScpwqjAeefvmtHUXbCkmGwdPlbJ4DJgXR/WKbxJuKo8h1FHldp649e5O4osIk+v6uPfr047HvG0lB1xwOcl4QEAQEgQMFgYM21+iB8oKkn4KAICAICAKCgCAgCBzECDBKzjQ+an4ChIWGv/XiyTFmuM3APzFgSiimQcrioEMIEbvtWk1VMUQIOo3RYApR0UCCgKqJclSmRKKigEFP4kNjcnpPBDUhbareEBjpcZjabF+XYd66tI2msihRU7wq21ZTkmDxOo1GkBN+v8cQgOm2IeDTo30/duC2eBYqaYSaU2FQHQLvDZdZqw/FgbTQGq3+VjDY3gylhLFyW1Jo+5osu6PCVrF1eetVWxa3WQoyohCqj81uu/lbEBRfoUdh1QkIjWqoRjY6q6zV25a36l9VnHTr1mWtg5XFie7iNZmm4tWZHRwVcV5Hpa1qw+/tMxbO6HUBrrsf5MVTG39vl7R9beafGDNVFkw9xV3nIb0xlNRhkH+tzqD5IWrkJEsYXKVvBj00Yq6orCG+U641tcK1yTV6UG6EQ9wyPAcUb4dIgK6+5e6HGNjksZVLFqkaJPc55NAhS/5s6G2RiMg678OG8BYZGO/OJNyG1DhMCUR1wu7cR4NqEgXRigfm2mc70SoHHjvmxFNHk5D4+N03JkWaX/OcktqG6bLm/dxQkaCQDvDbbuBhoNz7+dR334oOyrNtGhYzvVK0ITFxbakp9O5go1wLOwqq2TQ7wEBF3n8qfBCYRoueCMsXLZgfee6vd928WTXnU3abnLZKcL2xPsJCw+qC6XP0efqgcPyzZkyvtzu/Q+eu3XltU+02NleZAon3lu6GHwpTiJHgWr74T6b1a1AYsOfBaOLn77yTyHs2bVi7OgOSFvqM8DPS0JxqCJIEHbt060klzrjLrxtPFQ6Jhcg2SPqQ/FDSPZH8ePylyR9mt2qTe9s1F53L1FhKSi5k/6pHRLKdnn13qkvYdmPj6Yw1Q/JILcUaoOlHVYqaMmVP8ZH7BQFBQBDYnxAQwmJ/ehvSF0FAEBAEBAFBQBAQBASBSAS4e5sKARopRxcGURkkZbAkVv9Ny/HRi+EsVHpRtKO6wmQNaTLaBzU5vfw7UnKDdgTVGSRjqiQG3BkgmYxKkoLqDCoreJzKgLYI7h8GhUI6yIlEn9uoqSmN11RuS9a47GZNxZYUPZQW6e5aSxyUGFaD2WeEv0QI6gQvsi21dGZSpUC1QrPBfLQdNg2PT3Egl5NGB2KEY80DxZJhNPvzyjan6rcsbZNbWZQ0rmJrypg1c/IHrJjdtV/l1uTcYAB6i6A2Ff4aG7wu42b0OwkEhMdRZW0PT45u1TsSLyhc1qZf1fbErrVlCYcWr81si7Yy7eW209F+H9xnCQV1Gbj2wpL1GQNqSxM6YMzcuToMtRqkjyGrU6CnJSG0JIqs4VyjaSvfDUmhWJ17yvvm+LjGOF61ScC1yTV6MChNGqwBD4ykeRAx+7C3g1K4g3zMfy65QlEzbETUPfpmpknq2qtPfzWjaify/fB6Bp5buvBaeh2DsjQI7w11B3eZt+Q++g3c8cjTL5GUeOeV556KvAfZb8KppbhzPPI4iYzxdz/yFDb5V0x+eeKT0c/p2KV7Tx6b+vbrL6n1gbvsGRjetH4t1T27CtMXKWTGR5Nfe1H93m49Nq5dzRR49QpxBaR7HVPlIba4hPB/9/xgJ5Rj3H1P4/Q1K5Yupj/EiqU7ySsGuvm5O+86E4F03rMZoDT13kjWWKLmDr0rDj1i+LEzpr4/ubK8rDTy/iwwLU2129Rc5fvgvdaoNcBjVCvQjyXyWUz3xJRH8+f8OFstIM9rSXLxU42samrczZ1T0j5dd9t9jzKNW0HemgHqAAAgAElEQVTE3GJfaKzNeTn+nkf+p9NpdRPuu62BIXb3Pv0HUPlAooxjv/3BCc8PhvLoqQfvGK+sZRAeYTz5HqL7pBAWv/38varJO9cafW3UzMbDvi+dunSjCXhzY5XzgoAgIAgc6AjE+j+wD/T3I/0XBAQBQUAQEAQEAUHgYEaAQVIa+tZLaxEByCx8rxd4OZDBUkkHxcAag+NMQcQUE210eo0/LiWkScwIauLTQ7XwgKhAGJmVAQwSE1RhkKiYg8pdvtypzfQbuVAl+KBO2ATCgiSEnr4UCNwj3ZNR40cFQaCBokEDJYMBagWT12mOY3omqizQPh2+W1KY9qkps222U47qIwlClYXB4nfDQ8NuSfC4QWIkgUQIFa3OCiBlkxcqi5KqoqQglBWOmh2Jq9Gvo1b92Kn/ul86OL0uUzx++0FgGHB92qYFbd0gLr4CkcEUVjmuKqumZnuixlFpTcG4j4QXRy98JkJlEh4HSBKqMzJA2pyNsRsDXgP7TbwZZCowmDTFULM4G6FqGJgkzgeDsoBrjGtNrXBtco0eDDg0GP/mjevXMgh91LEnnKycRE6grEdfeHNKDQL13CFO0oIpkaJv7tG3/0AGb5dF7bjndUoqGEVJoNxLw+xb7n9iIo2dW7IYG7tmwv133MjUTvc99eIbZ19w+dVMWdTYtQw4v/DO9K/pKTDh/tv+j6bRkdduQ4olBmaPOu5Eqo52lTtBcDDw+thd469RMxynzwRTIH31yYcNPCrYCEkJYhitzKDCgEoDBoeVAHTkc5meiDvco/vJa/i+eI64K/dw7CRu7p3wwut7ginvZX/5yTRJ/GRfHn3+jfdnIrVXdpvctjS6po8C3+H3izaEiR72iZ/R77rfwMFDH3x60mSOV+kX7FLCyrVowiG632xTbzAY6BPCc0wDdc+Tz7/msNtrJz392P3R1zfXblNztRBpltgePRwi2+XvD2bOXXTq2f+5KPI4/S6Iy4J5c35sDG9ew7lRuqO4aE/fSeT961etDKvyaLytlo6KqoZ2IFmOO+n0M9944enHaJ4e/Xym26IPCsmKux6bOGnMuEuuYFtT3nj5WeVaTK/w/HI6asPEY2Tp3rv/AKaAY2oytbFRXcHjaumiSFYQO8UUvDFs+N+g7DoSam/iJ20JAoKAILAvERDCYl+iLc8SBAQBQUAQEAQEAUFAENgdBLgDlR4FYWPaqMKoc3h3M0os7u7mv9NJWDDgwe/9UZNhAm2wlyPn02YdfCe0Fk+tthb7WzOgCDgM57nLm9ceUffJgDrbYDqfIILz33jsZuYED8Qlu4zQKOyClMF7J7wqitdmabavzdA4K22ampJ4TXlhisZVY4ECouU5oZp4wSQC1qCSSFkU8OoLXbWWIrRsJ8lgNPscICt27FifoSvZkJEBMqUm4NclQkHRHSmq+uL7UbjPBAKlz7YVrdqu/7V99dq5+WWb/mw7r2RD+vba8vhOuCfsKbCzhLagliJdlMZTa9bCL6PMZPH541IdIEl8YbKEPhp49hIQH2tBcoTwnYGmVGBabUsOJvYZ5S02mkM/qYzpHhxjMLDezvomxn6gnlLWFtea2iTg2uQaVfMsOVDH3OJ+M1DP1DAMcN7xyP9ePPfiK657e8b3v5FYeO7x++9AXLNUp9fplV3okQ0rCoPuvfodMuuP1VtheRFOA8VSsGHdGhpGXwDT3xNOO3Ps8JEnnUZy4ZOf/lx9IoLrpcg51OJOqlzIdDwXnHbsEKoXbntowvPTvvt9BVUAg4YOO4a74pFiv0P/QUOOuOaWex6e/sMfK3v1H3jYK8889sD09996Nbo5phj6cvoH7x5xzMhRN97zyFMkU558+e2pNDWmsmLmZx9Pib6HihRsQm/39adT31fbhc7rSVgwMBx9b3vk7OGxj95+VVVdQWKFQV21e0kccAf7PU889yrNp/m+Pp49f/lDE199Z0/wjHxvJErGXX7t+HMuvPyaSR/O+I4pk1566pF7qWih6mPiGx9+zhRRj9510zW8b/ZXn00jiXHbgxOeI4ajRp8z7qX3P/vmjemz5jBwXxvhQwE+JEx80cyd7V1+w233zF64rpjvKrL/xJW/OU4aQU/+dPavfKeP3T3+GjUSQGn3/P9ef9OAwUcM433fgVAxQeLDdpqaq+WYjL/+9N2sQw4behTnEnG95Nqb7njx3ekzwY/UfP7Re29F9o0Be/5etby+v0jkNUw9pqiT9sZ7UdpYuWzRn/xeDsP5aE8VHmdqN65VphJTUwXxmtLtxUVUUH0+Z/G6M8ZeeBlTOz169853qRTFp+SxF976IJIc4/luvfoeAoP6Rr05FOLKBSlU9Ng5H3iMpumN4dJ34GGHf/Xb8oIv5y0vGHHyGVRnShEEBAFB4IBE4KDcCXNAvinptCAgCAgCgoAgIAgIAgcfAl7GEFAby0fEHZ3c/d3AmDIGoGIAmMGiZNRwGhAW+lcgmF7Url8glJgR0hnMoc4IIzPQqQQ7GQhhCh/6XjA9kx9BfDeVFLWlccf4vXoTAvNVSLPkgUm1NRJZkgZIq6SBGbcG6oWw+gIEB54Z3uOkpASKDlrzGexjSwobYvogjmcHnu+FOqIaqaDcthSnCwbZdhh8m8uRCgr9JBnAVFdKWjCmi6L6ASSERoe+WeFPMRRjb4cxVIFQqQIB4wZdk4kOrtcZAx0NpgDNuDXwxdC4HaYNcPYuNMV5ByRm2MNkDMdoMAaQiyowID7NMRvjh/ZEG9BqQnxuW71JsxkpoRZCyVJVtQ1H689CkkEkk4JQxmj/nPtui3NmtQSo/egavm+m+qm3ezqifxw31yjX6kFZnn3svtsZPD5z3KVXEgCmTfrfA3eMZ3CfwfGjjjvhZAbno3dr43fYm+fm+x575v03X36WqZMiAaSa4fm3p331yHOvhxUI3B0/7b23Xnnt2ScfZpB4T8HmDu5zjh/a75Qzz7twzH8u/u9VN9/1YHSbTJPD1DkvI+DeVBoaBuQZNB932TU3srKvT9x7y/WRu84j245D6iQGhV+d+MRDauNg6ht6O6h5W4DrsLFPMz+f9oHavelZ2VSkqQbEf54984ufvv3qc5ICrLxuxZKFf9z033FjvgNxsKeYkni4/+ZrLn3ipbc/uhUEBM3WrzzvtBEkaEgYtMY8YKqfsScecYiirKD65rnHIHm5++EJz7419Qv2gTvwn3n47luIX6TnBt/Z51Pfe4vvbNiIUafy2t/n/vjdOigDIvuOgPiiqe+89hLnJJUaDP4/fMf/XfnFx1PeVhvjNzOmfTj2kiuvv3L8HWH1BVVDTNWlqFuam6tP3HPzda98+MX3VOuwso1lMBe/64bLz482Y28P1QfnFRU+an0hYcACWBqQVXv6fmhgz7k5+aWJT/JdRbdnr6mppgn3o3feeFVjBugkIu989JmXaVL+5otPP/7ikw/drRh3K+1NeeOlZweAwBl0+JFHxycmJiljJSnJ1GlKGjW18TAVFY9XVlQ0GD+JHJKZaumilLZIHClEU/9Dhxz5zYzpH+0pbnK/ICAICAL/BgJ7ZavUv9FxeaYgIAgIAoKAICAICAKCQOwhsKiwJnJQDNgzHcadqOerjJYBpudQaWIaVlscqKbbKumguHOfu2aprLgENZ/jQ3ImTafDfct6n+gzGy2hOBAYs3BsIE71QuWua6YXYcCOgf4aj8O8MuDTDUYKqLY+j9FPE2uQASvKCtLcFVuTB/hcpnZRgfgGBtsR5xmc3t2/H4rr+sPUQQzEMChLlYWiHvkiId1e2qbH9hSoKzq4a82Oko3pHpAmx+CayDRUSsqdAI67UH+pG28iiIpSvSmgh2okPSm7Zqslwa2FyfalWqSzomoE6gynLcn1TXKb6uL4VGc7pLw6sXQT0l9VxpWZbd50XKdJz6v4qHW37Rb8TsEIid96jHv9lsWGyUUr9RcULDBc428Ykufcm4r6OwiLvW6OrDLf99mhiHXINciUYteijlbpAAOgD6NuwdpTFE/7rJ/7y4NopqwEhhk8VlIg0b/gtHPOv+S91154mn4M0f3lbnYGrhtLfZOE/DM9+vQf6AYJsmr54oVqxtZ7CwM+q0uP3n2R8SaTaZIQT95ORUB0wLmx59GToU//QYMZnKeZsloaqN3pK1MhOblFP0Jh0JL7GexmWp9tmws2qgWl2QZ3uTNrDoO//4R5MYPZVKqsXbl8SSDg9193+/2PXXDF9Td/+sHbrz965/ir1Yy/c9q1z++AlD8Qv2xbi1Ri0UHwyLGzbaZ52rZl86am0iZ17dmnHwLkWSvhm6GmOIlsk6qUTt269+LnRgh8YPdR7/8ZNzdXuQYOHTr8WHBRiRvhBUGFkNr7ysxu3YZEnlo6L+V6KpS8AGlvp4Ri+3w30WNTnsu5y/4pKdlaMt+auoZpufD666VTpFppA0gresmo3ct7uvXs059EWrTHB98B32NThAWxPXbUaWPAjaR9gvmmlo5uT8cl9wsCgoAgsC8Q2N0/OPZFn+QZgoAgIAgIAoKAICAICAIHKQJRhAV9ApgCgSlFdqkMIqCZgO9MfUFz1XDAOIYICwb0GSCmKe5IZcwgKTTZXYKVPY71bU7JCWTC0+Ib1DScPx6VO7apRGCApBTKgyA8GxbojcG2MJROBVnRGmbbpVAR/Ap/iPbwdxhEFUU0YbEXpx5z3beJam9T3TvjuBjApdfGD/CuaIV+HQ6yoEYT1BaAGemN/tOslUGzT1AvRQ3n9q4rVFpQWeMDYaFLzKot7DRkkw3ERHwwpHXay+LycLxVMKhzQWERTM2pKsC1tVBRVMGzYujWZa1TgUkQvhmZzkrr6owO5bOyO5ckm+O8ubgvD9eyfRdScE0pXq1PnfeeeZyrWsvAfWRx4sdlqF+CsGhgrroXcdznTUWsQ6bI6o46FvUmlY4wvde5qEuw9hrka9/nHZcHCgL7EQL0/3jkudfeG3T4UUezW8f0y89qTFmwH3VbuiIICAKCgCAgCPzrCEhKqH/9FUgHBAFBQBAQBAQBQUAQEAQaQYA78pmeR42s4C3MZR4fg+hx3AwU02CVQftdJeDXQhmg/dnr1Nj1Bk0ekkcMx8nfUH2oTFPEVFKsJgT/DUhy1AnkxM9QLoz0OE2WkvUZuSADzobBdOhvkhWKyqIlaotosoLjYF7uPFTFa4LB7lPRl5UgCjL0xkCmXh/chPRQf3gcJguOc4c/jcQ5DyILlTdMffUHqsto8duQ2skII28XCI/ZaKcryIteOJ4Fzwsvfuv1hoAXmBSlWnwFcSnOdQazPxHqC6YUKwdhkoX0UIXoA4kvts30U2ZaEae1C/6QkB6c4qrWkzAhkaQUki9xPAaFTE0Mp4XiGgv7BqgUrk2+m3opaRq5Vg4LAgcNAgOHHDn80edffx/Zu4rpc9C9d78BQlYcNK9fBioICAKCgCCwhwiI6fYeAii3CwKCgCAgCAgCgoAgIAj8Ywgw8E71gGrqBBzn7nsGnJkmKJYKNxVRXcId/CQtdhZooxlAz+vvn5rRIViO31QoMJjM4D+xah0BQiYUCl6dLpS6fW3msIqtKR1LN6ZrQFpovA6zBkF8GGnvNmR8D8ScqX+Ylml3C98TSQbuNmagnxVJrjRuEAVxBos/H0RCYlq7yj4ZHcraZHUsnQMigQoKpodS6y3JA6oeukFJ0r58S2qr2tL4bE1IewhSQ4Us8R4jiIoUo9XnBlnhBl4kIg6H2XY7W7Ir32T1pVqT3A58t5njvcnw0uB5kiwkSTjvtPifAmeldhOeHsD3SLKCY++BSsKIRAbJolgsfGdcY/XSw0QMlHOCWB2Uptux+MJlTHuGAFNS0XT65fc/+3b+3J++u/D0EYcz3RbTMu1Zy3K3ICAICAKCgCBw8CAgCouD513LSAUBQUAQEAQEAUFAEDgQEWCglN4MnVU6X45jNKaMJcKCG4oYMKdigrv988Jj1GrSDQjtx6UFaxMzg13dtdrFMNzupdWHg+Y9UemwQJIjsuiRZskAQ+mu8KuAybQRBtp7lBGW5Aifw0aiG2I6oOjnR78yhXSgnwULSY8OqFkwEq8FwaCFx0StJdENLYS+NdI1+a2J7q9gzg0FhnYK1BBMYXVIVKNQomjbep3GLKS8qjWafVZcH4oPaKfZUlxmWGUHQHjQGJxeICRIdqCSJFmBSqPu1fhsj0+qOIg5SYnfUalwIQFUWbNDt9Hj0qYwxRZ+R2/4IvY0pSZhEVM+FnU4c21xjXGtqRWuzcbIjEZukcOCQGwiYIuLi3/42dfePeLokaP+99CdN7332ovPkMDo0r1Xn7defOaJ2By1jEoQEAQEAUFAENj7CAhhsfcxlRYFAUFAEBAEBAFBQBAQBPYOAgwgMzBOpYFaWYyDDKBzd3c9Y8u98/h900qU4TaD6UwDxbFTWcBd/jCGxiDNIY3OoNloSwklw2zbgQD6DJxXlApUWVD5wMB5Er+HNFoDDLZr4eGQ7rGHVRV7Y0CKkoDkAzFnAJ+1ObKCz+a7+hWVhAUJgUE8iLRVGq0+2NFo9mtgiA0ViLEws0O5MzW38pB2fbduqSxKskM5MahkQ/ohzmrbTs8NVJAx4fHwt89tNFduTS6H4XYyfCu6VxUlLcjML1ua3Kq6AO0TD6onqBSYh/uygckiqDJ+MFm9CUgbxb+J2B/ix76R4GC6p36oNksismd5tRvw/VvUXX4idWDyXZUQA7xHbQymheKk4XvjWlMrXJt8EZyvUgSBgxYBkhUvvPPJzG69+vS/4ZJzTp37/TdfEYyOXbr3pNHzyqULRWFx0M4OGbggIAgIAoLA7iIghMXuIibXCwKCgCAgCAgCgoAgIAjsKwQYCGcgtBi1b9RDmYqGu+MZNOfO91gpDBBTTULlwSUcFNQHGvhVaAzGkEav12wyx4W6WhM1Nq1OuwXExXK/11AA/4bOSIXE9FF9kf4ozu/Tuyu3JS9FkD8HnxoP0kDtQSnEvcmokaQE34uimFBTXKg9bg2Hw7agaODO/HSoKdxGU8CN1E0lSVk1WqgqKszxHn9K6+pWelMgG9elp+ZWuQ2mQKqz2uryeQ1WpHLSgIjR+FwmTcAP03CoRlihIHEXr842gLTISMy0H4vfOSAnNqKXFWjnS2KK36nwxlgCwsLpcxnPAlYJMCVPQeopemv8gpqHStVKPiqMPrQ6V028320PpWq0wQwVh3KmuDoWdS1qLCoNuLa4xrjWuOaiPWO4NjkXJNXwHiwwufXAR+CeJ557tfchgwb/XwRZwVH1GzTkiBDK0oV/0GtIiiAgCAgCgoAgIAi0AAEhLFoAklwiCAgCgoAgIAgIAoKAIPCvIMB0NEw1pJaOhoFT+hcs6ZebeEATFtiVvwtc7NInCdAH9fTwQYT3qa6AmXTYvwIpoaxmm8YX8BuSqrbH5yLwHnJWWYclpDuytbqg311rqbEmuTS1ZfE1RSuy9VAXWLzwrdhdvwqdfqeMIUwGaLRV+D+5UTMg0rOBAe3m/q5YimtIWDCFEgiC0IyEDLs7q1OJD31fhv6VgnAJ2lKcbYwWXxKMtw0YO9UmRoPRn5yYVVON41sxthQoMYpAXgyyl8Ubcd8SjDkIcqIT+prBsfo8hgBwWQhcuoGcmN2qc0kR7j0W7aUgtVQA5M0InS7YunpHgrFwWevNya2rV6blVi6Bj8VsEBgpeGYB5x3a0+Na09Zl+cnmuCqoXBzz/B5n/1CwwXSLTJW1+84g/8rSavqhWFPKBcFFhTWcgVxragb3XJtco7GUlm0/fCPSpf0ZgQGDjxg28pQx57z76gtP/zx75heRfR0y7NjjN65bvdJeW1O9P49B+iYICAKCgCAgCOxPCDT3h8X+1FfpiyAgCAgCgoAgIAgIAoLAwYcAA8CNGS/skSHD/gYlUwqhTwwOM82TDdWOA/EmK8wTEA72ubWFXqd2obPaZHRVJ/cLBLS9kObJgnRIVqRNqnJU2ky1JfG+uDQnVQV6BOBD8HUIMHUSFAbb8ElD6cYKcaYHgwVqA43J5gsgyK9HKqmyYFDrhX9EU3A1+zcF2swAedId/chFP5JsSe7T41Id6VBWFOI5ZnOctxRkQZlWH2qDa0iGUIHBdEsJePsZUEEsiUt1OloZSorgbxHK7lyyDkSFAffvAEFRsXZu/jaMvQ3aHhry64K15XCxKA/1qypOPBHG40+36VFcgHZ7AM8kS5ynBxQpVhh8e4pXZ7WtKUnQb/y93WaYcWt7jVy1GceLgat3zdz8RGelrY3HYe1hSdAlWxJSl1ZvL4Cixd0zggGiJ8a2Jubo/jbN/m5/mlqDMUHS/F1g5D5BYNToc8ZRRTH55YlPRqLBNFGHDh12zNR3X39ZUBIEBAFBQBAQBASBliPQ7B8XLW9KrhQEBAFBQBAQBAQBQUAQEAT2KgJMj8St3qkqrTI9DVNsKDvAw9veI3aG79WO7KPGGBRm8Hce6u3hZ+KIOT6kMSKjkzUpNM+SoNcWr06Ld1SmJML3wYZ0UTnwa4AKI+gBKZADPwavu8aM/2OsReqkChwj8RDwuQ1bYD8dSVgwlU8rBPHpIVGGSoIkBGWChuoKBPRDMMGuQrqmAqRfMrhqzFAuUPDQbFmPK+gXwTRSTJeUyJRWIAEC8ekOvcniK68uSbChn/Ew1LbjWW6TzWuCWXYvjJV/m/RC5Xun3wTfKX0lqtHPNiAzEuKSnbUgJegxkYo0UU7014QUUsnZnUpWu6qsGLjej/NwF9ccgZGZQTy0L1qdlZcBTwxznKeVzhDM5/NAwoSSW9foc3sXabYsadPZ57ac6g1qg79P7fcp8CqBcXcG2qaZNvrC9FUhE0BFiiptT1TwFbti9DTrZj/pX3FAK30i3yxUFcpPEmgcF9eaWkoork2u0b1ikNLs7JILBIH9EIF2HTp2rqooLysr2c7/ru4qJ5x21liL1Wr7ceYXn+6H3ZYuCQKCgCAgCAgC+y0CQljst69GOiYICAKCgCAgCAgCgsBBjwADpfz3KnfaRxemp+mKugxVCaoe6ICRsOBY6xtOIDYenxbUJLUKtdKEzFXO6nibvdKGZE2aRCgMFAPqHBIN8alOk7Pakg6yQmtNcDthLP2zxehJQ5vGqNRQm3E9AvgBDYgJq8EY8MP3IhGplcKeGQGvwef36HcYzIEKt93U3WjzwS9CD6VHo1YFSlooGlzzonaoDHAvAWnSOjGr1paaU1WAZ22BomEtyIOUxAy7wWDx1SLFUxbIita4lilTeC9Nnvne+Z2R8/aoDIyX4rpSkBc8lqrXBmow/nDCrJxeRTZXjeWVbSsAUUA7EMd+R9Xj2nKoQ7qBfGBA3YpqA1lREwro4nGv3pbs0oLwSANO2fACSQHR0QqKFZIu3VDDZAmOgWmxcr5VIh0UzM5DVMAo5WN8mc0fMWq6TXz5LrjW1FJCcb7yfMyQNRHvVr4KAi1CwOVw2OPi4xP0BoMB/yXlfws1NNq+9Nqb79y0bs2qRX/Mm9uihuQiQUAQEAQEAUFAEAgjIISFTARBQBAQBAQBQUAQEAQEgf0VAWVLf2SAOLKvNOL+DJU59GOhMKjOoDCD/n8VEBZBvxYm05pad63+T53R0g8eD/EkGAJOQASVBJQLGqRV8qW0qTImZuvikPaI/hP0gQjCx6G2dGP67yAjesMnohUbhqLCakl0VRkMwWSQBnG2BHcNDK29JpvB5LGbXDC0rnTbLZtMQW8hfCVSjVZ/sc9prAJhcVwjQCt/V1BVoRQadS/X6ELr0Je2ICZ8MNL2JGTWzgOx0iMuzZEHYgXm4SFX3d8lTK3E+0ncEAO2OQCVZt+8hqoNkgiW8HUYGz6ZxioT6ZxsHQZu+aGiMOVHeFdYobL4HseZDmupx2mK374+w92+/5a1uCcV1yZDYKEFHlooMOANEipEPzqA2OiOe1gXo1I5wWdCvqKFwkNTFfD77FqdLi4q/xED+UNRqYrZjhoOVsZQoTcFU3RFm94rQ1TWZovkNzGEiwxFENiFwJzvZn5Jr4qxF195/dR3Xnspt12H/Nsf+d+L2W1y2t5+zcVjmS5K4BIEBAFBQBAQBASBliMghEXLsZIrBQFBQBAQBAQBQUAQEAT2PQJMN8Pd92qFyoF0VKYIipVAMYPz9VJged1ajaMScgODJiu9fTAnGHDAgyGYDVWEpqY0HooCnSYlp8pnS3YaoVoIkYwAQeCBIkKHIHxHEBZWqAkGQekQCob0YfsFXNMnLsldaLD6DHTVTsiuLYcKwQ8fiFZQGvg1Ib/JaPPm4LvDanJXBH06VzCoP/VvvP5eIFeWI33TAqRiqjTbvKH8Qwva4fkpIAqS8UkChYoJkhFOVAbH+TdK9G5+khMkQPi5FpWBdBI8vJfEQrzR6uua0b58I1I8FUFlkVPXjgZjaLd5YU4wvW3FDKSl2oDxDgn4DGlQUiQDi0Bau4oQyIt1Wq2lLQgO9oEG45xbSkkFaVFlMFtCBpMZ7XmB4a7pRhNxvjOSFbGoMiDGXGOReEROA67NXQ7df2N+yC2CwAGPwMfvvjlp6NEjT7zx7ocnsCoD+vTDd96Y+dnHUw74AcoABAFBQBAQBASBfYyAEBb7GHB5nCAgCAgCgoAgIAgIAoJAixFgULocVS0VDRthoJQ78jehxgJhwfEyjRJVAyWomXS0CBtu4whSOBkTMlxaZ5VvBRQPZrPNYzCY/UmJmbV++C7oYEztR8qlAEiKTQG/rrRiK+L7IS1IB30mKsQBIXsgtFOhAEVGqSXJ5YZ3RCGuKQ359UiXFEqE90UlVAgu3B+n9+t7+lzGLHt53FYoEfqBBGnxi4u40Iv72oAsoTl1JQiKOJAXh+I7g/tLUblDn4QDKBkNg/8kDByoVFjQQ4I54fl+6WnBYyQT+Ek1BsmOw+qu+QHpnzJhxl2xbWX2DihBOuE4g+1BYJgB/43UpbO6rR84evEKqCmS9EZ/jmd90w4AACAASURBVNmmyQVJk1hbGm8BqVMIsoJECIPz+RH9Zz+RFklr0RmM1UgNtUZndHUJeOpNN97H9xWLu6iJYdiLJAKTyK9cm1yjnLtSBIGDEgHk0/Ndd9FZJx9/yuhzDj1i+LFUVPz87dczvp8545ODEhAZtCAgCAgCgoAgsIcICGGxhwDK7YKAICAICAKCgCAgCAgC/xgCDBZvRt2Kyh3z0WUVDjDAf0AXeB9E9p9qEaoMGKwPqyF8UFgEER83mEOViRn+BKOlZi1UAwgga1OQBioUl+IyIy1ULUyna0EGWIMB7brCZW02wmg7PymrtshRac2DmkALEmJX0BnERMhVY3UFLPoEpFDSQ4FhT8hwWM3xXjzPmASCw8rETLgnI2g3ZwRD2mq0Wz9VVctQL0UiKHfZ5tTO8NCY365/YRnIlR51tzK1Ez0S6FGhpH0qw3dWkgA07+b73YBKAoKBcwbISeiQxOA9/E2igHhVwJNiQMfBm5Zv+K39ZozfDhJiDI4fiivswCdn9Y+d5vcauaoC5M0wRNjXuGotoarixASvy8RUUEzvlIJKA3KlhE07AIUObRm0On0XgKWBgCXSeJueI1R/kAyKRdKC74BrbVQELspXrk2u0VhUl6gMVw4JAuoIBAOBwFeffPQeq2AkCAgCgoAgIAgIAnuGgBAWe4af3C0ICAKCgCAgCAgCgoAg8M8h4EPT3LlOP4LzVR7DQDeD8H9r6/8/1+09apk72leiMkgf3ulPsgIpjjQVW/VOd22gHGmPesNToQ/Mow3uWstmkAsma6Lbo093hBCkX470RimpOZWnQ9mghdoigWQFAvPwtPjLMBvtZTorrS5oFUIgP5gGSm8w+WEaG0yEUkFjsvkMUB/UQFmRyBA8gvUM4q9B7dLC0fHdkXhAzipoOJCmKj7dfj6UFj/i92a8seNxbhAqA/wkaKi04E59khE8Rl+SjahMOUQVBc8z/RMNuUlUsD/rUDkHeA/7NQfES0pWx7Jce1m8t3htZj7GT9KDxMgWjEFTsjG9/bwpA37J61/4B5QVtTvWZ2QCn14gY4pwzVF1mEcG39kXVygUXOf3OJJhup2OikOccmFugsF8/qBKJBbJCo6Na4w4qxWuTa5Rvm8pgoAgIAgIAoKAICAICAKCwB4jIITFHkMoDQgCgoAgIAgIAoKAICAI/EMI8N+qDNozVZBaYVogBoljJVjKSDiD/Cz1UvBQaWEv0wVcNVqqLuKhEIjT6TVOEBUbQTB0gsIiFZ+Vfp2+ldHi74YUSKaq4iS3q8ZiqylJAOnxF1nBxhm8RzC/GqmQDCA5aFLt0hksbY2mAEQEIY3eEHB57GaQFeHnsdBUOXs33jOvDxt8M57vrjWvQnvJSC/VzpLg+QnExdE4QaKCBATJCe7UJ0HB77yPBAJVNVROkBRgyii2yWNUVfA6vnd6K/AaEhj8XoQ0Wdp2/Qqp7DBVbElZBAKnFuNjqqcUkDjHOSpsvVbM7kKFBkfWDZXKET7/Q1SmnKJagu0xWM/K79kAxhdCfq5gABYff3noUhETa6QZhrSrEGPixLWmVrg2uUb5vqQIAoKAICAICAKCgCAgCAgCe4yAEBZ7DKE0IAgIAoKAICAICAKCgCDwDyHAgDYDzY0pKH7GuVjyDmBgmAH8dqjVqEyBtKt4HNq0rcut2xOzNDnWJO92qCFAWgRTtfpQFdQT6W67OR1pl0hGhKqLEw0lG9I9CNAvhg/FUVBkKMSD0t56KDPyQ0GLE34PCbjO4vDpNfB30BjNfhAMFqSW0kXfw9RHNJeOJC6oeqAqRAnsN5gKjO2DHMlBWihnIKBLTGlTnYR+r8CFJCAY8P+p7n6Om+QD289Cha9GOEUT/2bhPGDhd95HYmE9KpUN/M7nU3nhB3ETgEJkC/ws4uDp0Xr7uoxi4NIbpE3HOlNtKjNIVHB+cUxUaNCUgkSIcqz+nIMjNzwsglo9TMvD8ftdYgqSGSQ4SJZwLLGmsuB4uMa41q6reweRH8SJ74a4SREEBAFBQBAQBAQBQUAQEAT2GAEhLPYYQmlAEBAEBAFBQBAQBAQBQeAfQoBGvgwu/4raL+oZDKQy1Q8L5QMHbA79P+e+u2to8LPgmLegzkftGDlmrVbvrijM7r5+nikpLsVryMwvTYGawmxNcm2DKgLpoIy2im3JQXgy6PxuowskQSlSHXUx2rxIB6XVBLwGqAN2kRDx+A5DbF3GLrFAUK9xQ4kB1UVYgfGXiGBXL4gxUzNFlsbMmKMu0yZQ7RHcnLoyI68ikJ5XziA4VQ1Keifu5GfaIQa++W65Y19RUJC4oBk3n0+iI7WutsHnIlQSFixUYfDvm2SdIeiEGXkNiJFeqJmOijhzZVGSAcRFAsaVh2sYZGe6KeJN9QCfxb6wNvgbCYoKj9/tNAa8bqTnqme4XYDrf0eNRbKCmCrSHK41vpdo8pBrk2tUTLfrJqF8CAKCgCAgCAgCgoAgIAjsGQJCWOwZfnK3ICAICAKCgCAgCAgCgsA/hwAjwwxcc5e9WhmJgwzuc6d9rBSFpPkOAxqM2iE8MEgkdHrj8IBPm169I84bDBo7mOM9geRW1SYYRnsNRn85PBmyi1ZmO0A4mEA4kFjoAU+HYGpOFe4NapCOaRtSM+kDPoMeZtqrcE0Sgve8btfueBwrh78F1QJqRTGj5nuhKoGkQwXqIc2BHyY/glo/VCBVK77rvLbb8HWLk7NrWhmtvuNBjWSENNpVUEYsqRsvFQtM/cTUUHwWiQoqKVipviA5oCg6SGSwD+wzCQiqL1xoqy/UIt2SsmuTbEnuMkelbW5tWZwFqpK28OWgikXxnSDJQb8QkiCdUam4iC5OsjfwrjDvTAXVQPBDHGi4vcvYojk8DrDzVPpwrakVrk2u0XoszgE2PumuICAICAKCgCAgCAgCgsB+hIAQFvvRy5CuCAKCgCAgCAgCgoAgIAjUQ4C7uxmgZqqe6MLgMIOkpagHrLoielBQWwShsiAJwx3tVBPsJCw4SPon+L0d/G6NG6bSKfCeqEAgfpPJ4nMjjO6s3JqcCUKgFdQUevIbIClCiRl2b1bH0hoE7wNIiWSH6bQD3g4hV7VlffWOxI0gEbYhBt8WRAWVEiQKWuIHwr8hWEl2UP3QooJnmLFHX4sUVdnrf22/LrtLiT85u3pVQoadJuIdEO53wTvDB4NupT32hV4VJEdIStCUm/3kO++KylRUDlSSFiQslHlCEoLHjWjPoIsPwpVD4wBRYYSx+Gr6eaAvJBmWotL8+0hUzieSHdFsBMkNB26wB/y+TBIX4fRaf42Y6gw+l32JtXRQHCXXFvHmWlNLzcaxc40ScymCgCAgCAgCgoAgIAgIAoLAHiMghMUeQygNCAKCgCAgCAgCgoAgIAj8QwgwSMpd/fQ2UCvKrvZd5xYV1mj65bYwS9E/1Om90KySXqcwsi2tDvyNVhsH4iIuCGTcNdbUsDE2FQdaTQGUEUYE4ut5CUBpUGtLdhWAvHAjZZQxo315ld4U2IGgfQieEqVIGzXFXmGz1uxISEeKqMvQVr00VM2MhX4TSlmAL/SFiE4ZFd3EKPRxsLPKumHzopzVVdmJW+A3UZmYUds14Ndvh3/GOluSawG8J36zpTiH4GYSN/SzYLsMijP90GbUHqgMljMd00l1D2FwnZ4aVATwepIWlcDAbDT7XGltK4vs5TYncEgGViSChqMy2M6/iUiO1Hcm39ko1Cohjd/rLvG5nR2iDLd5nnOU78ADsikmCAuuoahCooJrTa1wbXKNisKiEYDksCAgCAgCgoAgIAgIAoLA7iEghMXu4SVXCwKCgCAgCAgCgoAgIAjsOwQYuGewVC2QzF5wl31j5/ZdL/f+kxj4ZnCe/gw7SzglUUAT8LnhQ+GnosDG7EShgE4xpK7373peDqVCDcgJj8EYyEDqpXiTzVuL4L0LfhcMMpclt66OgxpDC7VFzeqfOhng8fAdzbdxTgni88k0/6Z6gMcb+9uBwf4BLYSBKoYskBY2kCXxVduSt6FPmZWFySRKTMGgdq3Z5q1u23dbN6PVazGYA26cZx+Ysokpn5JQ2xIRVLaVH9EvzoVwSihUpnbiuR2oW5Aay5Z/2KaytXPy59aWJpDMIKnBcVG9oShGVM3doagwG0yWoN5oLPB7nHk700KFSxkqTciZoopKjFgtxJVrTa3wHHETD4tYffsyLkFAEBAEBAFBQBAQBPYxAkJY7GPA5XGCgCAgCAgCgoAgIAgIAi1GgJFhBkRpztxL5S4eV0iNFjd6AFxIpQBJCY7/G9QR7DMJC7/Xo0HQ3GYwmqGUMDM4rygaGDSmuoKBc/4bH5YXASoqQiAqUkBeMN0Tg/1UJzDQvgZEQKJWH+oLBcbyniNWF+xYn/7Whvl5s0AkDMX5U+ra+w2fZ9S1qQYdiRU+l31prjCwz536JESY6skCL42L8BkAgRFvSXTnJqU5HDDLToYiJKOmNMFlTXD/Yk1yV6Cv9EkgccG+dOL46h5G4oFYKYW/eY5EBCvnyBcgHXwGE1zGXab1IEXy6vobqQxQJStwHagfQu9PCPi8eUE/uJm/CAtizfRdfE/EPBaD9goZQRzVCo8T75hQlzQyRjksCAgCgoAgIAgIAoKAILAPEYjFHWn7ED55lCAgCAgCgoAgIAgIAoLAP4gAA/cMVHMXu1pZg4MMwqt5D/yD3fpnm6aPBZ7AgP5C1NdQw/4AMH0OV7/bhZh5kGmIItMvEQdFjcLgsRtpkCoQWy9FgJ7+DyxUFAxEpZqBbfL6BJAZh5vjPGfk9irq2Xnohiq9IcigPxUKDOj3RG3KI4Smyy39m4IpnFbXtUe1BBUQNNduiz56LHGeYEK6vZPXaRxQvDqrfenGtE4VW1O6BQNaH8LhnANzUUlCKM/jGOhrwTRRBaicKyz0lViLSp8Kjrk3iBEN2rM7qqxML8V+cM4k1I2z7rYGHyQkXMDa4XHWtvW57FC31OMkSPzwuTR9b4n3R2PP2V+PK74enFtca2qF74W4x4yPzP76MqRfgoAgIAgIAoKAICAIHCwIiMLiYHnTMk5BQBAQBAQBQUAQEAQOPAQYBGVQmv4I7VGHRQ2BygPuumfAmoHsWCr0BNiESsKA6ZjCJRTwaXweJ1QWLp3B3MDvmgF6BvPNIB12pLWr1CVn10BqEVL+zc+gOtUI6XVYKt4QbKgKxIU9s0O5cfOi3CpnpdUH1QPP81qlMFpPAoCFbSmqCkVpwFRNzZlwkwThu+J1SltaEBLGmpKEKp/XkARjbL+71qIDnWJEyqs+iRlxW+LT7V6Mg/coxMBGfCdGfVE/QJ2Bej4qCRQSMvSvYKXBdmu0V1y4vLUH6pHjcIgqE5IaJBwYjCfBo6awoHLEB3VFmddRnQDT7bpLFTjChA6VK8QhVhUGHCNJrrDKJ6r8iN9cm1yjQlioACSHBAFBQBAQBAQBQUAQEAR2H4GW7oba/ZblDkFAEBAEBAFBQBAQBAQBQWDPEGAQmEFn7qx/B5Um1ErA2o7vVCCwKoHv8NNUTIP3rBf/wt11KgumT2LKnZVKF0KIq2v14B+Q4yjCS0E5TcIgE+mUvCk5VTsyO5SVmeM9VUinpBAW3AlPDPmbQX0SEsSYKgUG+vtClXF8p8M3btUZg9PwmymclEK8SQ4xBRJ9ISJTQFGNwd/FqE2lReJzaXZNskAJ8POTKaEMfq8+rrY03oaaCFVFmb0srhy+GmaoI9phuP1wHU2y+a6pPiGRwtRQDKiz7wyo0y2afSb5QBKlGu1uc9eaq8sKUtvB6Ds54NMz1dV1qPykwqLJAoydAZ+vzO9xJ0SkglLuIWFCkihmyDKVtUO8lXXGOcDCNch5xDXJtemA0X2sEjbNTRE5LwgIAoKAICAICAKCgCCwlxEQwmIvAyrNCQKCgCAgCAgCgoAgIAjsNQQYeGZlcP081FxUJVDOtD43oFJ5wZ3wsVgYdGdqozmoO4PFoaAm6PNqmJ4oFGC8vEExgLDw6A2BYp0hOBOqBKbyYdoeBpkZfGaQn8QBA/uRhtE87wHatSmtq4zxKc5S/KYCQSn8u4EKB8XkO/LBVIDQyJvG2CQNGtttz6A2SYI8VBIbDPTz/bJffpALBTD9hnrEqPHYLTkehynV5zbGu2otnfCpB9nwK65jv0ic8F4SF9zdT0NoEhdMkcVPzoc0VCNoET2UIz57eZwV95P0UJQU7CsxpeKkMf+KYCjoX+uo3KEP+lU9tb/DvSvYHxBMsRqwJ5ZcY1xrXHMsXINci1yTXJtaEB2NYVh3i3wIAoKAICAICAKCgCAgCAgCLUNACIuW4SRXCQKCgCAgCAgCgoAgIAjsewQYBGZUnoHlSL+GyJ4wmKr4N+z7Hv6DT6xTWTBA/xPqdD6Kqgqab/vcTk2gfhCdJAEVGSAhtGutSa4yBPzXuqot83BMSd/UCt8Z0Gf0nWTEfNQlqAxAK0bfDr0xmNW279YSk9W3huQHAv5IKxXmIKjQ4N8PJCWiC0kHpkdqytOCQW2qMVhIfESmp+UDSDJsxBCr6GsNAgMZsHTeysKURKgjkJJJp3hgMFUWVSfsewGqovwgocL2qRghmVEQDOiWggSpAWHhBmExKKrT9OpYhRr2CFEppT6X83efs7b7Xz7bu676BN9oiE4sY9G/ggPl++La4hpTK1yTXJt+UVg0gpAcFgQEAUFAEBAEBAFBQBDYbQTEw2K3IZMbBAFBQBAQBAQBQUAQEAT2IQLcSc/gNNPSHKryXKYJYgCdqZN2BdKZ2gZB1H3Yzb37qEOG/kdpkIQN/RqYRom1DQmLAFQWQXgqUG2h1evtSBG1VavVUbUQj8B+YvX2RD18G46MT3Nszksp9CMtFLFhei0G9HndctQC1M6oDDozzRNJDCuu1WV1LM0zmP0rYH7NgHWG12XcZi+LX4C28wN+fSqUCyP3YMQkX85EjUzlRSKE6oulqBXow0kgSmxQiZRrdKEtelMAmbCCmThHtQlTX3EMrCQnOC4qPEh6cCysJCECaIP9J6lADF2oy1DpC0LiRiEaiCuJlnol6PfPdturcsAQgdhoIKAgIcI22GZMFJV0UCSIjkXlGlMrXJNcmzGTEismXqQMQhAQBAQBQUAQEAQEgQMcASEsDvAXKN0XBAQBQUAQEAQEAUEgxhFgEJrpiz5DvVJlrAzEc+f8bNTVqLFm/stIOckEGov/hjp6l8rC5UAsHeoHg0Gn1WqXGCxxFnzGIbbudFTEtdPpQmmoqVAYFGj1yCW1U3VA3woG+qkuYJCf2P6ISjKACgkSBwz056e1rbCltK62Q5kQRE1wO0zJVUVJH25d3nqIx24aCQXE3516J+FGhQFgnxgY528yTMeArCjG80Px6Y6waTjIkxJLgjsLx9PwTA8+SUaw7wyUk7CgMoNpoUiA0FOBRALH2YrtoOVC3MfURiQXOG6eZ6GyhIbSkX4cu8YEBUsCUkFhnKrDJLHyM2pVjKaD4jzIQeXaUlPUEBSuSc6fWFtzqi9cDgoCgoAgIAgIAoKAICAI7BsEhLDYNzjLUwQBQUAQEAQEAUFAEBAEWoCAiioihJ3fDLAzNdK9qPdHNEP/gdNQueueQWgGnmNitzeC4MowQ1BbMOXRn6gMIo9WTngcNUgL5dPEp7eyhYLBEcihVA6lRUcE58t9HsMKeD9oTDZvHn5TOUEMmRKKZtUM2jOgT+Nkqg/G1LXJ4D+vIYFggNF1UG8M6FHBjGj8lkT3UFuS65ek7Jrfl3zZ4xW/13AJriNJwID17qaa5ftkSiGmceK9yv0gFrTtNNpQtcnq9UHlkeystvrjUp01SFBkAe2i1+rDqaRIIzBFFT0U6KHBd0/Cg3OCeJFN2eJzGxZWFSe1gtpkAH6rKSlUyQqQQl6tTtcLShZzKMz11Csf4NcsVGIaq+mgiAvXFNUsR9ThqhA9BINrke8wIOmgoqeH/BYEBAFBQBAQBAQBQUAQ2BMEdvcPiz15ltwrCAgCgoAgIAgIAoKAICAI/B0EGBimeuI5VO5sV4oSQGWaH16jmHSHz6ukuPk7z94f7iEJw13u2agV7FAQhtv0sKDxdiDg0xjM1hQE2Bm8Z0mBqkKHQH/J/7d35kGWnWd9vr1O9+yrpLG20WZJtmVLluRV3g1eMQSCY8CkEgiBImvxT6qSwB+pClSSKsKSUAQTKEIIBoKDDTbgBcuWV0m2JEuWZK2jkUaafXqmt9t9l87vaZ0zunPn9qy93n6+qrfOveee5TvP931V3e/vvO/7wmMX3Xls34YHUsuBWg2kRcL7TlooohIQLW6MUYj76hhRCDBF1MD5z5ZjNoTsmkQ2bFyzbvo9STO1Yf22iafyHQGAlFXn+j8Fx/NMiCUID6RwaoljmJkYWFNvDG+sjvYP1mtJQ3Xp1MTgcJ6p3tM76zwnuoJokFfGri/6WaaIIiIAAeP5XPGb9an+dUlnFVy9RFcciN0fezL2RGzOlrRb1dSuGG/WOupf3GtX0eeuiC5oWyvlOuI5WVu0VrGCNchaZE1yjE0CEpCABCQgAQlIQALzRuBc/7mYtxt7IQlIQAISkIAEJCABCZwDAd7kJ20RUQDtDec1dQxwVJ93nqJz6MuiHlqkHCJKgnbCcYxoUZuerDSn85L/yXmL+Bt/kFRIR57dsu6xr1zTVx1bg1iB8xnhA0YIBIgRt8SIcuA70QIvKzjiiEbAoJXpoxAnXp00U+8a3jhZy1XmShV0Jj6ME2II9SW4B2/zExlBQ8QYGRiq7R3aMHUsosXg+i0T16To9zZqa8Quz++IBLtjvOFP4zluLq7Jc3C9HTOVnldMja/Zs/+JHfvydKW4wfMR2dH5/6CZmaSPan4vkRUjEyOHepvNU/QI5hnFzRE8SE3VOWHUmQgs79+ZH4wRz8raam+sQdZiaw2S5f1E9k4CEpCABCQgAQlIYMUQULBYMUNlRyUgAQlIQAISkMCqJYCjHKf6R2IUZm5vP54dPxsjwqBbU57iyOfN9ntjOMxfbHGXT0+OxUYr9enqoaQyIk0Szn/EhO9LVMI7psYHD9eqA2NJDUWdh0uLM+FIFEUpSuB8RkQo+XXivDbX+EIiFuLMH16Te+/O8YQg4NU/V8c9wkvp8CbiAxGBNph7vCypnHpi/K+ypnegsT4RFz0RSHCgcxxv9tPPa2JEivCZCArqfPxBjLoYk3n2I+NH1vak/sbrBodrgxE77sx+ikRz3a3F/Vo3481mY7QxPTU2fmT/FfWpyVe0HcP9fy322djuGPOyGxs8WUusKdZWe2NusBZZk93KoBvH1WeSgAQkIAEJSEACK4KAgsWKGCY7KQEJSEACEpCABFY1ARziOOn3xSg83anh/D7lzfkuSguFY/ie2B/HHojNvvqf1EWVvv7+Sv/gcGxoe4puE0GAGPDuGOmeahErPrjnvktvSnqkPQU/OLY3/i8oxQx+65TqaGtkiV357bq+wcZQhIXP5TMFwec9LVCtOviqI89tGZqejH7R7K02Gz2NCBBEZOAsf1OM1E84zHmm/xf7TIyIByJGqLvAsa/ffOmxn9tx9eGXb7vyyPia9dMIOaTV4lk59qQIkdQBOTg9MfrQyN4nL5saHUnQyikIvppzqI/xdAyB5lxFmg7Yl+Uu+LCW5oqgYA0yh1iTXZESa1mOgp2SgAQkIAEJSEACq5SAgsUqHXgfWwISkIAEJCABCawwArzJ/+0YNQg6tVdlJ47zsojzCnu8M3aXND28+U76I2pO9JIGirRQiQSYjbJITYtOzuOdcavfVpsaeHvqOPRHZEDsIAqBSA2c9mUjBdCWGJEKtE7/J6xNlMPb89vOtZsnN/UPNqingdO+NcKi/Mx+6mbg3CYVFfUuykakwmlbBIoXEh1x36HdWydHD60bPH5gw3jqcJDWCgY40xlr+v+lGJEV3IvUVbfGiLzIs1bWp3D3th27Du9ds7b2hdTDIMqCFEfMJepZnCTcNBu1teNH97+mXpu6eGbmFA0GwejXY9S/2B0j4qUrWpuox7izhgDAmurUWIOsxa4ocN8Vg+hDSEACEpCABCQggS4ioGDRRYPpo0hAAhKQgAQkIIEuJkB9hWcLZypvubc3nNSkr8FhTQ2DbmsIADjovxIjquBEm5pIOqjqRGwSEaPdiXxZRIpNx/dv2JjUUIea9d7RfEesoP4DAkV7O20NkEQ5HM81HkptjL4IID+dk0mthABB4WzGCEc+1/5u0U+EkPtiCBZl39h3pjfzd+Y+bzr6/Ka1I3s3D6VuxiURIIiaoH+82Y9AgXBBRMV7Y3fE+N+Gex+OjLKjWe/rzcGDA8O1bX0D9eH+NfWd67ZNfCmFw++KcHFVjns5D59IipFmvfb01NjxF5q12vVt9UBKPn9aPA9RLt1au4JnZe2whlhLrKn2xtpD0GAtMt42CUhAAhKQgAQkIAEJzCsBBYt5xenFJCABCUhAAhKQgAQWiAAObpzRfxL7ubZ7ULfhb2I4yynKzFv4XVV8O4W3eX4c/t+L3dX6/HG2V6pjJ4IlqAdxSqvX+jZFZBhKlEJSIs1QoJp0Ua2NyAEaYkLHFrHi2cnjQ7sf+twNl0weG/pAvlMTgzoYpGmib6QQgj1bxoTUVIgM74zxtn7ZN/4HIb0Sb/EjPlBzgjYSOxH1EGFlS9JYVY48t7mSKAvucXH6T1onnOpcG8Hlshh1LLg/hbARRnpTcHtrCnXfkOfeGLFmS4pv37B+2/glibZ43bYrjrxlcO10oi1evOlMvT5VHT363NT48VcX/WjfECGCc577kUbqTGLLHJdZ9rvLKB7WEGuJNcU4tjbWHmuQtditHJb9QNlBCUhAAhKQgAQk0M0EurUoYTePmc8mAQlIQAISkIAEVjMBHMZfiOFALiMpqNvAW+HPFL9169+4czqI43KvTI2PVHr7+ir9Q+umUsviJOEi4sKag09tz6jJmAAAIABJREFUv+aSlx9o9PU3pnr6m78bVj8Qe30xmXaeZlIdj3jwpwee2v5E7M3V8TXvy7GIEognFOpmHEjHREOMQKQg+oF0UDi2SWNF36mRwXk4xnH+H45dFCtFEtI1IUiUjd+3pch3Ze/DOzdFrLguosPD2644ur5voEEdCwqGE9lBeiesJ/3ckMiM4/Xp/umJo8PrI3SkDnnvgaENUxvr030pwN27PeceHtpQfbA6WklKq4H3pDcb+voHbukbGOipT51SloIdpNG6M0ZUB/frZkc9a+dQMVZXZsvaKhtrjrV3Uu2Plt/9KAEJSEACEpCABCQggQsmYITFBSP0AhKQgAQkIAEJSEACi0QA5zGOeJzkpOhpbbfnyxtjOLxxvnedaFFEWSAAfCxG8e2T0j8lpVEiLUYqU2PHnk8x7q/n94dbAA2Ojwx/fyIkNsdBf1v2vyfWWlcCIaFVLChPxUn9fCIdDu59+JJtR/ZsWZPP1MJAdCDCohNn9r05RsoonN5EYZA6Ckc396T2BWmFOjm+iZwg3RA1I4icmG3pd2Xf4xdtjmCyM5+5PmIFjYiM3+C66dPxxnTfTK3af+zY/g3Pjh9d2xxcV1vb09vcMjBUu3J40+S23r6ZvX39tXvWbjrw/MzM9IFEp+ypVSfWVsePrc92tiZIW8NBf2fsazEiQOa9wHj7DZfwO1xZO8wD1hJrqrWx5lh7rMFuLTi+hPi9tQQkIAEJSEACEpAABLruHzmHVQISkIAEJCABCUigawnwZjvOVJzdnVIX8SY/aYF4KYe/c7sxxz6penbHfiVGgey3xWZrDTRqU5Xq8aOUYLhqYGj4hd6e3r5EWpyYDDON3h1x4m/ZvPM46ZVwTJNOqaw78Wg+44RGzCgb9RoifvRMpP7FxggV30u0Q+sb92eaaERMUCeCTjBmCCzch2gMxhHnP9dDpCgbb/d/K8b4vis2G0WTPlQmjw1X1m2ZWJti3GtS9PuZpHziOjD4wIvHzWxu1PrGq2NDh1Pz4rKNl4xuq1f7BydGhoeH1k/VE50x0j9Ya9YmZzamnsXWofVDjx18ut5o1GqVxvRU7tGInRQ8QaoqUlY9Hdtf9PdMz7ySf2fNlKm1WEvtjTFhHBm7bo4yWcljaN8lIAEJSEACEpDAiidghMWKH0IfQAISkIAEJCABCawqAjhKcYB3etMdhysO8isKx2pX1bFglBNlwXPjMH4sRpRFWXtidhI0atOVWnWs0mw2r41YQS2Cso1FyKgcP7Dh9REehhKNQLqlMp1TmcYJcQDBh/RKRC5UiVqoVQdqKbB9NGmWKKTdqVD3XBOQsSI11PoYERxEWVwX435EWfAsZQF1ohc4HjGFWhJEX3wxdiKKpNnoqRzdu+mbB3dvuyfCyaciYiBsMMZvi9RyVYps70/0xY7YjZOja7ZWj69pTE8MzGzcPtabwtvPNOozu+vVqUZ1dGpoenxq6+Sxgx+cGjty2/T48UqjPt0eXUEkCFEVfx7jPqSCOqVlPOZ69pW2vxSVWDusoU4vtjFeHKdYsdJG1/5KQAISkIAEJCCBFURAwWIFDZZdlYAEJCABCUhAAhKYJYCz/fdjX+7A4x3Zd1PsqhhO8q5rhWiB05i3/suC1cVzzlTqSW1UPXZ4IOIFNT3KHEeIBolSGBqcODa8JXUe+D+gTAHFW/NEW1BjguMptPxsBIHH9j+24+tPfH3XoYe/cD01ISi2/P5zAMo9Wv/fwNmNQxzHN4II44NQgWhBpAf35rkQNqiDcW/st1rvF/HkQwef3nb9sw9ceiT1Ke6JUEHESS3CymBSQV0cIWNLttsTjTE0emg91+6bHFsz/vS9lz36wqObxo4fbGwcP1K/beSFnlumxuqX9/UXvnfUnJfa/fn4q7Hfjv1tDLGCPndzGiTGgjXD2mENtTfWGmuOtWeTgAQkIAEJSEACEpDAghEwJdSCofXCEpCABCQgAQlIQAILQACnMU5THPWdnKeXZD9vxxMJ0M0v5+DcJ7rif8beEqN49WwjrVF19OiWnr6+xrotF4/09PZuJzNUik2PDW+s1pM2ac3YkbV7Nl08ipO6TP1Duh9qE8D1LyIA7KqODu156t4rNyRi4cqZRs9PZh8RGefSGKtOUS6IDNTQQJhAVCFNFM5yIjwQBng2UlYRnVGKGCfGMv2/IWLEL77sxn0U/Sbt1GT0hudG9m364r7HLnrz9PjgdYnGmEm9itHaZH+10tsYaEw3X5V6FVuqozPXjR7srYwd7kkkSk+iKk50j9RPpKP6UoyojqdiRFYwxzpGFHRRdAVjCl/WDGPGGmpvrWuum4Wbc5nfHisBCUhAAhKQgAQksAAEFCwWAKqXlIAEJCABCUhAAhKYPwK3XL6xct+zJ9VnxuGNKNEWXTB7z38ce1WMdEnUYODN/W51sPJsD8TujH24lXgzKY6mx0a29w8OPbNm/ebhnt7KxIYdY1+LYPGaweGkjZrqvy/H72obJbz3OK4fSjTF17931zXrq8eH/mlqX7zt5ACEsx7buVJykXKICAoaYgCOcraMK9EetKtjiCkPxR6Mvaa8K+JL/2C9NwLKxbHpnp5UAO+pXN0/UH988yXHt+9/fMex0cNrJ3p761unqxuj10yvmRytX3rgib5L+wd6K5OJl2hMI1bkpi8lFkOw+cOC53PZPhJjftUjTHTr/DmBtOBOdMWPxdqLbXMcLFhzjJFNAhKQgAQkIAEJSEACC0agm986WzBoXlgCEpCABCQgAQlIYMkI4DzGUc/b8BQQ+OUOPcHhSiFn3tDvujoWPG/hRCf6gHRKn4gRbXCizURhqFUnK+OHXriyOnb07sb05GcTebEngsV3hjdNHtnysmMwwgFdNgQD6lfsiQiwIZEKEyMvbLo9tStuPk+x4nQTpBQrOOYVMaIrGKcyfRWiBeNHxAWFtU9K7UV/picHK4n8OBT7XH4f6kmR7a2Xjfz41suOrOvtnzhSn5pYN350dOj4/pnUvaitHzt07NKJo1Op4ZHi3SO9lepYz+T0ZE+iUU50k3RXfxcjwgIOpJPqZrGrdXxgz1qBeSexgjXGWmPNrRYmp5u//iYBCUhAAhKQgAQksIAEFCwWEK6XloAEJCABCUhAAhJYEAKIFhgO7W1z3AFHPo7vrqxjwTMXogWpjL4Q+xex32xlMRNvfG16sjK675k1owd2Hx5a//zR7bsOHUlqqEYc/KSQ4tyDsfKt+S0RAw5XR9cMH31+U73Z6D2a33BQ8zuOfNz7pErqFNlyIQNdjuOzuUgZ88D/KdTdINLiZS19jMjQk+LivYdTPLx/amLwovS5ETvGhOgbqA8NrT82UZscn2pMVS+aOHb0YoSL8cMTlanxRqU63lNJ8EmlWa8Mt4gVX82p1PNgvvCMFARfTYWlWSM8e1kAvX0sWWOMUbnuLmSsPVcCEpCABCQgAQlIQAKnJaBg4QSRgAQkIAEJSEACEliJBHgrnOLQvxfjjfj29trsuDFGXYaubUUBboSFr8eIEDi5xZPfbDTeNDUx+RMHn5pYO3po5qk46r+bgygkjQOa8xAt4DmRYtWfffyrVx87vn/DNREGiG7AcT8Ye1uM/x0QEDYsAFBS1d4QaxWYuC+iBW/+n8gJlhRQiR4Z2NZs9lySJ7gsNS3+OjU2Pl2fnnmyt6/27aEN048kouTGZrOxjQLkRJo0avXKbKTIqcmd/k32/lKMWiDUrECsKCM9FuAxl+UlWSOsFdZMe2NtscZYa6dEK5GuzSYBCUhAAhKQgAQkIIH5JKBgMZ80vZYEJCABCUhAAhKQwGIQwO3MW//7YjjfP93hpryp/3TspSoFi9GzJbhHIVpM5tY4l/+gUxdmGjPbDjzR+7MPf37g4NRYz76IFmNx3vPWPAWm4XR3UkE9cHjP1u+MH13bSHTF+7LvltiJYt4drouIsH+BH5nxI8oDQYMIgIPpZ1I6rRk9tm/9I/1rputJdXVxpWfm0tSxWFebqmx+4mvNn6xVpy6anhit1CNWNGucPvucrY2IkS/GHo99o7AXskWs6PaaFe1Ddrq1wtpijbHWWHOrjc0CT28vLwEJSEACEpCABCTQTsCi284JCUhAAhKQgAQkIIFlT6BD4W0cy6QmIpUNEQbtjVe/2T+Ygt3VnN+1jtZb7/goz47TGef7n8W2xz7QCoToglq1Z8Oe+/t/LGLF+uvfWj8+vGlmsm9g5nBff+XhFOW+uNkkBVR9AymhIgqQhoni5e2N+5TFsYl+uJAIFq5DREVrsW3GqXyTn+gO1IZSeNoYceJofh1sTNX2P313z8j44eEnr33j9L5atdIcO9KzJc/3xpEXprbUp3PJk4tvlP0kmuQ/x0g/RU0GmCFmdL2w1WEsKWYPayJZWCudwiXYzxqbLUDeeg2jKzoRdZ8EJCABCUhAAhKQwIUSULC4UIKeLwEJSEACEpCABCSwFATK4tvX5+a7OnTgw9l3b4y36B+OUaOg2xuOd+ox8Df+k7F/2frA+O9Tu+Gtzz3YXzm0u6+yYUfzExEqHho71DN90TXNmRTY7p8an242arUDPX39FJ2eK/UTDm4c/IgNFyJYcB3Gkahvrse2VbDg+1CzUSd9VU9Pb9/2Rq16qD49lUiLnunqaPX6x7/W3PjMfUNrZ5ozr6QmRTPWmI0DOEWfeix7f61gQ4Hyu2McWU2EymqqV9G+BhAjrou9I8aaaW+7suOK2EPF2HQ4xF0SkIAEJCABCUhAAhKYPwIKFvPH0itJQAISkIAEJCABCSweATzSvPHNm/JzOZxxwPL7gbxJvjdvhK+Gt+hJ0/Tl2O7YpbEfaR0S/PgUnR4/0hPr++H8dnv2HR091Ls/UsHmvsGeyzbtnBke6Kt8f4ehRDhARKCmxEmXLcagFBz25vtQDEFi0xmmBG/4t4oejCnjhD03MzOztj5dHW6mevjA8LqHI1Zsnx4f7alVxwdTo+LqZr1xdXW2usVL5RVO1SpmBStqMNAvtkRZELmxqsWKrAkEJ6Jxro11EisAy9piDa3GVFlnmLr+LAEJSEACEpCABCSwEAQULBaCqteUgAQkIAEJSEACElgMAjhTqd1wX4yiyT/ddlOc0t+Ose2Lg7bZzamhimeHCbUeHolRUBrh4KT0UBzX4tS/PF8vJzqB1mw0704tiKT/SczCTApdz8xM9PT2Inzk48xIZIHRxDrcmC8j2RLRsY2fYkQrzBbuznH39/T0bM4xO/PDZD7zFj+iRPoyk0iHHu5J/YxO/4sM5Lxarl1L+qfHG/XpkanRkTdFoLiyMnLosUZt6uUJAUnv6DC3O2Omr0/mIFJKEVVxf4yi2tVYI5EVZzy5YNp1myIVFIJF6xppf07WFMxYY6s5CqXrxt8HkoAEJCABCUhAAsuZgILFch4d+yYBCUhAAhKQgAQkcCYCvIn/QIy36NsFi6uzj6gA8vD3rgKxomRV1n7gzXjqNVCrgaiIHz0TzGa99s9Gnn+6snbz9vrA0LqZvsGhrXFVJ5ihVo0QsTVCwYH+waGJmWajv1GvjfYNDE719vYN5YDp5GxKAe6Zvma9flltamI/xzbr08+tWb8l2Zz6BtAXmo3GsxEwjkYEuaKnp29DttTBOKlxs4gWzerokTdNHj+yKdfLeYgUMxnPVo3hFL3h0Vzohhh1KUiNRftU7KnYgdjhWG01CxUlaNZCRAsiYlgbKD+slfb2f+AVWw2RSWdaGv4uAQlIQAISkIAEJLBIBBQsFgm0t5GABCQgAQlIQAISWBACOFMRJV7f4eoXZ99/i/1G7Ntx0E6tItGijHq4J89OOp8tsa/HfvVMo9CYrlaqx49GkKhvHViTwImEXExPjK3t6e2pNGrTrx3euK0SoYGiEtON6alKs6+vLymbhnsHBusphHF0YuTQVdMTx6+NYLEvB10a0WFvb//AJyM47G3Wp26NCHLx8MatPf2Dw1P9Q2vXRsDAcY5GMRv6kYiKtRE8KtXRoxEpMrzZF7GEMT5F3Gh5FqImeNY7Y0R98MxEV3wjxm+rPqqiddxbim2/NvupdcJaaW8vz45vxhQszrRo/F0CEpCABCQgAQlIYN4IvJTsdd4u6YUkIAEJSEACEpCABCSwMATiaG2/MM5uHNmvjv3b2PvaDuCteoot47j+UgQL3hhfVe3WOz5a1pLYlQenNsUdsfeeFkJEiggJiBKVRFGkWHeyNEWkaCYVU//AmkrEiRN5pXr7+gnBmBUXUm/icLNWi2AQkYEbdCgowXX6uEZvX2Vo07ZKhIsc1ogoQiaq2ZNmP9enqi9epcM1WvqOMEEUBUXGmQufjpGqinEm6obPqzr9U6dxzjoiJdfbYm+I/esYIk9r++t8+eXYd2KIRSelhMo6Ou308UcJSEACEpCABCQgAQmcLwEjLM6XnOdJQAISkIAEJCABCSw6gQ6O0macrxPpCA7rL8ZujF0WK//OHc/nK2Js742NLHqnl/iGSYE0HdGCtFDUIsCB/1DsE7FbY7xZz1v2MHqpvRjVUJnpiU1Nvqgj1F9MwTQd8aJSjZgx++3FOhIt4kS74/uUp6f+xGxkRoSLyZGDs+IF0RWzdSlyT8SPRHK8GHExd/tafqKI9n+JUaOC/nMCtSrYUp+BZ22aAqojxHXZe1PBjbVRjhsC0HMx1hJraiJrzvoVp5uJ/iYBCUhAAhKQgAQkMK8EFCzmFacXk4AEJCABCUhAAhJYAgL4yyns/LIYRYIRJahlQMFpHNk/E/vnsW0RN8ZXY5QFTvuIFjimvxtL4evZIth/ESOV1p8U2w9me20xfrxZv6MonH3qkCJmzO49v7rVswJFY7Y4xmwkRaF+zIokZZRF203vyndECFJb/WaMouIbYqR6QjXhO4510hexpQj4+XXu1Kftqj1FdAUCBYxYG2WDJXVAdsdYS6wpGXbV6PswEpCABCQgAQlIYPkTULBY/mNkDyUgAQlIQAISkIAETk8AB/WRGMW3cbS+MkbKm9aGgx4H7Po4bI+txrfGi0gDHPqNiBc4q0kVdXfB6jPZIgQg9OCkhtdHCoDvynb7gkzCWeGjFCkqx3KP5IWqbI79TtEP3vJHkCAtEf0iMuBvYqT6opH6iagA7MVwD9ucBIpC26RQYy0wxq0NgY+1g6DFWmJNGV3hfJKABCQgAQlIQAISWFQCChaLitubSUACEpCABCQgAQksAAGc1LwdToHgtbEPd7gH+fpx1lPv4JRCGAvQp2V9yYgXOKKrhXCBo5/vRGAciOHM3hn7X8V+xAxEBFJvfV/x25ez3RqDK6mZ3lls2U+dDK5JSibSc9FwgJOCaLbAdtrHYwdjryvO4/6cwz4c5bzpz2fuyW+M6zMx+od4gUAxK07kWYpLKlaUIE6zhTFjiQjF2LU3hL4vxVhLrCkFoLOA6iESkIAEJCABCUhAAvNHQMFi/lh6JQlIQAISkIAEJCCBpSPAm/Y4skkbRK0GnO6t7bp8oW4Djm6OQbxY9Q3hIqJFyQEmiBY4qol0QDTAgc2b+JtiRFnsK35DPNgRo5YEzu2rCq4IC3fGiN54Icb/GzjJYU69DCI42H9PcR+2pO3aH6N2AlEW1NvASod5KWawPSFU5LPt3AkwDjAkbRpror2xdjiGtbTqCtSfO07PkIAEJCABCUhAAhKYbwIKFvNN1OtJQAISkIAEJCABCSwFAZzZRE7wRjhFpW9v6wTFuK+P7Ynx5r6tINASocAe+JUplvhOwW5EDBzcsHux1vaLkRJwRNQgCuLZGMIGzm5EDsajjITgWAwRidoJ7EeM4NhvFceXDvLy+icEpbb+OW4XRoBxoE4Ja4E10d5YO8wB1pLpoC6MtWdLQAISkIAEJCABCZwHAQWL84DmKRKQgAQkIAEJSEACy44ATlZSEFGTAUd4u2BBh38ohkOW321nSaAQDDo5r6mDUTYEBkSIU1pLBAe/H4211ppg3EqRwvRDZzkmF3AYc590X6yFTu2PijXEWnI8LgC0p0pAAhKQgAQkIAEJnB8BBYvz4+ZZEpCABCQgAQlIQALLjwAO9EdipBMi9dDPxUhrU6YlIk0RDtuLUnx4TwpvmxZqEcawQ42Jdke4jvFFGIfM+dm5X6wB1gKtjKghKua3Y38ZI3KmVYxahN55CwlIQAISkIAEJCABCbxIoCx6Jw8JSEACEpCABCQgAQmsdAI4XxEhroxRWJiGI7Z8g59izhti1ExYFweufwuv9BG3/2dFoJjr64q5zxpgLdBYG6wRGmuGtcMaUkQ6K7IeJAEJSEACEpCABCQw3wT8J22+iXo9CUhAAhKQgAQkIIGlIoCTlaLBT8dI/fRU0ZGyeDBpon4qRh0FHLX+LbxUI+V9F5sAc505z9xnDZQp08q1wVphzbB2WEMKFos9Qt5PAhKQgAQkIAEJSGCWgP+kOREkIAEJSEACEpCABLqJAI7WF2KfiH2qcL6Wb5DznLfG3hgjNY5RFt008j5LRwIt0RXMeeY+a6BsrA0ECtYKa4a1o1jhXJKABCQgAQlIQAISWDICChZLht4bS0ACEpCABCQgAQksEIF6rjsSeyA20eEeFH6+KnZ5zL+HF2gQvOyyIcAcZ64z55n77Y01wlphzbB2bBKQgAQkIAEJSEACElgyAhbdXjL03lgCEpCABCQgAQlIYIEINHPd8Rh5+n8+9idt9/nhfCdP/2H25w10UuWceKs8xbgXqFteVgILTyDzufUmZf2WNdl5S4y5395YI9VizbB2bBKQgAQkIAEJSEACElgyAr5RtmTovbEEJCABCUhAAhKQwHwQ6CAwlMW38dw+GNvfdh9S4rw7tj22PlY6dWcPa3P4zkcXvYYEFoVAh7nL3GaOM9eZ863poOgTa4M1wlqx2PaijJI3kYAEJCABCUhAAhI4HQEFC+eHBCQgAQlIQAISkEA3EpjOQ5H+5o7YoeIBydVfNpy3Pxi7Msbb5zYJdCMB5jZznLnOnC9buRZYG6wR1gprxiYBCUhAAhKQgAQkIIElJWBKqCXF780lIAEJSEACEpCABBaIALn4n4ptin0j9srYcNu9bsv3z8coNExKnBNpoco31U0PtUCj42XnlcAcUUFEV2yIXRNjrre2ci2wNr5XrJVT6lc4/+d1mLyYBCQgAQlIQAISkMBZEDDC4iwgeYgEJCABCUhAAhKQwIojgPjAW+QPx/4oVib2P9jyJDfn8xtil8SGYielhlpxT2yHJfASAeYyc5q5zRxnrpetXAOsCdYGa4S1ckKwE6QEJCABCUhAAhKQgASWioCCxVKR974SkIAEJCABCUhAAgtNgALCGLn5v1TcbEfLTQfy+V2xwRiVto0+XugR8fqLRYC5zJxmbjPHmetlK9cAa4K1Ua6Txeqb95GABCQgAQlIQAISkMCcBBQsnBwSkIAEJCABCUhAAiuewBypa3DEjsbI0393bKTDg742+/ibGAcvzt2TmgW4V/zUWPEPwBwsrOcc5iNzmTnN3GaOtzfWAmuCtcEaYa2c1EwHteKnjg8gAQlIQAISkIAEViQBBYsVOWx2WgISkIAEJCABCUjgLAnwBjk1Kr4Z+8M5zrkp+0mdszXGm+imhjpLuB62aASYk2czLzmGOcxcZk4ztzs11gJrgrXBGrFJQAISkIAEJCABCUhgWRBQsFgWw2AnJCABCUhAAhKQgAQWiAB5+SmovTf2QOzbHe7z1uzjLfSdMfL+2ySwHAnM1pgoIy7KDnaIumAOM5eZ08zt9sYaYC2wJk4qNr8cH9o+SUACEpCABCQgAQmsLgLm6V1d4+3TSkACEpCABCQgga4lMEcKm5k4dKfy0PtipMC5NsZb5605/V+d76+L/ZfYnthEzLfOu3amrKwHK+b12RbE5oW0dbFXxX4hhiDR2mr58tliLbAmpnL9s732ygJnbyUgAQlIQAISkIAEViQBIyxW5LDZaQlIQAISkIAEJCCBsyUQh2xZy+LJnPPJ2BNt596c7zfE3hC7PrY2djbpd862Cx4ngcUgwJxl7jKHmcvMaeZ2a2PuswZYC6PF2liMvnkPCUhAAhKQgAQkIAEJnBUBBYuzwuRBEpCABCQgAQlIQAIrnEA9/eft8mdivx+j2HB7e0V2DMeujhmJvMIHfBV2nznL3GUOM5fbG3Oeuc8aYC2wJmwSkIAEJCABCUhAAhJYVgQULJbVcNgZCUhAAhKQgAQkIIGFIFCkvSHNE47ap2Mfix2M3dVyvzfnMymjcPjyd/LZFjpeiC57TQmcLYFynjJnmbvMYeZy2ZjjzHXmPHOfNdAwFdTZ4vU4CUhAAhKQgAQkIIHFJOCbY4tJ23tJQAISkIAEJCABCSwlAXL1U59ivHDa/tdsqV/R2n4zXz6EQzdGnQtqYPAm+kl5/ueol7GUz+a9VwGBDgW2ESv4n44tc3ZHjDnc2iiu/dcxinEz91kD1q1YBfPFR5SABCQgAQlIQAIrkYARFitx1OyzBCQgAQlIQAISkMA5EyjeKKcIMSlx7o89Fdvc4UI/nH2IFdtiFDC2nsU50/aERSLA3GSOMleZs8zd9sYcZ64z55n7VaMrFml0vI0EJCABCUhAAhKQwDkTMMLinJF5ggQkIAEJSEACEpDACibAm+UHYqTFoUDxw7H3xoiiKP82viyf74j1xR6JjcUo3H2ilW+6G2mxgmfCCup6h8iKsve8gLYpdmOMCAvmbtnKOc0cfzRGZMXRmNEVK2js7aoEJCABCUhAAhJYbQQULFbbiPu8EpCABCQgAQlIQAKkxSmjJz6bzzfHKFJ8SYGGGgC/Ensw9j9iIzHOsUixc2c5EeB/OaIrdsb+QeymYl6XfaTINmIFc5zjiC5iHtskIAEJSEACEpCABCSwbAmYEmrZDo0dk4AEJCABCUhAAhKYbwItaaF259qkyeHt9OOxZ1vutSufb429v9j+QLaIGKTcOamd5s33+e6611ulBOaYY8xF5iQryF/2AAAZuUlEQVRzs3WuMnfLxpxmbjPHmevMedNBrdJ55GNLQAISkIAEJCCBlULACIuVMlL2UwISkIAEJCABCUhgXggUosVUHMG8gf71GJETb4jdHiNdzhOx62L3xiZjvJVO9AXO34Mx0knZJLBUBBArKK7NnGRuDhZzFYHt8RhCBrUt7ox9I3ZP7FDmvRFCSzVi3lcCEpCABCQgAQlI4KwJGGFx1qg8UAISkIAEJCABCUigmwgUDlwECOpUIFz8cYw30REraLfEfiy2NcZxOIj57N/Q3TQRVtazMPeYg8xF5iSfmaPMVRpzlznMXGZOM7cPKlasrEG2txKQgAQkIAEJSGA1EzDCYjWPvs8uAQlIQAISkIAEJDAVBM/F2FJk+4uxfx+7IkZtAOwdsT+LfT6Gg7iMvJjOZwsYO4cWgwARE0RSDMeoVXFl7N2xHy3mbdmHPfnwn2IU134ghqjB3LZJQAISkIAEJCABCUhgRRDw7bAVMUx2UgISkIAEJCABCUhgIQgU6aFIq7M3dmeMt9I/0XIvnL2kiCJl1AdjOIrLdDw4kHEk2ySwkARKsYKoCuYec5C5yJxkbrYKEsxd5jBzmTk9Xszxheyf15aABCQgAQlIQAISkMC8ETDCYt5QeiEJSEACEpCABCQggRVKgCgJbKjo/19ly9/JFDN+Y+z6Yv+ubI/EeOnn4dixGHUBGiv0ue32yiDAfCOy4rLYK2IIFT/U1nVEim/FmLs05jI1V4wAWhljbC8lIAEJSEACEpCABAoCChZOBQlIQAISkIAEJCCB1U4Apy7pnUifw2eKav957KLYbTGKHJftp/Lh78V+K8bf0g+meDfCRdM32Vf7NDr/588c6nQykRWIFZtipIH6vtjPx7a0Hcx8fbaYsy9kOxajoDxz2iYBCUhAAhKQgAQkIIEVRcCUUCtquOysBCQgAQlIQAISkMACEiC1zr7Y4cIBTOFi0uq0NxzG22Ok5nlz7PLYhjidfRloAQenWy89h1jBXNpQzC3mGHONOdcuVoCFOcpcRbRg7jKHrVvRrRPG55KABCQgAQlIQAJdTsB/qrp8gH08CUhAAhKQgAQkIIFzIkB6p4nYxTHqBTwT21VcASfwmhgO4vWxfxijADeFuJ/m2DifcRZPG21xTsw9+CUCrfUqECmuit0YI9KHucXcuzRWzkXOZI4yV0kDRYSFKcqcURKQgAQkIAEJSEACK5aAgsWKHTo7LgEJSEACEpCABCSwQAQQLChmTKonHMS8uf7RGGIFjTfff6L4fF22d8W+GMNR3Bd7LmY6ngUanC6/LOnHECR2xphb74i9JXZF8dxl7qhyLv7v7Ce64jsxUpoZWdHlE8THk4AEJCABCUhAAt1OQMGi20fY55OABCQgAQlIQAISOB8COH4PxL4RQ7zYH/uFGG/Al8W5uS6OZMQLjudt+O/FPp1Ii6NGWZwP9lV9DnOLyB1SQFHoHdGiFMZKMOXco9bKr8Z+J0a9CupWKJKt6unjw0tAAhKQgAQkIIHuIGANi+4YR59CAhKQgAQkIAEJSOA8CURYqGAdGsWMibLAIfz7sf8eG43tbjuWt9tJyTMYWxsra1r0RrjACW2TwOkIlMW1y5oVzCHmEnOKudXamHvMQeYic5K5yRxlrtokIAEJSEACEpCABCSw4gn4D9SKH0IfQAISkIAEJCABCUhgIQlEdMCRvCvGm++XxHj7/SMd7kn9AJzH/yr2fIyaA6SXmozxRnzHNodYspCP5LWXiECHAtv8PzYcQ6Rgbr0s9uuxTTEiLNrbx7ODKB7m1ldjuzN/EDBsEpCABCQgAQlIQAIS6AoCpoTqimH0ISQgAQlIQAISkIAEFpAA6XYeLZzE12b7ZOwHYziaWxsOZux9sfEYQsU9sbtj1B5oLmAfvfQyJdBBpCh7SrQ7oT2vi91ezKd12d4wx6Mwnz4TI0UZNhKrL9PHtlsSkIAEJCABCUhAAhI4LwIKFueFzZMkIAEJSEACEpCABFYRAaIjSLmDCEFdi4ti1LOgIPIHY7wdXzbEjctifz/2YPF5c7YU5Sb6Aic1xbmbeTOera3LCZQRNBEuKMjO+LNFvCKKgjmEEb1zU+z/xphD1LIoG1E6f1XMIYQv5iBz0TRQXT53fDwJSEACEpCABCSwGgkoWKzGUfeZJSABCUhAAhKQgATOh0A1Jz0XY7stdjSG0/k9xT4KIlN8e1dxcRzQl8YeiOGQfipG+h6czgMU5s4W0QIzZdT5jMgyP6eoYYJAgW2JITIQVUGasatjW2MfLrY8DXOHOYRgwTxjTt0V+0TskdjhGHUrFCuW+djbPQlIQAISkIAEJCCB8yOgYHF+3DxLAhKQgAQkIAEJSGD1EeCteJzJ1KpAbOBv6S/HHo+9OvbW2HTs2dhtBR4c0r8Y+/MYb8rjaCbtD6LF9hiObK5Fuh+uj3Axp3ix+pCvvCcuRIqykDZpwxAqEKUYa8acz9SreGfsR2LMkbIxdxC5aKQSo+g28405RhooRAxTi628aWGPJSABCUhAAhKQgATOkoCCxVmC8jAJSEACEpCABCQgAQkUBHAYIz5Q/Bgn9I2xr8Wejl0ea68rQCHl98YokkzdgVtjOKARLXiDHqc2jmiECtJGkRKoFC+EvkIIFEIFKZ+IjiDyBtGC8b24GF8iK66LfSuGiMGcYG60NuYOkRSfjf1tbKD4zlxjztkkIAEJSEACEpCABCTQ1QQULLp6eH04CUhAAhKQgAQkIIEFJIAD+bsxhIebYwgOD8VwWrc3nNYfiCFYUH8AQYItb9tT44Jr4ejmd4QPUkeNpv6BqX8WcADn69IRKxAWSPOEXVWMKcIT9U2IqEHYYntFDIGLMWdOtLf92UFEBeIGc+SbMaIuiMCxSUACEpCABCQgAQlIoOsJ8NaPTQISkIAEJCABCUhAAhI4A4E4pTsdgTjBW/S8OU8aKJzQ1Ln4pdg1xQl8J+0Pf3sTTUH73RhRFoMxhAtqE+D0vidWCh44vHFeI2ZY42KJZugc4172hjFFlNgZKwtlIzTcHkNsotYJQgWpwpgj/6Q4EQGCMT0So0g77cnYfyi+I1zcG2OOnDYNVFnUe4nweFsJSEACEpCABCQgAQnMKwEjLOYVpxeTgAQkIAEJSEACEuhWAnM4hptxaON8fix2IFY6qD+ezx+N8dsNHZhQaPlTMRzWz8RwcqOI4AAnnRDXIvoCZzaCxsEY6YJMFbX0E6ysT8H/UjtipSBBfZOLYkTJIECxnwLZu2IIVh9q6XopXCF2PBrjO3OG1E/fLs7nOtXMO2uaLP2Y2wMJSEACEpCABCQggUUioGCxSKC9jQQkIAEJSEACEpBAdxLAoRzRgrfgeSseYYGIC4zUTggMPxNDhMDKgsrUMeAtfKInSP9DKqFPxm6K8aY+tTBwjD8YuzaGWMG1SQ9EkW7EDB3ZizulGA9SO1F/gvFBrOD/qb2x1xXjwdgRGcOxPxgjtddrYggTjPk7ii5zDvVKsI/FiKqhqDYpxsqICguwL+74ejcJSEACEpCABCQggWVAQMFiGQyCXZCABCQgAQlIQAISWNkEirfgcTATcUFExP0x6lnsiuGoJi0UkRb/KEaap32x18dIA0QkBn+Xsw9HN2mAeCP/yhjXWhPDOU6x7udjd8V4g7+sgYEoYls4AogJZQ0KImjeEqNYNsIEIhLjc0eMSBkEKEQn5sKPxMoi2ggcRE4w9qSP+lyMyAoiaL4T210cy5gqRC3cWHplCUhAAhKQgAQkIIFlTkDBYpkPkN2TgAQkIAEJSEACElhZBIqICxzPRFngwMYhjRP6gRjREYgSOL15656oi/JvciIxePOefbyZTzQGdTFID8X1KOaMOEH6IIo3z4oWRXQHjvGOURfWODj9/JmjRkUZTcHYMI6kd0KsgP8lMQQkxApqlpAGirHiNyJl3lR858acz3gy1ow512UOMBcQPEgJxhwhnRSRFYoVpx8uf5WABCQgAQlIQAIS6HICChZdPsA+ngQkIAEJSEACEpDAkhBAPMARTZofUkURMYH9cgzH9fcXvUJ4KBsFuBEl2IdwUdZC4A1/nNkU5SZKg++lg/tr+YyAwe/ciy3FnnV8n9+wIyjAGZGCVFxsqUOCCMFnoileHkNsQKRgHxETRFAQWcE+ojFaWznG27PzszEiZBg3xAoMccoUX+c3Xp4lAQlIQAISkIAEJNBlBPiD3CYBCUhAAhKQgAQkIAEJLACBvL3fWqCZt+ypf8Db+a+OkfLpbTHSCdEo0IzggFOc1EE4wcs6GIgXXyzOozg3TvTp2O4YqaQQMEg5xNv81LlALJmxYPPZDWoxTowVYwR3aku8thgLIip2xRCUEIeoOULUDPUoNscQkBCa4I54wVggZCBQ0L4S+1KMlFGcR2QGURaM0WkLqRsdUxB0IwEJSEACEpCABCSwaggoWKyaofZBJSABCUhAAhKQgASWgkCRcoi/u3Fi4+xGVCDagi2O6/8Ye3fhvC4joO/Ndz6Tiui6ot9/mi3Oc4QKnOJEUuAEJzUUxZqpm4EAsieGYxyRA4d4ReGi88gXQgU/whrxASGJiAgEhptjr4yRCgpxicgLxCSEC0SiDxdXpeYIKbtgTQovGp+55udj/y6GUIUIQkQFW0Sn2RRQihIFMTcSkIAEJCABCUhAAhIIAQULp4EEJCABCUhAAhKQgAQWkEBLjQT+9i6FC5zepA+i5gEphnCU3x5762m6Qson0hThDN8dowA3QgU1FKifcF8MZ/hTMRzipJXCsc5vGM5xC3QD6tnjREWU0S98RghiPBCUro4hJt0S4zdqiCBcUGh7VwwhohyLfOzYvpy998QQjh6LkfaJ8UBsKmtVzKbtUrCYC6H7JSABCUhAAhKQgARWIwFrWKzGUfeZJSABCUhAAhKQgASWggAOaox0Tjit2fLmPfULvhd7NEbkBCmEiKz4qVhZlJn0Ql+IIVjwNzyObyIvcLBznV0xogBwjD8XI6UUb/7jOCeyA6Fibxz1HFvWSygd5l1d76IliqIUjKgxQWonBIqyPghCETxJ6XRZDCGJ1FC7Y9fEKK5NNEz5/xNjAVfSeJFGioiZ34sRaUGKL6JhHiy4kyqKc8vaIl3NO89pk4AEJCABCUhAAhKQwHkTULA4b3SeKAEJSEACEpCABCQggfMiUAoXiA5lPQNSDeFQ5zcEB4QJxAec3Q/EqJGAM7xsvO1PCiOiKx6J4WAnlRHCBIW5ib64Mcbf+2U0B8WeETKI0EAYoXD0gTj0y/6U25MearlHALREsLT2uxQnyi2c1sfgDBOECYqfl1EP789nmGJl5AXHwxWOpchR3oOxIIKCGiOviZEuilRcRF5wTSJfGBc4n7ZOxUmw/SIBCUhAAhKQgAQkIIFVTsCUUKt8Avj4EpCABCQgAQlIQAJLS6ClMDdv7GO82f+q2K4YkRcICT8TI03R64vePpktznVSPyFIEKlBwzlOTQve5sdZjtjB2/9EXyCOfDNG6igc8aSPQsSgcSw1L9g2V2rqqCLVE1ETCBMIOmxpiBPwQwQi1RMcKX5ODRCiWBAdOBbhgZoV5YtdREYgLBHJgghEtAUNjvD7WIz/qa6P7Y49FENkIoIGg6URFQU0NxKQgAQkIAEJSEACEjgTAQWLMxHydwlIQAISkIAEJCABCSwggbYIAf4+521+0gyRhghHOW/z4/R+XQzhgugAai6Q1og0UggRRAFwPG0ihvMdRzzGNUkFhXCB053i3IgdiBlfLfaXEQNlbQciMbjnbO2L4hrF5WfTKJW/lceX0RlllMhsoW/EmDM57AvBpvUe5TXK6Ij2e7XW4SjPK/sBm/J4aoKQWgsGb44hSvD8FNPm+dkPQ46HDYZgA3va/hhREggbRK3AkJogsEGouLvgwj0Qjjge9o0zPXNxfTcSkIAEJCABCUhAAhKQQBsBBQunhAQkIAEJSEACEpCABJaQwBwpjegRwgXO8LIGBW/+U8uCGguviJHmiFRROMuJCPiBGBEENCIucKDz9z4OeFIXEWGAuIGwQbojaixgRGgQLYADHiGEiIJPx6h1gZBB1AbHYOyjX2WjT/QRRz+OfBz2nI+AQJ8QBNhHxAet/P+jjDogooH+IQaUqZO4D/sQHxBe6ANRI2Ur+8B9MO5DH+jXB2Kcj7CAwMMzc8xNhZEGCy6IEDwz/Ogf/SnrVHAfIlD+sugTohH8KL79cIyUXdSuoE9lDYzxiBT0yyYBCUhAAhKQgAQkIAEJXAABa1hcADxPlYAEJCABCUhAAhKQwAISwAGOAIGTHWc8jnuc7U/FSEmEs51IAY4hVRFOdsQNHPakgMKxjsP/6hjiBmIF10Q0IEqBNEY46fmfAOf922OIHwgPOORx4pMSiagEBAciEEizxHeuwz247q7YYzH6RyFrzqW/r4zRJ45FQGh36HMMAglbnoG6DxyDKMN3okZeHtsdQywgfRPH8sykryJCAsGD7wg0PBepnxA6EBkQExAsEELoN8/MMdyD56TvHMO1EVxo3AOBg3ROpMsi9RbPwDMjWnAc4kpZm2K2gLkRFQU9NxKQgAQkIAEJSEACErhAAgoWFwjQ0yUgAQlIQAISkIAEJHAhBM5Q1Jq0SmWKo7IuBQ5zIhco8oyDHec+VtagwAn/Q7HSOU/0Ac56BAcc+wgDiA04+hE0cN4TccFxOPpxxhPFQS0NxINPFc+H8IEjHwGF8xBJEEcQPXDovzOGwICQgHByW4x+cQznsf1KcS2EBe7DcQgEiAL3FsfRTwQQ+sy1uQa/czxGeibOQ7ihfSiGSELtCM6l7zwLAkpZkwIm9BFeCCmw4TmIriDtE0LI7thfFPfl+fhOTQruzfHwhT3jcCIt1XIvSv4iIpsEJCABCUhAAhKQgARWBgEFi5UxTvZSAhKQgAQkIAEJSEACEMBRjtMeJz9CAw1n+j0xHP58xplPlASCAlEKpD8iyoBoA87Hic9xu2OIFggipHbiPFIxPREjSuG9xTkIBogQr40hDODwR9hAzECI4HcECESPXTGc/4gBFLbmXq2tLA6OuNHaEAG4JtcgaoHoEa7B+RxL3+6I8cx85t4ICQgU74oRIfJXMZ6F50Uc4TiuwbMjVpRFtYk8QcDgHP4f2htDtCCaghRZPFNZkwOBokxHVe7LLpsEJCABCUhAAhKQgAQksBAErGGxEFS9pgQkIAEJSEACEpCABJaAQKIxcMTTyjoQpGgi0oGoBMQInO7swxFPuidECVIi4fhnH5ENRB1cGyNaguO/HaMeBM79x2MIEkRoICYQdYAQgi1EQ1TASOmEqEGEBILGdTGECOpuIKTwfw19R2zhOek7USgILaR++psYYgn7ECg4nuekaDlCD/vK+hsUDG8t7L0Qz+U1JSABCUhAAhKQgAQkIIEOBBQsnBYSkIAEJCABCUhAAhLoUgKFgIGwgMMfUYGoBJz9RGnglP/RGKmfSKGEgIFogRhBdAYRCdTMYD+RGmXkBMcQxYCYgaOfFEw0HP6IBfPRWq9FRAQiC/+7UIcD0aGMxCAyAiGC1FE8E1ESiBocw37SQpEq6s9iiDk8E6ILUSEIIQguNQWK+RgyryEBCUhAAhKQgAQkIIELJ6BgceEMvYIEJCABCUhAAhKQgASWNYEIF/zdj+Gwp9A1Dv1dsVfFEAeIoLg5Rvoj0i0RcVHWfeDZEDz4jjDAuTSEC5z+XI+GuMHv89Far0XBbsSW1vvyO4ILggON1FZ8J6KCtFWkuLo/RgQGIgq1KHYXfeZ6iBsWy56PkfIaEpCABCQgAQlIQAISmEcCChbzCNNLSUACEpCABCQgAQlIYLkTKKIuSO+ECECtCkQKHPzUiuDz22O3xhAuqBmBEblQFvdG5KA+xZ0xIh8QOziP/y3K1FJfzuf3FCxI3TRX7bzW3/42x701VqZyKmtrIDoQyUG/vhkrC2ETLUIkCLUvMISKbxX94nn+rugXn6npgbhSN5qiGBU3EpCABCQgAQlIQAISWIYEFCyW4aDYJQlIQAISkIAEJCABCSw0gSLqgloXpHoiJRTREUQosCUFFIWvSQeFo586GERZUCMC8YAC2J+OIV4gbhDNwDHUk/h47Lux98eIgOD8XTEiGzifRo0MIjN2xxBOuPZnYhT0/kiMuhnUliDqAxECkeIDsa/EEEk4n2tzDOeT/unpGCmiiL5AOGFLSihqXkxHqEAAsUlAAhKQgAQkIAEJSEACy5iAgsUyHhy7JgEJSEACEpCABCQggYUmEOGCW/B/AVEQGDUvSB3FPgpdT8cQCK6OkRZqLIZI8HCMqAaEDQQPRAcEEEQDhA6iHvhO9AXX5TM1KGhEb3BtIiyIgOAedAThAbGE7wgSCA4IERz/ihjiB/UrSP/0VAwBhOvSZwQJUj2V1+XapH0qbulGAhKQgAQkIAEJSEACEljuBBQslvsI2T8JSEACEpCABCQgAQksIIFCsJjrDggUtFLEQAzgM+mYEBOof1HWxkDkQDQgooHfEBU4n+/s5zP7aOVnziXCozwW4YPv7Ed8mK01EaMOBb+RlqrsQylOcL3yusXlX9ooWJyCxB0SkIAEJCABCUhAAhJYtgQULJbt0NgxCUhAAhKQgAQkIAEJLD2BlgiMMqVSWcB79juplkgvVaZcav18Nr1vE0y4dut9+Fz+z1L+dtLvChJnQ9ljJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIIGVQeD/A3Xdt+WbMXRnAAAAAElFTkSuQmCC" }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO29d3wc5bX//57Z2d6LpJW06r1YknvDxpgWaoAQAiEQkhCSACGFQBokN8lND/leCAk3JDf93pRfCKElhGIcmsEYV7lJlqxi9bKr7X1+f6y8tnGTDUa2NO/Xa162ZueZObO789nnOec85xEkSXpEEITzUVBQUDgKsiw/J6jV6olEImGZbmMUFBROX9RqdUAEhOk2REFB4fRHnG4DFBQUzgwUsVBQUJgSilgoKChMCUUsFBQUpoQiFgoKClNCEQsFBYUpoYiFgoLClFDEQkFBYUooYqGgoDAlFLFQUFCYEopYKCgoTAlFLBQUFKaEIhYKCgpTQhELBQWFKaGIhYKCwpRQxEJBQWFKKGKhoKAwJRSxUFBQmBKKWCgoKEwJRSwUFBSmhDTdBpzOiCoJt6cEu91GIhphsL+XYCBIWpan2zQFhXcdRSyOgNZk54Zb72TliuUM9nQwOjqOzmimsKgEs9nIyEAvbTu2sXPbZnZv38rAwBDpdHq6zT7tMNgL+MZ9P2G0/TV++N0forxDZzaCWq32JxIJ83Qbcrqgt7n5r1/9L8//8UEe/dtjJFJv+YoLInmFJdQ0NFE3p5mahibc7jyCE2P093Qz0LcPr9dLNBLguccfIRxLTs+NnAZc+5lvE9vzPLUX3sJzD3+ZN1r3TrdJCieJWq0OoFar/YCsbJntE//xkHz15eedcDurM1eua5ovn3vZNfIfX9gi/+yXD8smnXra72c6t+//7h9ynkUjv+emL8gffN8l026Psp38plar/YqD8y0snFvNU/9cc8LtJsaGGRge49Jrb+KVv/6MOz7xCYLRxCmw8AxBVJNrhlF/nFgigU6jnW6LFN4mis/iLQjIpNPyCberW7iaL3/tXn5731d5fu2rp8CyMwtR0pNOxEgBVqMJ/1Bwuk1SeJsoPYu30Lq7j9VnLz5sf3l13ZHXeRRELrnhM9z1hdv4+q0fVIRiEpXGRDo5AUBBUSmDvd3TbJHC20XpWbyFX/3o6/zgoV9SNfdpNm3eisHiYsUFl2JIjfLFT99B4qBOh1pv5vav3YdLGOXTN11HKBKfPsNPM1QaE3I0CIhUVRbz1z1d022SwttEEYu3MDHcxe3Xv5dlq99DdUML0aCP/3vgG+zYufuQ45yFFXz9Rw/y5j9+w/1/+DMnMXKZ0ai0WuREEoOrBFNyiGF/bLpNUni7KNGQE99qF66Wf/PYs/LSRS1vz8OsM8l2m2Xa7+dUbJbiefJPH7xPXv2B2+Wbb7pmSm2MVqds1GsP25+XXzDt9zPbNyUacsIIXPShT3PXnbdy7yc/yLr1m9/W2c69+hPceddn3yHb3l1ElYRKPPrXR1SrSCXgkksv4KnHn5rSOW/83He47torD9kn6N38+bkXMKpO1EIBtVp9oo0UjoEiFlNEpdZz+zd/ysqmQu74yAfpHRg5fiNBxfs/8km0koBKa2L+gvmHvBxPxDAaDIc1MzsL+NSXvs2Pfv5b3nv5xYe8llfexG+eeokLz1kCgM5kY+nZq9FppMm/7Sw753zMRv0h7Srnns2fnn2V+XMqJ6/hZumKlUhixm1rdrhZturAefYz9+xL+f5Dv+XcVcuz+ySdhR/+9km+9e2vTf5t4uqP3MaCeXOyx4gqFWVzVzPR9jID46HsfnteCbff831++NCvueg95x5yrdiR3o9klIQsYjAcGnotaVjMiuULAaiduwSzQXPQqwIf/dKP+N9H/45RqwIEzrro/Vz+3ssOc1KX1LRw021f4Kpr3n/YvSsciiIWU8DkyOd7v/wLyb43+OoXvzRlR2ZZyyrOXtxIPCmTW9rI9Tdee8jry1atprRpBZUeV3afzpLHD3/+a/ZseI4ffvPraGy5Bz4kQcUd93yLl599ioaWeagNdn74P3/isutu5vprr0RnyeX+3z/CORddyRfu+tyBC4la7vra11n73PPUNjRichVz///8gfd97PNcdO5yHJ5qHvztH7ngqhv52EevzzYzOIr43Odu5ec//iE3ff4rSJNP2iU33kHb2kcoqG9BQODO7/2cHIOKO77yzQOXVInYnUZ++4tfZPcZHYV8/6cP0/rSE/z4u/+J0Zl/4OEVNSyYP4clF1+L9aAHv3HFuYS9QT744QN2gcAtd32d4PgwANfc8gUKcqzZV0uaz2Z+uYH24ShOq4nV13yKK96znAtv/CxFTtOB9//SG7j361+lr3Mn+pxK5s+tP/6HOotRxOI45JbUcf+v/49///H/8d8///UJOTIXr1zN80/8FRmwuPIIjY9mX7MUNNCQk+Zb3/0JN37849n9H7vr22x86lc8+9wLaKxugoN7s3MqPPXLKZRG2bqzh2QyzjWf+hKbnvwl//vnR3A6crnxc//BK395gJ///JeY7c7sOc++6iP0b3qG/tEQyVSCj9/9Lf76k3t56pnncbryuP2e7/Kn//cV/vTnR7DZDwjXxdd9nI431hJIqon5x0jJoNJZed9VF/HXv/8LOexn/gXXYYvu4b8f+gVp6cCvf2V5FVvXPk73oDe770OfuYdX//Yz1v77Zcw5JYzva2P/21k9/zzkvo385fGXeN/7LpvcK3LDTR/jKzd/gJYLP4TNkPnlL56zkobcFJt3ZsKxVquNYMCfvc77rr+ZJ/7vN6hFCZ2zmA9dcyHf+NLdjPiC2aGTKbecL959K3d/4gae/edTBEZ7efX1rQBc8uE7WbWsZeof9CxBEYtjUNq4hPt++lMevOeTPPn0iWd1Oh1uhgd7AahrbEKj2z80ELj5c3fz+4fuY+MLT1I5fxUAZS1nc801l9G6aRMA51z6fpaddVamhajmE5/7HA/ffx9avQWjw8M580v43z/+DaNeh6moluUNLv74l8cwmeyEg+MA6G353HTj1fzsgQfQ6czkV7RQYQnwz+fXYdTr8LSsJFfu4+k167CYbQQCYwC4ihu45porKW1cyH/+4Ds89INvIwOXffgO1v/9YaIaE7FQmk/ddjP3/+AHCBorqnQAAI3Rzic+81kCgXD2vahoWcV117yXzW+8CcD5V36QxUuWAiBKOm654zZ++dBPefHZJ5m/bDUAy9/7Ubzbn2H77jbWb9lDc0MNolrPZ77yNUYHe5AByeCgsrIYtSbTGymsXUR9ATz/0gYMBj3XfvJu/vzgdwhE4liNWkKxBCDw8bv+g77W9YwHouhsRXz687cjAEZnMde9/yI2bmo94c97pqMM0o5CScMS/vN73+a/v3cvhtxy3n/TObhcOWi0b3GayTLxWJRQIMCEb5zxkSEG+vbRv6+bzs6drLzwKlK23Vx67mIMZhMLFsxnzuprKLGrcL/3enLmjNGzfT1Nyy/ktts+wf/++jecdf7FiPktrFpYjVpvYO68p1lx1c34Wp/h1Td3cF7de7jgiuv5xq1XE0um0evMrL7kSr5xyxUkUjIT3hEKyhuoa17EJ+7+Gr//4ZcZ8YXRmgxcdvUV3PGBC5ABg87MBZdcyu1XrUIGxseGKb/sYuYs6uS2L3yJ73/2Q9z6nV/y1AN3s3nHXlZd8REuXl7NZ27+Dq7q5dQsWc1jP/8mg+MhEJPI+kKa5y3k2tu/wuaX/km+LtNvKGtcyte/eS/PPf0MKy68GHtDlJaqHHT6i2lqeYmLbrgDKeblkg/cRFiTy/Ytr7Pqig/zvkuW0j8e5wM3fJRFc8p54fcJ7vnxL3n9kZ9x8UduZ978hZx33a0M7m3nuptu4ekXN3Pr5+/mvi/eTAIteZ5i9JE+vv3v1wEYGPKydMUK7PWrcWtD2IpqaWyay9Wf+jKaVAoZgdvu/R5/e+jb+COzdwLg0VCpVKovp9NpJXH/Lay6/DoqSwpw5uWj1ajxjQ7TuXsH7bt2sLdtF53tu+lq301X5x4G+voIhUJodAbyi8pYuPwcCl0mHv/zH/A0LKGhuoj7v/Vl1r3RyqXvv5bhttf5r+9/F8yFnH/h+ZjsuZg1Se77xpdZ9+JaKuadTWWRgx//x5dYv3EHl19zHXvWP81vf/d/mTiWLBAY3M1jj/0TGTDacjGmhvn1bzKvRyeGiEoOzl29kr/+/Aese2MLAKJKQ8+2F3nhpczDY3eXEOjZyN+ffA4A72A3pvxaFi9o4tc//gatO3az7qUXueKmT3PDxz6OgSDfvffLBCNxkskkFoPEr3/2INFECuQUHV19XHbVlaz5y8O8vKWL5QsasZXN5eaPXse3Pn8z/3ziCeqXnIfHpee+r3+RLTu7ufzq97P5+Ud46MEHKaxbyJJF83AVlBLz9nDft79JW0cPF199PXaLiaq6eh7/zX/xzHMvsH1HB5e//1q2v/QYD9x3H2UtK2hqqOThH9xL+959QBqjxc4jv/oJQ6M+AHZv38Z5772Wie7NPPCj79Oxz8tlV13FK0/8nrLmsxgKSSwp1/FfDzz87n/hTnNUKlVcybNQtlOyeZrPll/bMyR/4QufkfXa0332rUr+00s75f976jnZZTWcBvacfptarfYrwxCFU4IgCPTuaae6sZlk4vSefas1u7CYtdzzyU8yOhE+foNZiuLgVDglCMDuN55hY3eM91563nSbcwwE7vzeT9F5e9i4fc90G3Nao4iFwilBBmRZ5k8P38+l1330yDN2TwOaV1+NM9ZJf0ieblNOexSxUDglyLKMKAj4+nYzkrLjcZmO3+hdR+Sjn/okP/3RD1Gk4vgoYqFwSkil0wiCAMjs2tVBZVXpdJt0GMXNZ8PAJjr7vQhKOeHjooiFwikhFouj1+oACPjGMdns02zR4ax+z+U89+SjIOpBjky3Oac9ilgonBJCw0NY8vMAsDlzCHq9x2nx7tMyv5kNr29AY3eT8A5NtzmnPYpYKJwSYhP7SOhLqKysZvHcKrZub59uk96CCrtBYCQQo7y2lu6Otuk26LRHEQuFU4Oc5Gf/7z5u/+o3+eMDX2cscLpVykoTT4kYdFouveoDvPz8M9Nt0GmPssiQwqzlgutu56YbrmH7un/y3f/8rlIa8Rio1eqAIhYKCgrHRa1WB5RhiIKCwpRQxEJBQWFKKGKhoKAwJRSxUFBQmBKKWCgoKEwJRSwUFBSmhCIWCgoKU0KUZVkRjBlKZtbnASRJOmzfu4Eoimg0muMfqHDaIsuyKIiiGEmn07rpNkbh1KBSqUilUtm/BUFAlo+cqigKUFEAK5slaspzUckT+CZCbO6Al7aBL/huWa1wuiGKYlQRCwVMerhwASxrgNqaKornfxqHZzmCINKzZx1qIURw8HWe+deTPP1alM0dkFLKP8wqFLFQYGEN3HGNg6qG5ahzVuMsew+IegRBICcnh0QiQTKZIBELQ2Qve166h2eef4mfPQ6jE9NtvcK7hSiKUZUgCPfIsqxU+Z6FXLgA7viAk+pz7sNQcj2eyrOw2lz4/X5isRgmkwm/34/JZCYtCwx5U+RVX4nLGKTeuZWtnTJ+pRj2rEAQhKQiFrOUSxbD52+swN74ZexFq4jHEzidTkRRRJZlQqEQQ0NDbNiwgaKiIkwmE0ajkWQKNM5F6FRh5uZt5o3dEJgsMjUdzlOFdwdFLGYpdcXwnbtWoS77AjmlZ1FQUIBWq0Wr1dLe3k48HqesrAxRFLHZbESjUWw2G2q1Gq1Wi0arJad0FalIH2XmVl7YfMCHoQjGzEQQhKQSNp1lSCr4zDU27LWfYmhCQ05ODhqNBrvdng1xOp1OVCoVkiTh8Xhwu92Zat2iSDwep729HY1WT8P5P6ZpTh3vXX7g/EeLtCic+ShiMctY3QJLV1yEwTmHSy65hEgkkn3A/X4/BQUFpFIpurq6GB0dJZ1Oo1Kp2Lt3L9FoFJ1OR319PZIkodYakQqv54OrwWqc5htTOOUoYjGLEAW4/CwtYs7FFHpKGRkZYc2aNciyjCzLWK1WZFlGpVJhMBhQq9WIoogkSbhcLmRZJp1OE41GCQQCqNVqCuuuIq0pYHXLdN+dwqlm1oqFMyeXRcvPpmXhUlTSsV02ue58APLyC6d0brPFikZz+ML0U23/VtyFRSfV7q2sngtnLarF7F5AOp0mmUyyYsUKkslktgcxMDCAwWDAaDRit9sZGRnB5/Nht9vRarWk02mGh4dRqVQkk0ms9hwcNR/nwxcqvYuZzqwVi1QqRU9XJ7u2baaypv6Yx+a6CwBwuHKmdO6CohISifhh+505eSduKJCb5z7hNqIoolKpDnE4NpZBTmE9ksZELBbD5/ORSqUQRRFBEEin05SXl2fFwGw24/F4cDgcQMZ5qdFoKC8vx2g0olar8Xq9hMQqFjflYtIfaoNarcZqtVJQUEBBQUHWF6JwZjJroyBOVw7deztIJhLZL7CoUiFM/puIZx72opIyhgb7kSR19sHLpFCnYXLRO0lSk0ols2N/Sa1GlmUktRqr1U7AP0E8EQcBBFGkuLSc/t6erKDsP++ceQvpbNuFJEkEAn7kyV/7E3EaqtVqysvLqa6uxu12EwgEaG1tpa2tDaM2jqTPJZJMEQgEyM/Px2q1olKpCIVCxONxzGYzwWAQm82GVqtFEARSqRTpyRXGJiYmiEaj5ORkhNNsNpOSJbSWYgzaYQDy8/MpKyujtraWmpoaKioqsFqt9PX18Yc//IH169fj9/vf3geo8K4za8VCpzeQTCTQ6Q1EIxHmzF2Ap6SckaF+9vV0Mdi3D4B8TzGuPDdtO7bR2baLytp65sxdyOY31uHzjuPKzSMvv5Cujnb2de8FIJlIAFBYVEIoGKB5wWL6erspKa/EYDCi1xvwT/jwjo0C0DR/EbnuAna3bqW8upaevR1ceNlVtO1oxeZwnlA4UpIkSktLWbFiBbIsZ4cY4XAYQewknQgxMTGBIAhUV1eTTqfx+XwEg0Hy8vIIhUKEQiESiQSpVApJkrI9j3g8TiQSQRCE7N8Gg4Hc3DzkcBxRAI1Gw1lnncXy5cspLi6moKAAu91OXl4eZWVltLe3s3v3bkUszkBmrVhIkhqA2sYmhgcHsDmcJOIxujr2IB3kw4hGI/Tu7UCt1iCI4uRQQkaj1bFg6Qq69rQRjUTo7+0GQG8wEgmHsv+3O1xsXP8q9U1z2brhdRyuXAIHCQVkhEuS1DhcOYTDIfLcBax/5d+UVdYQ8E8wOjQ45fuKxWL09/ezYcMGCgoK8Pl89PT04PV6SSQh6u/CUeJgeHg422OJRqN4PB5kWWZ8fJza2lp0Oh2hUCjr7EylUsTjcWKxWHY4sXnzZlpaWjDodaTHB4knIZlMsmfPHmpra4nH43i9XiwWC4Ig0NXVxYsvvsjw8PDb/fgUpoFZKRYFnmLsThe1jc10tu0iJy+faCRMb/dect35jI0c+DLHolFEUSSVSlFSXkkyHqd105vo9Hq8Y6P4vONo9frsKtx5+YXYnS7UGi0qlYpYLEp5ZQ2BiQmGhwaQ1GryCjxIkkQymQQgHouyc9smEokEDqeLYCDA6PAQ7sIiqusa2b1965TvLZ1O09raSnt7e9YPkUgkSKfTjAcgOLoDKTCO3W7PDitee+01LrroIuLxOGq1mkgkgk6nw+/3o1KpMBqN9Pf343K5cLvd6HQ6ZFmmuLgYQRCIjm9hZGSYSDxz/S1bttDZ2Zm9x/1DmP1io+RinJnMyolk+7v1s+1LW+iCn38WhKrvsuyCT6LT6Uin0/T39yMIAkajEavVmn1/BgczPZr8/Hz27duH2+1GkqRD3rfx8XGe+58L6Onczjd/D4nUES+tcIYjimJ0VkZD9ucVzDb6RmHtFgjv/VU2VyKRyMwJGR0dxWQyZXsio6OjuFwucnNzASgsLGR0dJT29vasD8Pr9fLK2kdxiNv5+yuKUMx0ZqVYTIXyqtrjHrNg6YqTOndNQ9NJtXsn+PNa0MTbGe1+KSsWyWSSkpKSbJ5FKpXC5XIxPj6OLMtZZ6derycvL49kMklPTw/r1q0j2fs7dnTDxtNt3WOFd5xZKxZmixVBOPLtG81m0uljV3fJyXNjttoATih3QG8wkp6sXGUwmtDpDVNu+07QOwJPvAbJoaeIhINEo1EGBwcZHx9HFEWsViterzebfxGJRPD7/aRSKQwGAxaLhcHBQcLhMImxl9FG3+A3/4LZ10+bfczaWac2uwNRFHG4colGwllxMFmsLF25mu1bNlJSVomMjCvHTcB/aKWXsspqggE/giBS3zSXCZ8XV54bq82OWq1BUqtxOF0YTWZ0ej1mqxWnKxe7w0kiESccCmJ3OiksKiEcCuIu8JCIxyksKmXCO35K731XLzSXTNC88CLSKgt6vQFRFDGZTEiSlM3YNBgMWSes0WhEpVIRCAQIBoMM7n0Vofs7/OWFOC9sPqXmKpwGzOop6sVllbgLPeS68wmHgoRDmQKTjS0LUKs1aLVabE4nhUWljAwPEJzMC9Dq9CxefjbxWByHK4eAf4K+ni5qGpowW6zk5hcgiiKunDz0BiNWm52erg7Ov+QKAn4frrx8NNpMpKSgqJiyyhq0Oh2hYICS8gp0egOD/ftO6b0nkvDaVh/NpQEKPKXEUnqCwTCSJKHRaDAYDPh8PrRaLWNjY4TD4azj0+v10r75cYLb7+GpVwL8/tkDvQpBEBDFWdtZndHMWrEQBAG7w4WnpIy+ni6GBvpIpVLo9IbJ3AgnANs2bsBitbFn1/ZsW6vNgSAIdLTtxOF0gSwzNNhP84LFBAN+RoYGCAUDpFJJNDodQ/19WGx2YtEoiUQcSZIIBiZQqVRodTrisSixaJTd27dS09DEm6+9dNwh0Mnec05ODkajkWg0Sigq8/zLOym19VJR7CAWFwiEk2i1OrTazLyWQCCA1WrF6XQSCATo7dzKhifvJNb9Cx57KczvnoX0pFLk5OTQ1NRES0sLVVVVNDQ0UFZWhsFgyIZNDy4crHBmIQhCclaGTiVJIsedT3QyG3F8dATIPFAtC5YwNNCHIIqkUykikTC+8bHJdmryPUX0dnUCmbkiWq2OWDSKRqcjnUqSTCbxjY9R1zSX9p3bqaypIxwKUVBUzJYNr6PV6RCETDRhfxgyHo/hHRuloqaO8dGRQxK23gkEQcDtdlNeXk4oFGL37t1EIpnyVjoNXH2OhRveW4PFWYrWtRiDexU57kzxm1Qyid/bm3GI7v4x23Z084fn4M22Q/0UHo+H888/n+bmZurq6mhsbESlUqFSqRgfH+fxxx/n0Ucf5bXXXjslYqhwalEK9r5L1DQ00bZj27SEawVBwOVyUVZWRjqdJhAI0NnZSWIyJX0/ViPMKYPz58OiRjvOvDI0piJ0eis9+/p54unXeeb1AJ0DRw6RajQaqqurWblyJfX19dTW1lJfX09ubi6yLCMIAo899hi33XZbNn9D4cxBFMXorBp+nCokSY1KkohFI0d83e/zTj4wIrKcRlSpshGRqSCK4kn/GpeUlNDY2Iher2dkZIS2trbDhAJgIgQvt8Kbe7Q4/hHGot+IVr0RfxgGxyEcO/Z14vF4NnNUp9ORn59PRUUFy5Yto6mpCbfbTWtrK3q9/tgnUjhtUXoWbxOjyczyVefR1dGOqFKxq3XLUY+trmukbWcr1fWNtO1onfI1GucuoHXThhO2zWAwsGzZMsrKypBlmVdeeYVdu3YdfZEhUaSpqQm9Xs+mTZuIRqMnfM0jndNsNmO1WlGr1ezbt49Y7DjKo3DaMWszOI+FVnts3dTqDv1ljMWi7GnbSdvOVvSGo1d/sdodBIMBYNLZmOeecuTgRHohB+NyuZAkCZVKxbZt22hvbz/mUEilUpGXl5cdPhyMRqPBZrOdcM8gnU4zMTFBT08PHR0dilCcwczaYYjN4aTAU8xg/z7sDhdanY6xkWGaFyzh5TX/orKmnt7uTorLKunqaCMWjWB3umiat4h/PfE3mHzoct0F2VmhqWSS/MIiRJUqU3xGkuja04akVrNw6QoG+/swmS2UV9ViMJhIp2WsNhtWuxPf+CjhUAhXbh6CIDAyNIhGq81OxDoZfD4fbW1t7Ny5k5GRkWzOxNFQqVS43W40Gs1hQqbVaqmrq6O0tJTOzk62bNnyjvQ8FM4cZmXoFDJDAkmtpqSiisCED73RRO/eDhKJODl5bqLRKHmTFbK0Oh3NCxbTs7eD8bFRAhO+7Hn2h181Wi02h5Oyymq8Y6O0LFjC+pfXAlBZ20DAP8GOrZtIJZN4x8eQZZnc/ALUag1GsxlRJVFcWk4ymURGRpLUlFfVEvT7icfjJ5WoFY/HCQQC+Hy+I/op3ookSSxcuBBBEAgGg+zbdyDfI51Ok5eXx4IFC6ioqMBut9Pd3T2l8yqc+czapQD0BiPptIzJZCEUDNLb3UkiESffU0wkEkZvMNCxewcqtcSObZsyWZfxOLnufPw+74FfXUFAo9FiMluYM3chPV0djAwN4h0bZddB08rbdmzL9g5ceW6GBvpQSRI2uwOVpGKgr5eevXvQ6Q1otFrktMz42AgDfb2TodgDodT8wiIqaxuYt3g5K8+7iKq6BtRq9RHvc3/xm6lGYQRByM4TMRgOTUNPJpNs3LiRjRs34vF4+OAHP8jVV199SO2PZavOA6CkvGpK19tPeVUtpRVVaLQ6tDrdYe2rahuO2d5qs2Ox2g/bX3GccoknO0entKLqiAWJrHYHOZP1Wmcis65HARCNhHEXehjo6yUcDCBJasKhIIP9vdidOexq3Yosy3R37MFisdHb1UkoGCSVTmFzONEbDIwMDaI3GLI9ijdfexmAcDiIDHR3HDqzanigD4D+3h6SiQQ+7zj9vT2k06nMCmDBIK+sfRbIPORB/wR2u5Px0WFMZgsTPi8AA3292XOaLFZq6hu58rqb0Bn0dLbtZvOG1wj6T24R0v15EbFYjGQyediK66lUijVr1iBJErfccgt33nknHR0dvPLKK+TlF2aHOdJxCiAfjCAImYxWSSIei1JRU0dfTzdWuyPbm1JrNMc8R2FxKWYjIO8AABkfSURBVDu3ZXLOLVYb/sme3/7kMhA40uyVg0XWYrXjn/Aewb5MBOtgzBYbZos1e5395Obl07O3I3tfM21m86wchpRWVJNKJmnb2cro8BCJeBzf+BipZJJgwJ+tvxkOBQmHQwT8E8SiEeKxGP4JXzY1PJlI0N/bfciXxjs2SiIeOyxbMToZVt1fdzMY8BOLRYnHY9nrxaKZbM54LOMLGB8dIR6PEQwcuQRdPBZjYF8v27dsZOub69FoNJx78eXMaVlANBrJJptNFavVyvz580kmk3R2dh4yDNlPKpViZGSEG2+8EYfDkS2ek19YRNA/wYTPhzMnl1g0jEolodXrKPAUE/BPZB8eT0km58NTUpbdZ7XZkQGj0YTPO4bBYMQ2mUnrKS4llUySTCbI9xTjcOaQTCaIxzPOUlduPiNDA0iSGrPVhs2eybLNzS8kLaepqq1HbzBkk+tUkkRD8zxisRhqtRqjyYRao0GlUuHMySXgn6Cyth6DwUTLwsV0d+7J3n9pRRWu3Dyik0lt7kIPcjqNzeGksLiEUChAXn4BJRXVpzxt/91k1qZ7a7RatDrdMT9MnU5/XIfgO41KkhAnf5E0Wh2p1Ildf3xshG0b36CzfTfzlixn6dnnkkwkGBkamFL7/b+GyWSS1tZWAoHAEY+LxWJs27aNYDDIq6++Sk9PDw5XLr1dndQ1NhPwT+DMyaNp/iJcuXmMDA5kJ+LluguwOZzk5OXjys1FrzfS3bmHmoamyahPGklSk06lMVutRKNRGudmBMxdUIRao8FssdLb1ZEVGqcrh7GRYRyuXExmM1q9gVg0wpx5C0gkEkRCITrbd2Xtn7twKaKoon9fN2etvpDWzRux2u3MW3wWRrMZrU6PzeHIRLp27ciKeUV1Hel0GlEQUWs01M1poaNtJ/VNc0mnUuiNJpgs1LyrdQvyDMpUnbU+i+HB/my39WhU1NSd0DmdOXnUNja/HbMoLq1Ao9Wh0xvIfxtrhYSCAf7xtz/z+4cfJDe/gNu/+HUKi0qO2Uat0WCxO4nEU0yEoljsTiqq66id00J5VS3uAg9qdWY4IMsyGzdu5P7772f9+vUkk0lEUSQWjVJUWk4sGsFoMhOY8BGNRA4RZXehB5vDicFoZMfWTSQScRLxWKYXJGSCTFqdDmdOHl0d7ThcLv797D8RBBGL1cbOrZsJBvyIk2UB9keMIJN+b7ba6Opow+HK4eU1mWGdIIoIB0V3UqlM1Eqt0fDGqy+SX1jE6PAQ0UiY8dERRFHMTCbU6YhEDiwTrzMYKCgqpn9fD8GAn0DATzgcQiWp6enqpLyqlo62nZnFpdMzawgCs9RnMRXeGq505uQxNjKU/fvgMTVAgaeIbZs2kO8pRk6nT6oLajSbiYRDlJRXMjLUf/LGTyKn07zw9JO89uIa3n/DzfgnfDz5yB9JJhIIgoBWq6OorIJFy1Yyf8lZaAwGRJWEMycPo9kC6RQB3zjesTFAJhwKsmHdy2x49UV6uzsJhULZa40OZ96bnds24/f5CNonGAz4D4uW+H0+qusa2bDuJWwOJ/4JH1abHZBp39lKRXUd8ViMCe84lTX1WYexRqMlEg5htdsxGE3ZCuomswWLzU5VXSPxWBTf+BhVtQ0MDw4wPppZ/8Ris6PT6QhP2huPxenubCcWjTI6NEi+pxhRFFn/yr/RG4wUFBXjzMmlv7cbpyuHkcnQuG98DJ1OTzQSRhQF2ne2Zoaw3jHMFgvPPvkojS0L8Pt9mK3WU15q4N1m1mZwFpWWo9Pp0RkMBCYmyHHns23jG9TNaaG3q4O6OS307O3Irv+xv3Cvu8DD3j1tNLTM49/P/APIFOltmreQbZs24B0fxWZ3kOMuwDc+ll0ewJWbqV+ZSCTIyy8gFAzgzMljV+uWrA9k1QWX4B0bJZVK0rr5TSpr6kmn0/gnfEiSxMjQ4AkPTQ6moXkeqy+6nJfXPMOi5StZdNYqVCqJLdu28uqbG9nZP0LKmoPOnksy4M04OSN+5FQSKRmn3pPHsvnzaW5qJh6L8uLz/+Ll5//F3j1thzkBj4QgCDQvWEIsGjluz2660Gi01M1pIRQKHjLbeLYjimJ0VvosBEFg6dnn0tfbTU1DE2+88m9y8tzYHU52t26d/GXqx2S2UFZVQ/++HkxmC1W1DQQmfCQS8cxYdtJZqdXpGBrow5Wbj6e4lGDAT2VNPZvWr8tes6ikjPqmuSSSCZLxOFa7k1QqmRUTOOD4S6fSIGREyJmTSyqVoqF5Hm07tr3t+164dAW33PlV0BnZvGMX9/1/T/CSN02/qYBkaTPp0iZiJXNIuCtIFdaQKmkkmVtKorSJ/rSW17bvZO0/H8ff3838RUv4wIdvwZWXR2f7ruwSCEdDVKkoKa+kr2dvViCnG09xKQajKetE1ur0VNTUsXPrZpJJJYdkP7PYwanDbLEyPjrC2MgwyUQCT0kZkqQmEg5jtlrp39eDWq1Bo9USjYQz3WW7g3AogFqtIRaNZh+OXHcB4yMjFJeVY7U76OvpYmJ87ECURBCYt3gZYyPDGI1GRoeHiETCOHNy6evpytpVXlXL+OgIOr0BT3EpiUSCCe84npIyvGOj+P0T2UjJiSAIAqsuvJSvfOfHdHZ388Czr7HNGwFHPn3OKhJFDQj5FYi5xQgGK6SToNaBwYygNyE4PQgmG4K7FMFVRMySw57Wzax7+jE2v7qWqtp6PnLb5xkdHqRncvr+fnR6A3aXi3AwiCzL7Os+fYQCMtEdi9WeLUCUSMTp7mhXhOItzNp6FpBJ9w4GMrUlBTKJWqlUCpVKJB6PI6fTyDJYrFZCoRCynEZOy5mELAFAyD64Dc3z2L5lI3qDMRNNSMQzPYSD/B4Go4l0OkUiHkcQRVLJFCaz+ZByfVabnQmfF6vNnvHiR8KoJXVmOcR0ZrZqKHjkCMXREEWR62++jcvffz3f/9pdbGrvwHLJx6mub2RJuYe/b+ukXzBCInMvsncYOTCGYLBkTqAzIWi0oDch2N1kvJBp0rvXk971OumNz6KK+Fm4/Gzu/sYP+Mtvf8Gff/swAO4CD2aLlfZd2w/LORAEkdLKKva27z6h+3mnKK2ooqujnUXLz2b9K/9mzryFbNv4xpTa1jY2H3PC4ExkVk9R3x9zh0y6ztEeQu9Bx70Vnd5AOp3CaDIDHLMbfsiv6WQOxlvreu5PvNr/L0A8HsvmE5wogiBwxbU3svqiy7jrkzfQ1dGOxeHihuYSto4M8OvfPUvI50VOJpCjAUgksqIhqLWg1qDRaHGU1aI3GBnc9SoxRxHoTchBH+jNYLSSCnp57cU13PWJG/iP+36KwWhkZHiQN9e9TNvOI8+uNZnNyJOLD+kNxne8t2FzOA/5jN/K/gmB+6MqiVgMo8k8JTHWaLTHPWYmMmvF4p3AXeDBaDKxcf2r023KEVl53kWcf+mV3P3JG7Meff/4KA/c/UkwWCARg3g0M+yAySRHGUSRK1eqmFNtRNN8H3/6zf/Qvms70VgcrC4EkwNEETk8AaOZzFSL1YanpJS1//oH511yBQ/d9x369/Uc1bbc/EIklQqD0YRKkqiqa6R9UljUGg0FnmLCoRChYCCTgDU5W1Wt0ZBOp1GpJDRaLUaTiVAgkB3+QaZye667gGQyidOVw8C+Xpy5uXjHxohOhkJj0QiiSkWBpxgAQaXCaDKj0WpRqzUMD2aiUUazBZPJzNBAH6UVVVkHtNFkRhTFyQS0KONjo9idLvw+Lzq9PrOG7DHE6kxEEYu3QVdH23SbcFSsdgefuvMrfPPuT2eFIksyDv6jl+5TkSZHyiUxKrL5hWe59bN3s3MyajM00MfQQD/JRAK9wUXxRReQl1+Ib3yMDete5qXnf8zmDa/x+Xu/zcb1rxI6SvZpYVHmIVVJEoN9+w5JvU7E46jVGlRSjHxPEeVVtTz75KMAlJRVMuEbJ99TTEFRCUG/H+/YyCFZlgVFJciyTHllNalUisraejRabXaxa8j4KjzFpQwP9lNYVEIkFESj1bL8nPN48q9/yh7XPH8RBqMJw24T+Z4iTGYrGq2W0spqikvLiUTCBP1+NFodRaVljAwNku8pwjc+zubxAw7umYAiFjOU6z92K207t7PzJMbWuWY9Dm0u/UNh1rz5CG27dzM0sI9wMIgrLx+L1YreYGRsZJg9u3YwMjRIOn0gvX3TG+vo2dvBtR++hf958EdHvMb+9O9EIpOnkFdQmH1tf5q3KyePdDp1yLBMJUk0tCxg57bNWKx2vOOjtO/cTmlldTZatL88QCIRR6PVgZwpvnyw3yQSDjNn3gKG+vsoKC7FNzbK0EAfu7dvy0a5IONr6u/twe50sX3zRipr6+nu3INOr0dVWUMsGiWVSiKpJXq7OnG4cmnbvg2LzXbC7/vpzqx1cM5kTBYrv330Wb786Y+dULhVADyOjJN2jsfBroFMNGfIHyEcP7ECPHPmLuCe7z/ATVecRyQcPuz14rIKEok4arWWWCyCWq3JhpHLKmtQazSEAn7UGi3xeCy7Sr2nuBS1RsvI0ACyLKM3GLHYbIyPDOObTIJyF3iY8HnJLyzCP+FDlmUmvOPk5RfQN3kend6AKzePYCCz+LPeYCQSDhGYmDjER+Rw5SCKKlSShFabSQyLxWLI6TRanQ5JyvSIAv4JikrLGRsewusdw2gyz6ikLFEUo4iiGCEzWlW2GbJd+r7r5If//KQsiuIJt9VIotxYaJe/cOEc+eoFpXKhzSBLonDC51GpJPk3f39WPvfiy6f9/VC2t7+JohiZlXNDZjKCKHL+pVfwxF//eFIVtuLJNLIs0zEaYmOPj+GwTPIk5jmkUkmeeuRPnHfJFUes/aBw5qH4LGYYVpud8uo6Xrrz1hNuazA5yM8voazYQ6/sYlG5lvyghHe4B99oD6NDe4hHpx7iXPvMU9xwy6cxmsxHnWZ/0giTs84U3jWUnsUMY9nZ59K1pw2/7/BCLkfDYHJSv/AcPvDV81jygWYShUtwFtXiN1dhK6jAXdmCp2IuVQ3nYra6p3ze8dFRBvv7WHzWqpO4k0yy29FYsOQs6ua0nNR592M0mfEUZ9Lwj3a9/a8dD09JWXah7JmKIhYzCEEQWHHue1jzz8enOAQRcOZV0rLig5S3nIvFncRa3InGNIIgiCQSMdJyCI15H6VLvBTNMVLZcDZanXlK9qRSSdb+60nOPv9iJtNep4zeYJycdFd4xNdjsejbnozmLvAwPNSfnb4uyzKu3DxUqkyHW6vTHXXJxf35Gfux2R0nXaHsTEERixmE0WSmZcES3lj30pSOd+VX07jsfRgcLiKhNBufKKX12fmkYsXI6RQCAnrbCM5CHemUhsb3DGIvHaOsZjkq1ZHrfr6VN9a9xNxFS9G/pabnsbA7Xay64GL6e7tJxOPUNDQdvsyCnCnfl19YRFFJOa6cPOrmtKBWa6iorqOgqJi8gsJD6ngYTWbqm+dhsdqormtEbzSiUkm48wsxW22ZwjaiCkEUaFm4lMLiUiRJwnJQj8GVm0dOXj5anR6dXk9tYzMGowmNVkttYzNanZ6G5nkndL9nCopYzCBqGpqyhX6Ph1pjoG7RSnKrUtSfu5m8ms0YrTY0GieJeDSbN+EdDDM20IvW3EMskqD+3Bi5VTFKqpcxld5Cd2c70UiEiuraKd9HeVUN46MjWO0OLDY77kJP1kla4CnGZLbQ2b6L0opq7E4XZquVhpZ55LoLKCgqxuHKweHKpaFpHipJfch5JZVE49wFSGo1yDJ5BYX0du+lpLySaCSC1W6noXkeWzeux1NcSjwex13oyZ6jpLySsy+4GLVGg6ekjKLScnLzCygpr8JoMlNd30gkHD5iuPhMRxGLGYSnpAz/hI/UFMoB2l3FVC4dwdO0EZkw9rwcPI3jqLV6JEmDWqvH6AiRFjYgM07IKzLUnkf7Oid6hxeLw47OYD3udRLxOMGgn8LisinfhyCKuPLc6A0GDEYjWzesz84dcbhyiMdimC1WJEnKTPqTZURRxdjIMO7CIro725EkiQmf95BZvWqNBmdOLipRRdvOVlKpFGazFa1Oh5xOM9DXkw0WatQaAv4JBKCnsyN7jlx3Ad0d7RgMRopKylGrNURCIVo3bSAei6FWa9i7Z/eUF5A6k1CiITMInW5/bt2Rq1lnEQRc7jKMjhAancjoXjfe3mpEKTOxC0EklYwx1j9OMlGDkKggOLIXT72Io0BGbXDg75/A5ixiMOw7+nUmryUgoDuBlcxCgQDr2tagVqsJBQO4Czx4J5dD2LFtM1W1DcRjUXbvyCwFuXv7Vnr2dqDWaIjHYpOFlwMUl1UgqsT98/YwGE3ZBC+DwUgymaC7cw+u3DzGRoZxunIJBCaIxaIYzWY6du9EktTZYssA615cQyqZJBqNUFRSxmB/Hxqtlu7OPegNBlLpNIIokpuXP6MK9oIiFjOKdDo9OWvy2CFFvcGG0a5lrE8mHnXh7W1ATguk4ilANRmSjGNzC7hrQkR8+/D15+Ed3EVBbZj2N8bxDmswWXKOa5OcThMMBk6oeO1bHZd7du84cI+pFLsPWpNl//8Pmy0a45Bp5IVFJQQDATrbdmbrjOz/t2dv8MjnOAIHTw7rnJxev7/Xc3Dm50wTClCGITMKlUrCaDQd9ziN1oham0JSF5JOppAJYXD2gOgDZBAERE03JfN24SqOUFDXi634dUa79UQDIjrpAnI9500p2UoQBIxGE6rJqeDTRTQaIZ1OHbbWh8LUUXoWM4jMA3H8X/BYJEDEr0cQYgRHPWj0Qbx9erR6F+m0jCjIyKlihjs7QZYxOSTKmk2k4kG6NtSiM5hQa0TSU6wHmk6niRzUlZ8OxkaGGRsZnlYbznSUnsUMwjs2ilanQxCO/bFGI34iwQCDu+oJ+1NUr9yMpWANkeA4AgKynEaQTXi7z6N3Sz0TQ3GSiTROTxyENDqjjVjIRzRy/KxMURTRaLV4x44+JV7hzEARixnErtYtFBSVYHM4jnOkzMhAO2HfKBPDfqLBFPlVEjVnbyKZ3oEgqhBEEVHUkIo7CU3IBMZi9LelMJg8pFNJIhNj+MaPPy7PcefjdOXSvlOplH2mo4jFDGJ0ZIjBvl6a5y8+7rF+bz9R/zhabTkDbQbKWpxULFBjtEdJJePEI4GMT0LWYXY4kNMyJrseBC+BkX34RnsJB45fCWruomX07O3A551ZVaNmI4pYzCBSySRrn/lHZjXz4zgfE/EwA91bCY0PIamKiYaSvPlEmPB4HSpJg0qtJRYJEPBG2betjkRMQyKcg0rVxcRQN31dG4+7VoggCCxduZq1zzw1uTShwpmM4uCcYaz55+P85HePZFfOOhaDvduw2NxoLWkEjZ/eLfMxOzL5ECpJg6hSI8tpQuMBJga07H1dhXdggq6214nHjj/71GA00bJgCT/9wTffkXtTmF4UsZhhDA32Ew4FaWyZz4bjzBFJpRLs2bGWeGwho535WHLVhL0jpJJxErEwRlsOyXiM4Gg/vVvTjA6tY2yoY0qrjwG0LFzCyNAAo0oUYkagiMUMIxGP88K/nuTqD32UDete5ngJWol4mI6d/0ajNWIwOdDqLahUakRRJJ1OEY0EiIS8RMMTUxYJyAxB3nf9R1jz9BNTSj9XOANQyurNvK2gqET++783yg5XzrTZkOsukB97cZPsys2b9vdD2d7+ppTVm6EM7Otlx9ZNXP2hj02bDR/48MfZ+PqrSiLUTELpWczMrbKmXn5kzfpp+WUvLCqRH1mzXi4pr5z290HZ3plNFMXIrFwYeTbgHR/FbLWx4tz3sP7ltUet+PROo9Xp+Ow9/8lrL77Ai889/a5cU+HUIwhCUhmGzFBkWeb3D/8ElUrFbXffi1qjOeXX1Gp1fOYr3yTo9/PHX/33YYshK5zZKGIxg4lFo/zk+9+gpLySb9//C8yW4xerOVlsdgfff+g35OS6eejH3znpxZwVTl8UsZjhTHjH+cqnP8bY6Ag//cOjLF15Lg5XznEzPKeCIAg4c/JYtup8HvzDo/R27eXez31ixheuna0oyxfOEkSVipXnvofrb74V79go6195kddffoG+nq4TXoxIVKkoKiljycrVLFy2ErPFym//+35ee3HNSS1spHD6I4piVBGLWYbJbOHK6z7MslXnYbU52LDuRV5d+xw7tm7C75/gaAv3CIKAxWqjoXkeZ62+kHmLlzE2OsIrLzzLY3/+/ZSqTCmcuShiMYvRaLWUVdaweMU5zF24FJPZzNaNb5BKJjEYjZjMVhAyC/6Gg0E0Wi2NLQsI+H1sfP1VXn95LV0dbSTi8eNfTOGMRxELBQBUkkRxaQWNc+djNJmxWG0kJ1O0JUmNf8JL0O9n26YN7OvufNfCsAqnD6IoRgVJkgLJZPL4hRsVFBRmLZIkBUVBEJRguIKCwjERBEFWQqcKCgpTQhELBQWFKaGIhYKCwpRQxEJBQWFKKGKhoKAwJRSxUFBQmBKKWCgoKEwJRSwUFBSmhCIWCgoKU0IRCwUFhSmhiIWCgsKUUMRCQUFhSohkSn0rKCgoHBNJluXn1Gr1+dNtiIKCwumLLMvP/f8aVmdl1Pb+AwAAAABJRU5ErkJggg=="}
,{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)", "background-pattern":"" , "items": [{"x": -626,"y": 96,"w": 2749,"h": 510,"type":"text","text": "","text-data": "U29ubmVudW50ZXJnYW5n","font": "sacramento","color": "rgb(202, 222, 236)","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -656,"y": 602,"w": 2803,"h": 770, "type": "color", "background_color": "linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)", "border-radius": 0 }
,{"x": -611,"y": 599,"w": 2740,"h": 776,"type":"image", "image":"png", "image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuxdB3hURRedLemhhNB7hxBCQuiC0jsoTYqCKIgFFRW72LAgKKiAP0hRBAQUpAtIkSJIh9A7Um006SVt/3uSvTg83ia7SSDtvu973+6+N3PnzpnZwN7z7j0WJYcgIAgIAoKAICAICAKCgCCQDRFwOBwWTNtisThSM32yY9bd6ryIVzTAGe8cLzXDSd9kEDCsR8Ia88FrjbVP7bpnl4Vwsb9vQqrhkPBFIFyzCzQyT0FAEBAEBAFBQBAQBASBO4CA/G/yDoAqJgUBQUAQEAQEAUFAEBAEMg8CzoAs/l9syjwkF4BNIqALmyAsbHSCrIgzGyM5+5kHSfE0KyJgQgDhe8K/I/GKM4GM0w4hL7LiZpA5CQKCgCAgCAgCgoAgcBcQ4Ce/7sJQMoQgIAgIAoKAEYFcuYPyCCqeIVCkWIlSIWHhkXny5svvWU9pLQgIAkYEctIfIZyCTELAlc+0hIMzK5iouFPjpKXPYksQMEOAyTf8fuR9zO9ByHnRic/6fUsy2RmCtCAgCAgCgoAgIAgIAoKAICAICAKCgCAgCGQEBGrf27DpoJFfT1l34J8rC9btOjJqypzFPfo8218IDNerU79pq/uBVdSJiw4+J839ZV2lKlWrZ4Q1FR8EgcyIwP8mz1r02fipszOj72npM8oDaadCkFU/UzuW07aVXm104hWnZDqnFljpnyYIGPe74TN/N/T9y9ewn3HanSfvb76f8D2SQxAQBAQBQUAQEAQEAUFAEBAEBAFBQBAQBDIwAm8PGTEWAfe1+/++vHTLgT/xecqCVZu2Hr8Qv2rX8XNNWrfrlIHdTxfXatxzX8MtR/+NBbFTs16DxqXLVazUrG2HzjOWrd+5/uA/V8Mia9ROF8dkUEEgEyNgpeO3fX9dev+zr77NxNNIE9edAVoOyN4SbE2LgKsWAIZtJiyEtEiT1RMjqUXABUGhk3Y6oZeQNWFyurqeWvekvyAgCAgCgoAgIAgIAoKAICAICAKCgCAgCNwpBGx2ux2kRKfuvZ5E8P3NQZ+N4rHKVwoLn7Zo9VYQF03btH/wTvmQGe1OX7J2O07gp/vvHxAQOHvlln2zV2zea7XZUJJCDkFAEHATgXIVQ8NAnj7Y4/Gn3eySZZs5g68IuPIT4yATbgZlUztxFwFhfho9teYzdH/HMmWh05edpPdedN4sS4v3zmuKXnH6ok+GnpQ4JwgIAoKAICAICAKCgCAgCAgCgoAgIAgIAoJAVkLA28fXF5kBzdt27KLPy8/fP2D60nU71uz940LuPMF5s9KcUzqXciGVqyCo2vbBh3qa2UDGBe7Xb9qybUrHkH6CQHZEoF3XR3rjuwNNmOw4f33OJhkQN8mENM6wMH1qPSvg7yQmQDjYnaRDEL0WpDPYeeag18J0lqCzDJ1lnSfe4xruoQ23R1/YAIEBm7AtREZW2CwyB0FAEBAEBAFBQBAQBAQBQSAJBER0W7aHICAICALpgEBEjdp1fXz9/LZv2bBWH/7a1atXPnnn1X4BgTlydnq415Pp4FqGGzI0PLIGnDq4d/cOM+c2r1u98vy5s2cqV61eK8M5Lw4JAhkYgcoR1WreuH7t2gEX360M7PqddA0F9+Pp5ML7dzJAfrO4v1Pj4k7OK81tOwkEb3r1o9OfBshJZ0E6C9OZm85cdAY6zzzO+370ihMCzdHOE+/5OmygLfeDDdiCTdjOibGcY2JsOQQBQUAQEAQEAUFAEBAEBAFBIIshcEtpjSw2N5mOICAICAIZFoEwCq6fPf3P33//efKE0UkE4E//89efdRs2bTl+5KcfZdhJ3CXHgpyZJnF0mA0ZT9ef6NKm0cnjR36/Sy7JMIJAlkCgCmm/7N25fWtcbGxslphQ2k4iTZWCLRaXvEfCOCzAjWyOJNqm7QxTbw0PPoFsyOc0hc8ge/CKElB4Rak+b2Xzjldx0TnoPYDAnPH3HCQFDrxPbJdoD0eAsy1+q+A69ijsgRjBGDhOO6/zZ+dleREEBAFBQBAQBAQBQUAQEAQEgcyMgBAWmXn1xHdBQBDItAiUD6kcvmfHti2uJnBgz67tIiSdiM7FC+f/xWu+/AUKHdy7yzTL4uC+3Tsz7WYQxwWBdEAA+i9lyoeETvlm9PB0GD7DDWkkCYg4QFCdWQYOst8xv2n8NCVI7pijZJiyGkAugHxA9gPIhBgnVsAJhAI+g3iIVwEhVmX1t6igey3KFuBQ3pQkEX3eobxy+Kjzq2PVhc3x6sYx/B5hQppJDj3DBbbwGSTIDedY+Iysi2jy5wK9XrI0uWnjTk5fbAsCgoAgIAgIAoKAICAICAKCwB1GQAiLOwywmBcEBAFBwAyBCqFVIpYtmPOjK3QQpKeqUAgGZfvjMNWrAQjAbO2qXxZne0AEAEEgDRAIDa9WA0L1u6I2b0gDc1nVxN0oC5XhsSNCACQCiAmcyIq4KaBN76/SCZICZAWIijgVUNFLBTUiyiK/l/LOa1FWH6WuHXIov3JEXvg5EkiMmNMO5V+W8igqWdXFzRZ1dpFSdkqqiL0CO3o2nUXZ88Sp+Ot2FX8V15FNwQQGxsZvGfxbmYv8vE6v1+hMKDVFBIZkXmT43SUOCgKCgCAgCAgCgoAgIAgIArcjIISF7ApBQBAQBO4yAtCuKFaydFlXmgxwJ1fuoDxXLl+6eJddy5DD7YrasvHqlSuXa9/XqNmEUZ8PyZBOilOCQCZDgDO4dkZtEsLCZO0MGReZJvshLbehUx8CBAXKM4GkIOYhgUwAYYDfEMh2ADmQWArKt7S3Cm5sUQFhRDIE2YisIDpjP1EZOS0qV13qVYAIiTMOqn8VrwJr2JVvGS8iIhyqwMMWVXqgVV0/6FD/rqOaWN5EWsRalYWG9i0ep2LP2lX0P7HKv7Sd7nmpuKsOdX6lQ8U7iOxYb1ex57lkFMgOaF/Ar+vk/xV6vUbEhRyCgCAgCAgCgoAgIAgIAoKAIJCJEBDCIhMtlrgqCAgCWQOB0uXKh1jpOOCivBHuVQgNi9i/e8e2tJixzW6339e4RZu9O7dtMdPMSIsx7qSN2NiYmHWrli1u0Kz1A7lI0OLCv+fO3snxxLYgkB0QgH7F2TOn/vnr5Ilj2WG+MsfkEaAAP+tFgIDAe7xCBBuvOHGAsABxAU0JvEe7eBXc1qZ8giwqMNyqvINtKvbqDeWV065yVrUqn6JWZUMShj1eWaoSqeCwKEd0vPIuTjZhwkrX4igDo1S0CqxlV44bFnVxS6zyKWRT8dFEcBSJV45Y7wQCJPYSNf3XoQo+RPkcF/xV7jpKXSCS4+IWGvPsdeWIhz8gV0BigLy4SPNCpgX8xSsyL0SzJfntIC0EAUFAEBAEBAFBQBAQBASBdEOAf3ykmwMysCAgCAgC2Q2B0lQ3PiYmOvr40cMHzeZer1GzVsH5ChRcPG/m92mBzcBhoyd8Nn7q7JfeGfRZWthLDxuL5v44DcRLg6at7k+P8WXM1CFQLqRyldRZkN5pjUDlqtVrIXspre16Yk/2hSdo3bm2FNC30AliIpjOPM6TNSpQ5okzTPAKIoCzKvyUPYddFX/JroKb2FT+LjYq/0REQ4l4lbOmXXkVorJPVR3KVjhOeRW8przyOpTdK17ZKYPCK9BK768ru280fY5Vdj9qn9db+Ze5QWWiLqjc91ylVyI9gmOVb1GUjiK+Iw9pYBQiD0palF8FK51eKiDCVwU39FJFn6bUxIZ+1J6Bgq/wHeWiMBeeVzDmijnfOUTFsiAgCAgCgoAgIAgIAoKAICAIpAYBISxSg570FQQEAUEgBQhA6PbIwf1742Jjb3vKM4CEK15+d/DnJ48dOTz3h+8mpMD8bV3y5M2XHxePHD6wLy3spYeN1b8sXnCJhD3aPvhQz/QYX8ZMOQKtO3Tp/v3Pa6Lsdi+UkZEjAyBQsEjR4sF58xfYvS39CAvZFxlgI5ALFLgPohecxAQkHKxRAWFtfGcR7McrUiH0ID8RDzmuq9KDAlXsBSoHVZxIhVCr8i8Vq/zK3yAy4TJlTFDPHCSw7Yt+sAs7/NuDRbRxDWMxCYIMiZzKj8pF+ZCmdq5aRFxERFN2xVUqH3VdxZwlEoKyM6yURGGJpawO0rew5XOooCZEWjzqrYr191H+5WFb9x32kXUBH3BgrkHOuWeMhRAvBAFBQBAQBAQBQUAQEAQEAUHgJgJSEko2gyAgCAgCdxmBkLCISDP9Cohsj5g446cChQoXfbR9s3rIwkgL117q81CHAoWKFKWEDiomnjmP6BvXr//047RJ3Xo91a90uYqVfj+4b0/mnEn287p1x249IJyO0l7Zb/YZc8YQ3IZnu7ZtTrcMC9kX6bs3KFiPGk0soo2APg4mJ/BdxW8EEA0QssYrAv64nqhXEdzcqoJaBKicdawqR6QXlYIiG7ZolbNogLLaQBhA9wKv0JNI7JN44BWfYRP/xoFYwHuMxxkcaAOf0JdEu8mulUgJa27Sq/jnqrpxCr77Kp9i1MbLrnIVpN7gIuIdKlcDyrwoY1eXtlxX/3wfrW6cYL0NncSAH/AvjnDAdZSJgoC3HIKAICAICAKCgCAgCAgCgoAgkAEQkAyLDLAI4oIgIAhkHwRIyNVSqUrV6vv37Nyuz7oOCUr/sGTttkphEdVe7N2tHfQm0gqVa1evXsnMZAXjMGPy11/hfeeej/dNK2zEzp1FAFkV1WrXrR+1ce3qOzuSWPcEgdDwyBoOOnZv37rJk35p1Vb2RVoh6ZkdZ+mnPPSKrDsulQRyAJoUTCgggA+ygDMscA8HMiwSdSCgNVHyDS9VqLONMipIt6KGTdkDSGjb14fIBZAP6MvZGExEwD5OJipgk7OumKDQ++I9iAn4CS0KP2Xz8iE9DF+VM5I8LkFZF5Qo4RVE4tuXSRvDRkLelOFhJx2NuCvxqmAXH1X+80DS1iCffOEDfOLSVvqcE0pfARM6gY2UivJsW0lrQUAQEAQEAUFAEBAEBAFBIM0REMIizSEVg4KAICAIuEagWMnSZXPmyh105tTff4VXr3XPo0+/8OqUBas2jZoyZ/E/f/1xslvL+6qtXfXLYk8whLYDiBCzPigHVbJs+Yqu7EHgOx+ldHgyXnq1PXJo/97N61avbENP7Pv5++Pp2Cx5ZKXSScVLlSnn7e3js8vD0kPJYYDSaVly8e/SpEKJND1+5PBBqrL2rztDJrce7tjQ26R0X3g6jrT/DwEKxCNgn5tOEABcnglkBDIncA9BfSYXOLCP7Ar9vVL5O15XVebmUoFV7VSKKVp55SH9CdKlUOoynSA1cKIfv4cTeI8DGRXX6GSigsW8OcODiQ7ch29cQgrX8ZmFtEkDI6cPjU1lqaialW95KwluxyqHFeLcDpW/vV35FKQMkIZ2VfZ9i4pY7KPytiXh74R/NnieXCaKxwEmwCa3EyvZPoKAICAICAKCgCAgCAgCgoAgkE4ICGGRTsDLsIKAIJC9EACpMGne8vUzlq3fiZkPGvn1lG9nL/3t+TffH1KkWIlSE/732eB+PR9sg6C8u8iUrVCpMoiODQdPXVux4+gZZGkY+77zyZfjJ8xcvBrjm9nt3LPPMz/9tv2wTniAVPlk9MTpq3YdPzdn1db9VWvUqcd9Ubbq2Vff+ejnjXtP/LR25+8hYeH0qOvdO2ZOmTAWweoWDzzYzd1R72nQpMXQsd/NBPajp85dUqVazTpmfa02m+21D4aOvK9Jizb6/cYt7++A/ihH5WpMlNz64PMxExGI5TbA/LG+L74GLOFDUv5i7Mee6f/6ks37/9hw+PR1iKR7eXkjOHfLUbNu/UZvDR4+BiQA38idJzjva+9/OsI4vt6xxj33NRzw8RcJGSquDv+AgEAz4svTMcNIzPnLSTMXDp8wff7bQ0aMxXj3P/jwo0PHTP7x068mzRj42egJ0HEx86NRi7btpy9dt2PTkbPRM5dv3A2tBWM7YLx8+++n6jZs2hL3gN0jT/Z7edLcX9Z9M2vx6vouhNmxRvBn8aZ9J1fvOXl+3PQFK5544fV33CG/8F0DvuNnLFzZpHW7Tq4wTM0e0m22at/5Yfy9WLP3z4sL1+0+in1Zr1GzVu7u+aTaJWR5hUdWd4dEcmc93PU7NfsiLeadXW0g+E4ngvEF6ERAnvUiQFSA6MbfGZASiWWZbJQpERhhTSj5VPpDu6o0waLKj7Cp8Pneqs4hb1VpWg4VGEZEQU7SjkjQpeHsBbAB+F2BzyzMjYwMkBScXcElqLgkFC8LkyL6MultdEIF7zFWIrlhtccqL0rE8A8l33NalIX8d1go44IyLSx03bcUERWkoVFqgLcq/Z6X8i3Cpa64/BSXu4KfsAmMCgAzIS6y67dG5i0ICAKCgCAgCAgCgoAgkN4ICGGR3isg4wsCgkC2QAAC25PHjhy2f/fObX//efLEiMHvvTH2i8HvT580btSx3w8d6PnU868s23rwr35vDBzs4+vHwqAusale594Gk+ev2FCydLkKU78ZPfw61X168+MvRhs7nP7nrz8R0A508UR6lciatWNILAPlYdAXwfxpi1ZvadC89QPQHUBwePCoCd8jeF6xcnjVGUvX73igS/fHNq9bszJf/gKFnn/j/SF3cwGXL5o/68K/58526t7ryeTGRfAYAer/TZ61qFqtuvedO33qH5TCGfXdnMV58xdkgdmbZhBQ7froE8+279bzcb7Y+ZE+fUFWgLR4deAnw5u2af+g2bhtOnV7BOe9jZu3xn0EhQeNGD8F64k+wyf8MM9VJgueXv9s3JRZz7327qCojevWLF0we0bD5m3aNbu/QxfjWCA1Oj782BOlylUIwT1K1skDQqrrY08+h/E//3raHDP/kMlTqEix24L/3BZru2TzgT/MguKejlkhtEoESCVosJCuc0FoV2BPFy1RqkyJMuUqYM/SlG8T4IaPwwiHa1euXP5+wpiRaP/ki2+8a5xPuYqhYSBssGfJrP/oKXOWvPjWh58GUTYRMgce7NH7KWMf7GsQIcB13owp344a+uE7IDCefunNgf4BOVASxuXRiexNXfTrFuBbrXa9+m98OOx/rhqnZg/BJvbsRyPGf4cT+3wk/Z1Ys2LxQuxLV0RMct8D4318p0E8Jqdf4e56uOt3SveFp/OT9v8hQAF3fM+QjRRMJxOgHKDH3/w45V3YrnJEOFTpgbGqeP94Veotqyrc3aqK9fNWuWvblHfpWJX/QbvKSzyuPwlh27wQ1EfGBGdFwB5OLikFnQu9rBSXlmKtCiYiOCvQjKzAJNgeZ11wPyZX0B/X2K5N2exUlsp+XXkjkcQapxzxcSrmPJWwKmdVPsWJiKmqVJnBFlXiZSI5gnkOeGUBcPYJWAGznE4MZVsJAoKAICAICAKCgCAgCAgCgoAgIAgIAoKAIJA1EZi9csu+94aN+sY4u0JFi5XAk+dRJy46QETkCsqDYInpUbho8ZLIfpi+ZO12BKzRCAFr9EW5Kb0TnrxfFnXob1e2YGPe6m0HcT84X4GCaIsTQWFcw1PesIsn5PG098dffjMVT+LjHkpZIQh8t1fqlfeGfAGfyoVUrpLU2Ahio907n4wch8A22pLgeTVcwxP5xr7d+zzzIu71eOK5l3AP5MbmI+dikO3Qst2DD209fiEegWSzMb/45vu56Av7uM+2nur/xnsgLXBPJ0J0Gy+/O/hz/T7IjpWUMQOCRG+H68gM+HX3iX85YwYExW/7/rrUukOX7v/7bvbPsIMMGb0fCJG1+/++7CpDBGXBsI5bjp2PK1i4aLG0GJNtjJk2b9nUhb9uTm6PNGjW+gH4jiwG+IP2IIqwP419sf4bfz9zI4BYOOC+5ei/sQ8/3vcF4INsCSPhhwwm4PbD4t+2YY+zPWRLIIMoKd9A1sCv+b/tOAwyp1nbDp3xGfuA95TePzV7CHaw5thnIMrYLshJjNnigU5uZxUlNSdkb8AeyBVX7TxZj5T47e6+SG7fyH3XCFCg3U5nETpLOM8y9FqKzpCEzytzhzh2PlTRcXRIiGN//1DH8eHhjpNfhTqu7Al1XFhd2XH1eCVHXGw4xfxDiRsMd54R9IoTn/m1ivM9XsMM79FXb89tKzuvR9IrzqrOV/7Mr2jv6p7uC9rx+JWc/oWR7xGO2OhwR/SNqo6Y6EhH9IUIR8zlSMfFrVUdJ0eFOTaElyUscCZikvgKjIAV4wYMTTMUZf8JAoKAICAICAKCgCAgCAgCgsCdQUAyLO4MrmJVEBAEBIHbEEjQk6AnzLdtWv+b8eZfJ08ce7f/04+9+nTPzhVCwyKGf/PDPLOSQOj31pARYxCEhjg3laA/h2sUj08IyMdRKoduGwH03dvMhXUR9MYT73+eOHYUfV57/5MRIEBe7NX1gYP7dieUruLa9W8NGT5m8bwfv3/zud4PX6Un4HGPgtvFz54+5ZIM8XQLoGxRjz7P9k+u3+L5M39AGwReXbW9p37j5iAe5s+YOvH9V5/rc/3atatoCzFz+I+MAmPfipUjEspbrVj80xzOzqAkkx2vPf1ol0VzZkz9648Txyjebar3QfYikTkD+yhj1Pfltz/4/tuxX3712cfvzZg8PiHzxSzDAjomD/V++nlk2syeNnE82nHmQKxhLYsUL1kaT8b/uuznn5Cx07jVAx0RWH6n/1OPLpj1w3c/z50xzWycSuFVqyOQv3PrpvVmeCEQDoJqHWmnYA56m5SOyTYqhkVEkrBzkoQFTSk3MmH2796xDWsVTwfv6VgCwehzrXsbNNm+ecPaNh0feuS+Ji3bDni+T48p40d9AdwgMH+DFpv7gMQAQUhJHjF9u3docfb0Pwn7FXgg62LV0oXzXO0h4NLv9fc+3hm1eUP31vVrrFm+ZCF/30Bg+Tq/c3r/1OwhlN4C8fj1l0MHYT+w3dr3NmwaHxcXh/GT+264c79SlcjqyHrZv2fXbWQQ+nu6Hinx25194c5cpM3tCDiFtZE1lBd/TpwnGnL5p3hVqIdFFX3WpnLfZ1VWH4vKVTtW5b43TuVuQO29Y1XOepeUH3GXVluMslg5WM8ZDbpeErIfWEibr+M7i3H1kk7IYkA7/t3B2hQ3v6ou1pLLN3G2hd5M17/gdrj/X3krC2VZ2LxIZ8ObSlh50Vz8qFxUbByVhSKdiwdtlG3hp4LqAxrYR2YIXpFdoWd/wF5ewjWHCHLLN04QEAQEAUFAEBAEBAFBQBC4OwgIYXF3cJZRBAFBQBBQrAWxY8vGda7gWPrT7BkD+vXpjkB27+deetPYDsFLaFWMGz7kA4qfH+H7FSpXqfrnyeNHr1y+fImvgWyAxoSrQHVxYk9QWmff7h1RkVQyCaWLxg3/9EMEaGEDT7oXL5X4tD6uDRrQvy+XjkIGCAiYk0d/P5wWS4tSSv/7btbPSQmE8ziYDwLrqK9vNjbm/TZlVQCPQQNevPmkOre9euXSJc5M0ftXJAxRnuvksSOHO1BZKOgWvEtkAEoboR3xO7eVMcL1oOC8xEUUKfrbiqWL8PkF0iU5R0zOFx+9/Wpiv9vLH/G4L7z5wSf/nj1zevigd17ja8AAWQIH9+66JXuFSZY1yxcvBJn10tuDhoFE+mXh3JlJjRNerdY9CHiDfDHiBWKmz/OvvY3r0Acx3k/pmLCD0kPI+HG1/3gslEPDXvrojReeYqxBppWtWCns4L5bMUB5M+hf/H5w357nXn930Lejv/jk57k/JhA1ZgcyFZChMPjtV55jsgLtEGQHhpvW/rrCrB+IvveG/u/rQxTVf6Z7+xZMVLTt2O0RtN+zI2rz+XNnz9yOV8r2EAiUd53jjf18yPu63XsaNG2xd9f2rZcvXbzgap6eXEfm0MG9e3ZG37gOYeTbDk/WIyV+u7svPJmTtE1EgALq+H89SkChJhJ0bljrBoF4rHesKtTLpnJG+pMOhVUFVraRxoNDOa7EK1uOa8qn0GUq+4SAPTL1WJuCSz7xbwZ85jJNXPoJ10BK4JVLPDGRASKAbcFNJjJYiNud5dNJEm5vLCXFdjHeDTpBXLKwduIc7F4OZfWnfrlBzBBSNWyqwtgAVbinXdlzQdMDNkG4ACsmSRhHYIoSUfLbyZ0VkzaCgCAgCAgCgoAgIAgIAoJAKhCQ/3SnAjzpKggIAoKAJwhEkHj1RYp8JiesDdICZ8+nXniFyy/xOI889fzLCJROoxr/fA0B7iYtH+j4049TJ+n+IADv7ePru2OrOUFSpkKi8PG+XdujoJ9w/MjhgxD/ZhtUc74qtAiQnfAWPcWOp/r5HrIh8H7blg1rPcHArC1KO0GM+ZeF82YiaJ2cPZAm61evWIrAp7GEEfoi8wLXvxwycABnVug2/fwDA28YgrXAqVSZ8hURwAaJ0/u5lwcgQ4IzTRDcJlqiIHQFjP6VrxQWjmub1q5eAZKjaZsOnYe+9/qL/KQ/a0cY++IJ/4gatetO/Gr4p5y1Ajt9+r361hWKTq9cvGCuPhYyb3gclJdC8H7Y+wMSylfhIM4kQaPCOE44jQMixixAjVJSyPpBMHz1L4sXGOeW0jFhByQYXrcnsUdAzJDwe1+MzUQZ+qAEWf6ChYv89OO0W/Z05YhqNXEfmRXECf3z1bBBt2lc8BywZn1eePXttZQ5AmJHnxtE0JHJgUwN45xBsqDUVnR09I1+jz7YhqA5jzZUia00l2XauGblL8Z+qdlDHR56tA9KvX3wWr8nmLSB/WASAcH3GNomxvFS8hkEFUioPTvMs148XY+U+O3OvkjJ3LJ7Hwqk4wBZAQ0k1o1A0D1Rn8G7YA6V934f5VPAQpkVpE1BVQfjr8Uprzw3VAHi4fzL+pCQNogK1qZAP12gWicI8G+BnvXAWQ0gIXCPCQb2Q8+6YDv4DeJKv8K4nGaEhX4tUY8jkagA8QC/mazhe4m/eWxeNGdkXARSf4LqxokYFRBhUQW7WJUlQeYDxDTKHjKBgXniGuYCbEFayCEICDU2E84AACAASURBVAKCgCAgCAgCgoAgIAgIAncQASEs7iC4YloQEAQEAR2BqjXr1NtFmQqcpZAUOjOnfjsWNfJr1WvYhNshgFurXoMmKB3EwXDU54eo9LEjhw7gaXPdJgLieLLelbhu2QohlROiM97e3gic4yl/PVjaoFmr+3F/0pjhQ1GySreNkkv4HLVh7erUrHKiyPC470CWoCQWlwNKziaPi1JMxrY9n37+Ffi75KfZ0433oHuA0xjUBxbwBeTO/Z0ffpSImhwQRef+EIDG/RNHfz9ktFmhUiKRsGPrhnWP93t5QNTGtatXLvmPbChBItO4f+Lo4Vv6IigPEoFLQaENRKZBuHz67msvcKCcx6tQqUoEskbOU0rGY8+8+DrWBaLqfB/jYG9R4s0tWS8oAcTEi+47Mj+e6v/me7i2/tflS1Em6Pa5pWxM2Imsec+9586cPgWyxNV6Nmzeuh1KEH0/4aubBBzIhNc/HPolynkZMyCYHAIhNXLIwDeJU0CA0vRo/kDHrgj4TzR8L9C4bsNmLSEqb8QY95597Z2PkDED8kDf931eeO1t1g7ZYVJeK6V7CGWruvR84pmttG+M2Sj3NGzSAve3bUobwqJMuYqV8HcFGSJmoHmyHin12519kdz3X+6bIgA9owA6EajnAHtiloPFy6rytY1XOcKp7NO9VhV3I0Z5F6H6X1Xpcz0blX3Cdx+ZZGjPItQgGThrAuQAkw4YHIQAZzRwWSi88skloZi84IwM9OUyVS6/u9rs2JfklpwzPUAyYEyULUSWBEoB4jPmh5PLWkXTnIm4oEqKuer7qHzNrKpQby9VtC9hQaLdiVjw/IAJEy/AFhgnaEfJIQgIAoKAICAICAKCgCAgCAgCdwYBISzuDK5iVRAQBASBWxDAU/t4Wn17EuWg9A4H9uxMqC8PMW6+jtr9KNMEvQIETjs+/NgTPyxZuw33+z7cvjnq9+s2QFgcoLJC+tP7+n0Ef//564+TTVu3fxABzOU/z5+t329+f6euyFCY+s1XI/TrCNxDOwFBcATQU7PUjVve3wH6CeNGfPphUsFn4xgoCYRryLLQ76GUT2kKys6cOmEsyBpjv7JOMfHfDyT254OySRJIh707tm15+PFnXgT5g2wYvs/ZKL8f2r/XaBN9UdYJ15u0atdpxOD33tDblKlQMSGTxdi3Tv3GzaBHgaA5hLJBPEGke9SnH749d/p3E24fJyxi97Ytm5q1ad8ZmiWTx44cdus4IaFYDz2TAhk60NQgt3cZ7T3QpftjeKof111lQWDPejomjwMSLCqZQDswOHvm1D/r16xcBuKi/zuDho2c+OOCTb/9uhx6FkafWQz+6OGD+7kUlqv91+2xp55DWa2Nv61arrdBRhKIPrPsCuyfjg/3ehKZHchy4n7InGnToWsPztihrKStZvsgJXsIYt5Y/6mkw2G0Wbdh05a4ts0kE8TVvJO6zqLwrggLT9YjpX67sy9SMrfs3Iee+NczK5gcQHAe2kbxyjt/vPIpaFNeBezKr4xNOSgG71eOAvbB+B2A9ih3BN0LHJwtAdKD9St0/QmGmss/MTnBvynwGe0R9IdtzsbQyRCQB6wVwRkQPDb+brOeBPpwf1fZGLpeBmdBYC6cEcilqZhYgX0u7+dQNpqidzmH8i3hpQr38VGl3/NX+Tt5KXsQ+uEEhlwWiwkZPyfm2XnbydwFAUFAEBAEBAFBQBAQBASBO4aAEBZ3DFoxLAgIAoLAfwhAYwJPtO/YssGlfoWOl9ViTfj7fFXTpEApFQR3USJm7q9RB94aPHzM2pXLFndrUS8SxIMR7ypVa9amQOdtAt/crkpkjdrnzpw5hcDj6GEf3VJaB2RHidJly0OA2piNAE0A6DboWQQpXevmbTt0gf0VP/80xxMbZ5ziySjfo/er16h5K3x2FcyufW+jprhPQtCb9H7lqSwVslaQSQF9C/2Jf7QDCYLXAyZCxeVCQqvs37NzGwLkKFVl1ChBX5ASf/9x8jiPiQwBkAXIPvjg8zET56zcsq9SlarV+z/+UPtxIz750IgFfEKGDcYhMfH+IFR0vRIQWCBvmOji/hgbT8If+/3gft0m9mKvZ196A3oduG6WMZDSMWEPGicIwm83EZjX/cCe3hW1ZSPKYC3asOdYNxKdHvP54IH9Huvc1izjg4ijhKygH74d82VSmUoYG3jO/n7S10Ys723UvDWuGUka4PTmoM9HUdLG9eEfv/u63u+ldz/+DNlH61cvX4ryWUZxcrRN6R5q8cCD3VDmbYWWlQN7WKM69zVuBq0aXX/Dk++JsS0RFpGYx6F9e24jsNDWk/VIid/u7ovUzDE79YWeAp2Fac4I0CO7AMF41ibhgLtNlR/qpfJ1oFJQdeKoNFS0yl3XQoLarEWBgD+yHdCPg/8gGzirgskKzrZgiJnY4GC+nuXA15DpAFsg03kMvOq/P9gO22WSAqSFTjqj3W1ZYE4/9WXnUlHIhADhAi0LZFrghD1cw+t/BIuNsiq8CxCCJWJV/s6KiAuLKvORnbJPQKowjhgDGKEvsIYId2HRtNChl/eCgCAgCAgCgoAgIAgIAoJA2iDAT06ljTWxIggIAoKAIGCKAIRuEWDdtW3LRncgKlws8cn3U1rJn4jqteuixM2Hw8dNRvkYlFDasn7NKjN7efMXLITsjG0uAsYIlgeTJkMQqR2TrnHUmuVLFup22nXp0Qufl8yfdVtZJTzhj3vQnHBnLkm1CSVNAmSBmAWnk+rnSxkGuB9D0Ve9HfQaUCYJT+Cb9ccT6xBQ3m7Q9ShfqXI4xfT3dH30iWcnj/vyM2NWCslbhCLQe+TgrRkW0EkoRU/s42n9dl0f6f1Mjw4JT8TrB0SijURCOK0l2pBWxpsIgH/95dBBE78aMRTaFWZ+cykkaIpg7X6YOPZ/ejsIqMMX4zhFipUshXYouXXL+nbt0Ss3sU7zf5wyEToE+3benjGQ0jExDsgwvG7bvN4lYYb9B10InPVoXX6eN/P7r4g4oySR380wQAAfWGMdFs2ZMTWp/cGZCWakWst2nR9CX2OGBYTfoZExfuSnH5059fdfbL9h8zbtIHaP6yC8jHuA26VkD4EkqUslsFYtWzTfmBFUl8pBgZAzfjdT850rTxkzh/bt3WX2ffNkPVLqtzv7IjXzy059KVCOp/3z04lsAdaqwHsE1DkwH61KDvBSMZetKoYSxnLWu0oaDgjU44QeA4L7CL7jFTYQ1Mc9tsNZFFwWiQP9TEjokOuC27iODAecrFWBv9U4Qa6wj+iDsfS+aM/30R5lmHANfnLGBttkvQ3j0rOfaAfigkkTzijhDAsmYxIxsAfEK2tpq7p2mMpo2S0qX3ubir0Yry7vwO8lzMVY8gr2CtBanLI0uYVcMfrj9mf6b4IRx4S+9J1z24Y0FAQEAUFAEBAEBAFBQBAQBDI7ApJhkdlXUPwXBASBTIFA5YjqNY9REB3BaXccRpAUJZL0mvaoq4/MgB5tG9bq3bHFfa7ICtgPr17rHrxudxEwDousmRBQRnmnb/437GPdJ9S4b9a2Q2cE7SFYrN/Dk/wo44Sg8v7dOxLKUaXmIL4k/znKGvHUBsW4y6KPMbME5X5AwJjZA3EQVrV6LWSN6ALiaItSURQP9w6pUrXadAMZgPsoCXV4/97dusYHrmM8BNJBlOzduW2rUYMAwtiY414DIVCgUOGi6P/ZBwNebl6jQtFRQz96xxVZkehfpTC8IrA/5evRw43lv7hklXEc4q2oUL1Sf/1x4mZ2B8Sh+zz/6tvIIkGmx/7dO7eZleNK6ZgYL4wIC2AF267WljFYMPP7yW3qVSkDYXdXZAVslC5fsRKw3rB65TKQTkntmfBqtepAf8KovYI9UKZ8hUrIaDDqkVDmykso+TSJiCO2jfUbMPiLr+DXxNHDP6WElTBkPJiNnZI9hKwYZB1sWXc78disbccuIDl3bt243tPvh1l7kAyktxK+f4/599aT9Uip3+7si7SYa1a34SQrWEeBtRb4//TICkAAPkZZ/b1VYGW7ylUrWgU1vE5kBYheBN3RhoP+CO4joM8aDwwfZz5wkJ8/JyWUrWdbgAxAWT38m4cxkOmA8fGeNSFAHHDmhF5KCmOy2DXaw1/Ws2A/uMST2XKDYOAx0BfkjF7yigke9GUcEjNOrLY4FdyCMi06EMFT01sFVPJR/hU4qyJBldvZh/Uw8DmPc03MfPHoGn1NHSAnjKdHRqSxICAICAKCgCAgCAgCgoAgkMkREMIiky+guC8ICAKZAwFkWOyI2uRW4BHlltp36/k4nqxmUWBoYFBSQQBEiN3J0kAAHWVrzErXADHcxyuCr8sXzZulowh9CjzJ/ys99a3rIaANykEhiGvsk9JVQIA4KDgfnhL26ECpHHQwll/Kl79AIf3peN1op+69nsTnHyd//ZV+HaWW8CQ79BFwTy+1hHYIkqM8lpluAQLYaFOOSkp9O+rzIcZJIECOa/t2bbtF84AqPAXj+vRJ40e50hjRbbF2Q9ESpcugHJLrcW7NlMhDgICc0ct6de/zzIsQFZ9EGhgQ8jYTEk+Yk1Pvw9Mx0RflkUDwJKVLwhgsmjtjml4uy9VGqBhapSruGbVWzNqDbEHmjvFe556P9z1NaUs7ozZv0O8hG6la7Xr1l/w0a7ouxI2yayiN9cYzj3Wj5KaCPsTm/Xni2FGj3ZTuIdZUOUgsm24TRFIICcqDZDAr1+XRl8XZGJk5+F4fIu0Zs/6erEdK/XZnX6RkbtmwT6BzznhlAkJ/vUFkhUMV7OlQuRvZVWDCnykO+COYz6WOOAsCZZpw6qWSOHuByzJxZgYH+I2w60QGZ3Dj7xx8ZPIBRAoyJjhTgn3isUBq4ODSS/jMgtnsG/dFO1e/Y9iero/BmhzIIoF9PbtDLz0Fm9dJ3+OG8i4Up4o9a1V5mluVX2n4YYa1vhap3orEUSpkWThf8T7hlEMQEAQEAUFAEBAEBAFBQBDITggIYZGdVlvmKggIAumCAJ6wp4o9FTavW70yOQdQ1mfgsNETQE6M1MSbc1I0EX1jKOsiORu4T0+Y3+NKSBn38aQzXudMm/R1PB26zUYt2rbH52UL5vxoHKtB01b349qqpYvmu+NHcm1QXgfkCcVRcyXXlu8jgNymU7dHiECIYvFt3ENw14uIHWP2Ae4hAIySTSgDZNSv4EwClMmZNmHMSKMfeJocpMWh/bfX/efALe6t+3X5EmNfJiyMoteeriePM2/Gd9/qYuA8HkpWIXvHmHEC0W3SYkcd+YQDpcJ6PfPSG+NHfPoRyCgIcpvpn6BtSsdEX2hnoMRWUmv6HwbRbu3pipXDEwgL0m35Obm9UqhI8RKniAXR2yEbpnxIWDj2mpGwqNeweSvsH11Lpc/zr72NbKIvh7w/ACQhC7z//ecfJ4zjp3QPFSb1b9iiKma3+Prc6+99zALqZropyc3f7D4yVHAdRJLZfU/WI6V+u7MvUjK37NSHnuRHgBwi2xDKRtAd5AMC6fg/vV35h9hVoV4xqtSb3qrIE/HKnvBPByLeyDLQsyv47z6TCWgDMgFkA06uQaSLeDPUZvWJ9GuwBYKASyiBqNBFtnURb7RlYgE2ztB5ic6zdIKwYG0MngdIFl3wm68bt4GeeZKITaIP8AWEBWwzUcFlp+Av2iWUHFQ+xalHoWiVv6O3KvhQjPIvw9hw1gnPCWuR07k2Rj88+qyVfpIaUB4hJ40FAUFAEBAEBAFBQBAQBLISAkJYZKXVlLkIAoJAhkQAWQlwDKVsknIQmRUjJs74CfX3Px7w0jO6DsPVK5cQwFF4wju5SYL0qBgWHmnMPuB+IEPw9DY+/zzvx+91ewjM39OgSXNkPqxZsXSRcax6VOcfpYuSIkOS80+//9PMaZMwp/5vf3SzDE9S/RFUfuOjYf9D0HnsF0Pe19uifM6/Z8+cBkFktEH2h6HU1QiDmDLala1QKUHIGcFqs+wMLrf0+4F9twXgue+MSV+PNvO7TIWKoSCEjhw6sE+/TxyCcz19k11PzJmJj+kTx48yHyck1Mw/lH+CmDj3ef3DoV+iBNeU8aO+YH0LM8IiNWNiLGQs6ELReLKfNTHYF08wQJ8KpL8ALQ5XBIuOC4ia2JjYWwR6X3l38Ocb1qxYBsJrh1PDBCXR0K9SeNXqeGUio2W7Bx96+qU3B/5C2UeTxiSWiCpAk8Lr5UsXbivrltI95E+ZLrBJXNlNXyF4Dz2Ma5R6Q9WbtrDeBPvqyfdLb1uASDt8Pkab0cyGJ+uRUr/d2RcpnV926EcBcQTGg+jkEknn6T3KOcUqe+6rKkdkrPIvHa1yRpDyfR0KsFe0KltCsgMC8ExCcNkm7P3EvomkANpwIJ4D+bpWhVFb4Rai24k/X2NBby5BBfICRAvEt3UChMfnrAeMi+8E/i5iriAX4BO+cyx+zUSIMe1AL/PE24GD/vzK5AdsYwzj7yC9fRyV0LIpr4IkVB4M0sJHlXydepXCdxXzAG7wH2vAZauCnGuU2u0oKRWpRVD6CwKCgCAgCAgCgoAgIAhkagSEsMjUyyfOCwKCQEZFQA+a16hzb0PUwD9Fj2ab+Qux20effuHVeau3HQyrWqN2/8cfaj93+ncT9LYoG4RgOj/1zvcCAgNzPPZM/9fRn6+FRkTWQAkp41PkfL9qjTr1oEWBp8ZPHjtyWB8HgVIEl9euWrZYD3SjDYvyQqvBqAGR0nWYNfXbcdDiQAmsdz4ZOQ7zcWULc3rzo89GNb+/U1eILkOLwtgWZZtq1WvQBOQE33ugc/fHmrZp/+DMKRPGQqzc2IcJidnTJo43GxvZC7hO8N+2fugLnBbO/mGKed+Q0Iukt2AsrXXs98SgsXE9sTYffD5mIjIf2B7eIwAPAkrPKOH7IJnw9L/Z/rpO6RXcDoLiyBgY9v6bL0FfgjgfBO3UKcPT/biWmjGtOCxWq59/QEKpFOyncdMXLMf66hixELgRA0o6KPXqwE+Gs3A290G7vTujtriz15CFwsL1aP/4c68MAMmFNQSBtCtq0wZk6fy298+LKH1FFbryot15Yrxw/cMvxk7CXoKuBogw3PP28cZT2IoD+7ofKd1DF86fS9DiKFysREm85iMhicFfTpj2+YdvvQLiAsQgNC7Gz1i48pPRE6e7M3dXbeirhafyFUg9szaerEdK/HZ3X6Rmjlm5LwXCkYWGv4+cJYH9iPQJHxVQxVsVfixQFetrV8VesakCnf1UDqr6Z/fVBbkR0OdyTJzhAHtow+LYsM1BfSNZAXj1wL8xAwD9WHuC9SNY5wHj4j3Gw9gI+uMVJAre4xX9kfnAn+ETZ3zwPEAMMDHBGRTsF3/WyzvpPuM92oDswXiwwyWpMJZ+4H6iWLeddEB8STLJ4nND2YNjVNFniMTICyIFbf5bg/8yXXI418pg0v2PziwLJi0k08J96KSlICAICAKCgCAgCAgCgkAWQYBrzGaR6cg0BAFBQBBIfwSgdzBn1db9IAQgTF2/acu2JBVxOLJW3fsotuyFwCGCkHgqG5kQEVS+KS4+Lg7B+3FffPLBWRci1Ivm/jjt4d59XwBBAbtVa9ap1+nhXk9Cf2HgK88+zjPnp70rhVWtNnTM5B87N61TRRcpZkHuBTOnTTaixWV3Vv+yeIHxXv6CBQvj2lFDtkBqEEfw+LmenVq//9lX34K0gNj4wtnTp0CrA9oKeMocmhkRNWrXfbDH40+jtBaEwN97qW8vs3Fnfz/pa8oQaTF0zHc/Tp80blRlEtnu/ezLb27d8Nuvn773+gtmfUqVrRCCYO361SuWmt3n7AYINev3QYoUouj63B8mf+NKTB19jf1gY9nCuTNf++DTka9/MHTkV58Neg/leNp07Naj9r0Nmx7Ys3P7JVowHgv+4T3mY+Yf9htIC7Nxjh89fAhloIaO/W4mSn3NnzF14qqlC+fBDnEKCQ8tXCbnjXZTMybWFPu9YYs27UhD5XjT1u0eRDmiJ7u0bayPgwwiiIT3fLLfy3+TKDiyeuo3a3V/q/adHwZBN4dw5fYgULDPt1FJL3f226bfVi3HXur17EtvgMzB3B9qeW+13v1eGXD4wN7dPYngA4kxmXQ88Pn033/9Cbszf9m4G+2x9557pFNr+MTjsZbEi299NPQwZdvoZF9K9xCJba8EIfLKwCHDf6E90aPPc/1BxFG2zG7oYkBPY9LcX9Yh2O9q/7qDB9oQb4YSO+qRJ59/Gd8H4FyfSry1rB1aAoSaJ+uREr/d3Rfuzic7taMAOILn0IPgQHuijoRvsRsqfzt/la+LXV076FB+5SzKHnRVeRXggDoC8lzuiP/Pz4F6Fq3GfQTxkS0AYoAPLqOEzwjoM5nBRAYH+fk62jFpwcLYrBOhB99hF31ZfBufURaOS1PBDyYq0B/tkA2BTDHOLGE9DbOgPvzRM0Tgl06+6KLd/B7zRh8mB5gYAfF9Vdl8LCogxKq881hV7EWLyhFmUedWwE+0B8mCdnjPZae8aM1iLU0SMjFSc+gZH5J1kRokpa8gIAgIAoKAICAICAKCgCAgCAgCgoAgkJ0RQDkd6CWMmjJn8apdx89FnbjoMJ5bjv4bO/fXqAN4arp1x6493NFwQNbG/DXbD7Et2Pj862lzqCx/QnknPhCwR5vNR87F9H9n0DDjWoyZNm/Z4k37TupZCNwGZXA2HTkbbVZWCeVcYLfDQ4/2uRPrW7Neg8ZffPPDPIxvhtnsFZv3durR+yng62p83Ptw+LjJNzE6dj4OT/YnVUpryoJVmxC4dWVzwqwla5Zs3n9bdkUwqTAv2rDnOMSMzfqiNNcWGn/QyK9Nsy96PPHcS/o8YavnU8+/gkwS3R6yIr6ZtXg1smLMxql1b8MmrtYFT+yv3HnsLO4PGzdllo5DsZKly+I6SC2j3dSMCVuNWz3QccPh09dhf+mWA38asyV4PJB4a/f/fZlxWEMZD68RiYNsHt2ne6kUGfaznnmS1B7EmuD7Bbsrdxw9wyTd9z+vicL3Btdgk22A9Jm5fONujP/pV5NmGMfnds+++s5H2J/G/ZLSPQS7ffq9+tbW4xfi4Sv2Lko/Qfgen+Hr4FETvkeWSmq/c8jSmb503Q7GGvNAJotu1931SKnf7u6L1M41K/WnwDeC3yXpLEdnKTpLJ7z/rUyoY98LoY6/p+IMd5xZEOqIORtC/FcFOsPoxPsI5/tweq1KZ6TzGt5X0trgPj5XdrbHaxVne/TByf35M8ZAn1Dnifuwo7fF+Di5D96jDWyXcvpakl7L0lnGea2i8zpeyztt45VPjIsT47FPeNXH4XsYh8dkH/T5MC54xYl5Yz7og7nBDsbFPeBZ1hFzMdRxeVcVx9YmlZzrUYFe8R7rg7XBGuE91kwngDzeljQeC3BDhJvPm0Lczvsiyu0xstJBEBAEBAFBQBAQBAQBQSCjIyBpxhl9hcQ/QUAQyNQIoMQPgs1DB77+4l6qRw8BZJIvuASRXWOZIHcmiiA4gq+UqOG9f8/ObefOnD5l1g+6GSg7dJoGMt6v16hZKzwdrmtkcBsQJwjeGoWp+T4yHfCkOSWEGMtuuOO+W21ApFQIrRKBJ8xJgsEPJWz+oJJaZv66MogyPwhuQwz7r5Mnjrk1sItGyIYhN/zc0U4wmoAPV5HCoGVM6G2KlihVpnS5CiEoVXRg764dKcEVJE0Jyjz549jR31HqyegDMlRAriCTwHgPZM6eHVGbf/zumzGeYJTcmLAF/QyUnfr37OlTRmF3fSzgGxoeWQPlq/bu2rbVTDQdBATKLpll/rjyG98ViGFjr2MBQMIg+I+sjpef6N7RVYm25HAAceRpSbTk9hCIJazTQdoDyCQBaVL9nvsafjygf19P1yYp/5GJUy6kUhheSRR9L/RojO3dWQ/ukxK/3d0Xya1DdrlPQW9kVoDERPAbp13loWSlwMo+KqhxnLpKVf2CGlKxI9945VsylrIBODOCCU49u4Bh44wJZDUgIwGfUYqJS8Wy+DS310WycQ1tkRWBE9kPLNiNewm6MHTowtj8nu1zhgXssP6DnuWAdriOdhgbmRW4xuWi+PcL+nCWhNmWYE0NvQSusT23wXXOPoFdLmfF7XHvioq7FqcubrCruMtWdXa+TZ0ciywsZFjgb6+OZQJGlGWRkNmU2gOEhQmuN80mweOndmjpLwgIAoKAICAICAKCgCAgCNx1BISwuOuQy4CCgCCQnRCoQUFHBIU7N6tDIrr/6QlkJwxkroJAeiIA4uKFAR988lDvp5+HH6/1fbTLkvmzUqUHcafmUzmiWs0hoyf+AILmCBEKHRrVqHSnxkpLu5nV77TE4E7YIrIiP9ll3YrEgHrBLlZV4GEKmF/1Ud75Y5TVz0vZ/C4rv4r0SqWLUMIoMcDPmVrox4H9xFJSiYF5JhZ0HQcmDThgj2lxKSI9cM+BfQTpMRb3Yx0JLg2F/q708lizgrUsWIxb7wv7XHKJfWF/mcRgYkFfAt3XpPT6MDYTOmwXnxkfYykpjBGn4q7HqugTsepilJ/6a8JFdfZnkDYg/4ADl6viclaXiLQwfbDAkz2DbArNV+5qLBPlsmyUEBqeoC1tBQFBQBAQBAQBQUAQEATSGwER3U7vFZDxBQFBIEsjAC2GtvXCywpZkaWXWSaXQRFAGTNkOEGvYdo3X42Am5RR4pZw992eUrdeT/WDr1Eb161BdhQlUGVIP424ZFa/7/b6ejoekRUoAwbheiYbolW+B4iseIhEoItblU++WBKBptfCDhVQ2UFkBYLsyEhAoBzBfF1HAsOzILYezOf26ItsCdZxQBs+0df4gBNIBA72MwnCbXAd96E5gSyDpA74iewEFgNnsoBfWZwbvoG8YMFttGfbeiaHcazkfuew74wPslJwjckT47wTyRGbr035lrEpn0KxKl9nX+VfHvNlsgA+wlcmigKda5kMTIdkgwAAIABJREFUFEnf1oS4GQPRtEgVotJZEBAEBAFBQBAQBAQBQSAjI5Dcf+Qzsu/imyAgCAgCgoAgIAgIAqYIQKNi2qI1W6mCk9dDre+rfvnShQsozaWLZWcE6AICA3OgBNTL73z82YiP3339/VeefbxI8RKl9uzYujkj+OfKh8zqd0bGlH2jADee2EcgH0F/nHaVo2pOlbuuj7r+p0VdP2FVXgUtRCOQ8HbxK8piA/EAgWdkVyCQrYtOc0CfSz5xFgSXjsIriAPO5EDQXicO9FJEGIeD8RgHnznoj/cI3PM4l533XUEOuyz8rZMjuMZkBPziNkyE4JWzMmAbbY1lr9zJINfH5BJVTAKY9devWZXFalG57yWyqLyFMl7gI4TOuZQWiCbgyOvn71zTVG0/kBbO00GvZiffv+01VQNLZ0FAEBAEBAFBQBAQBAQBQeAuI2Aq4HmXfZDhBAFBQBAQBAQBQUAQSDMEnnjh9Xee6v/GewtnT5/ywWv9nrhx/dq1CqHhVfdmsOyK4qXKlBtOQvPQr3jqoQeaIiMrJCyiGjQmoC2SZoCksaHM6ncaw3AnzYGw4Kf8fZQ9V5zKdY9d+ZW3Ku8ClHORx6LsOeKVNRcC7Tg4ewJ9OBMBBAQ/jc+ZA+yzHnzXNR3YDpc1Qns9IwP2ke2AAzYCnPdZa4KzPJgMcOfBKC5NxWNxX/YdRAAIGMyBtTS4DRMmKVkLxkAnKYxaHWZ2maBJJFICaliVbzG6Fh2rjnwE8gTXmTRCJgiXmsKagsCQQxAQBAQBQUAQEAQEAUFAEBAEkkHAnR8SAqIgIAgIAoKAICAICAKZAoFX3hvyxdMvvTlw3PAhH7z1fJ8eICsgEh5erWadjEQClCpbIeSbmT//avf29u5xf6PaICsAcHj1WvdAfH3fru1RGRHwzOp3RsTSzCd6Eh8kAILbCNQnEg2577Mq/4qUB1GASj/5WlX037HK4h2t7P6s98BB8jPU/l86ERhHQB79kaWQ1MGBe868YKKE++j3MR6C8CwCjiwKBOSRWcFaEvAbR25nO3eh56wOJhBgl4XGMR7mwr5hTjw3nfBwdyy9HZe2AtmAsUH46IQOZ6vofRhbL+VFrtjzWVTBXt4qIISzKpik4CwWYOLnXNuU+Ch9BAFBQBAQBAQBQUAQEAQEgWyFgBAW2Wq5ZbKCgCAgCAgCgkDWRaBT915PQlz729FffDJ62KB3eaYIsucKyhO8fcvGdRlh9n7+/gHDJ/wwD3Vbnuratolepiqy5j33Hti7awfxLCjvk6GOzOp3hgIxCWcooI3/lwfRyaWQEKiPV4X7eKnctW0q9hLRF5Q44VcqXtlywRKLX6McFE5kP6BPYacNd0sjmXll1IbQiQv+/cDkAvzV20N/A0SCJ78zmHzh7A6jDgfuwyaTM1wGytMxjHPVtT84c4O1M1h820wvgvU+bMpKvIp3UauqNNGHNEXYb/RBf9bnwPUg5xpnli0pfgoCgoAgIAgIAoKAICAICALpgoAn/8lPFwdlUEFAEBAEBAFBQBAQBJJDAJoKLwz48FNkUYwcMvBNvX3dBk1a4PP2LRvWJmfnbtzv+dTzrxQrWbrsB6/2e+KPE8eO8JhWm81W696GTTKKn0YsMqvfd2NN02gMzkpAZkGiCHahJ+xU/ok0EyjuHViJKAAvh/IqbFFWOwgKZFLg//JcpqksvS9CJ5MH7riVFKlhpg2B8RCsx/j8ngkWZIdwwN6TzAcQBKyNoZd9Yr0KzIP95IwHXYvDnXnqNvT2IBaQKYKTxcSBJ+tauBIORzZFYrksq51IC1u88i9nVSHjdM0PjAN/YQ9rCvICayyHICAICAKCgCAgCAgCgoAgIAgkgYAQFrI9BAFBQBAQBAQBQSDTI9CgeZt2IC0mjRk5DCWV9Ak1aNGm3d6d27eeP3cWJXPS/WjdsVuPo4cO7Fu1dOE83ZnqtevVz5krd9C6Vb8sTncnTRzIrH5nRCyNPtGT9wh0Q6wZQXMEy/2UX0m7yn+/l4qn7WyjzAorxbu9i8RRcBxtIMqNYPo/zvcgKlB6CIQBB/PTeupctomzJ7g0EsYx6mK4+xsD31UmJsyyLHgsznJgu0ymuJNFkhQOwAsluFh3ApgCf7xSSstNAXPYMGZa/EfoWG1EKgXEqBxVvFXe1nr2B/yHfRYlD3SudVqvjdgTBAQBQUAQEAQEAUFAEBAEsgwC7v6YyDITlokIAoKAICAICAKCQNZDoETpsuUxq4NUTkmfXcky5SpUrVGn3orFP83JCLOGoHaRYiVKHdy3e6fRn/bdej5+7erVK+tXr1yWEXzVfcisfmc0HJPwpyjdw1P4ICISxZrztrMpW4BDWei/61cPUADd+1rCk/yJB2cBoDaULtLtTgBfD7zze7OyR2bucqkjjMnZFKwvgfYYP7nsCn0sBPIxF8yLdSSMmR2wq5Mk6I+2IDu4D9p4Ohf0Ya0M4M7jctkpEECcrcIloBh/nisLn5OHXpRtkV+pPI0YNxYjR1+sKcbAGmOt5RAEBAFBQBAQBAQBQUAQEAQEARcICGEhW0MQEAQEAUFAEBAEMj0C165cQUkXlTN3bmgA3Dz6vTFwMDIu5k3/bkJGmGRcXGxs9I3r15FJofsTEhYe2axN+84LZn3/HYTCM4Kvug+Z1e+MhqOZP/TEPQL/CIRzeaJoFdQkXuWIpFJD3nHKcSNe2XPFEnmBdtgbrOcQTO9BHCAzIzmSgIdOLGP0X3DfWMLIFWTwj8s2IQAPkgJjIwDP2QlsWw/qJ0WEIKAPv1nnAb9L8NnYnz9zuSi9Hd5z+SYeyx3SRp8nZ0EwoQA7yGJhkoJ1NfBZ/+3Egt2Mp43IJYcKbmtXQffBBtYKtrnkFf5GJRA+zjXPDNtTfBQEBAFBQBAQBAQBQUAQEATuOgJCWNx1yGVAQUAQEAQEAUFAEEhrBNYsX7LQQcdDvZ5+HmRA/oKFiwz4+IuvGlKpqDk/TP7mn7/+OJnWY6bEHnyEr5G1694XWavufb5+fv731G/cfPiE6fNjYqKjJ341/NOU2L3TfTKr33calzSyn8cZ2AYh4Z2gieBb3Fc5Yii4bbEpv9JWFRhJoXIbMhHwf3cuY8RkhScBencJCuPUOPsAQXtkHrBANfzBexAYZqWouIwUEzKwy0LXIBr+y1BItGHMkkB/JiV4LLaBz7pdvu7JsmBMHDrZAVyRuQIihf3jzBFj+SqeX+KrzW5XviWtqmB3O5FNwMkovM16H1hzOQQBQUAQEAQEAUFAEBAEBAFBwAQBT37gCICCgCAgCAgCgoAgIAhkWAT69Hv1rb6vvPWB7uD+3Tu29e7Usv6Vy5cuZhTHCxQqUvTrmT//itJQ7FM8HQNffqb3vBlTvs0ofhr9yKx+Z1Q84Rc9aY+gdj6njxCtjld+ZS2q7Md+yrsABcD9rMqe5xqRFpyNgIA3DgTrOdjuaorJZRxwRoSxv9l1BN6RIQAf+WDCQP89wdd0MoHt8TX0hy3WwEAGAsgBfW66T8asENxjooBJD+7LmSZmWSTJ4aSTEWjL2SM8Hr8yWYNXFh5nMiXx3qUd19ShV73UucXISsHcMEcmXyBYjuO0pUlCJoccgoAgIAgIAoKAICAICAKCgCCgISCEhWwHQUAQEAQEAUFAEMgyCCBrofn9HboE5siVa2fUpg2zpk4chxJMGW2CgTly5oJmRUhYROSFf8+dnTfju28hDJ7R/DT6k1n9zqi4EmGRl3xDKSI81Z8Y0C/9vpfKWZ3KC9njlcUnVuWsFadsPgie4+CSSRxM17OlXREQ6KcH/T35/z9rViCzAuQAZ1LADzNSgNtzIJ91HNAW5AzbQTvMAWWTEMzHe5AhPB+0Y7+ZDOAsDx4D9znDgskQ2EE79Gcfk1p+HTM9a8TYR2/HvvF6cD8uGXVDxUXHq9MzlNrdnTUyuHwU+4l5XyXC4kxSzsk9QUAQEAQEAUFAEBAEBAFBIDsi4MkPluyIj8xZEBAEBAFBQBAQBAQBQUAQSHMEiKzIQUahZYKAN4L1DuVbzKrKDvNRXjlIuyIuTuWsHa28grmMEPvAmRXJZRHomhJmQtbuzAlkH5dqQtCdCQH05QwD3Q7aIJspJ50gIlgUG4QMa1/oZaDgF2chsDYFEwCsWcGZDyAgcOoC2Ewe6CQCExwsms3+JUXo6HoUxvkYS+gyYaLrhujjo/9Vdf3362pDONE8l7F+yLJgcgVzRpYFXv8l0uKSOwshbQQBQUAQEAQEAUFAEBAEBIHsgoBoWGSXlZZ5CgKCgCAgCAgCgoAgIAhkJARykzP4vzgyLBJLPgVUtJB2BYls56HSUOUsypabywjx0/scJGchaldEBOyh7BJemTRgIsATDFjHATY4OwL99WwHtseEAETAmZTANfRDfxAfLCjPQtYsbs3khG4L79EffXUygzFgPQ+eJ9riHmwatS3YZ7apv+K9ro+h4+PqtxL7wGW3+DN0RhKJHe8SVpWjBuau+4N2wAZrDtvYA3IIAoKAICAICAKCgCAgCAgCgoCGgBAWsh0EAUFAEBAEBAFBQBAQBASBu4gAZVcgYM1lkTgYb1UBVWzK7m9RVl87aVg4SGibS0DhKX0O8rMANDzmgDnec5AeGQ7nndPBeyYSPMmsZnKDxwLZcFUbA+Z1soRJCc6GYM0L9IHvTEigD7I0mCDAK2dt6BoSPD4IDtar0DMkGAv0QSYFcAJZgPE4A4XHwHX9gD0mYPTrnv4u4qwMtgEfkEmSSF5Ybb6q4CPABaQPY/XfWjs1Mpx7weCifBQEBAFBQBAQBAQBQUAQEASyLwKe/sc8+yIlMxcEBAFBQBAQBAQBQUAQEATSBoFcZIZLLXGJoRjKrohR9nwWZQ+KV9ZAFqXmgL5OODBRYRS8ZnFn9DlHp15+CZ67Ii104oNnyCWnmBxACSsOvnMb7sdt+DOXSOLr6IdDL9PEQXy9VBL7x+Wf0B5z4YwSI/poxzZBAgFTXega7Vn/Q++LfmZzdrW6xjJWaGf2O4ptJpbxKtAR82Gih0tk8XzRFv5iL8ghCAgCgoAgIAgIAoKAICAICAJOBISwkK0gCAgCgoAgIAgIAoKAICAI3CUE6Il6/P8bgWw8jY8gNjIAHMqn6HWVt52PijnjUNGnYugJfT0rgb0zIypwD3YQqEf5IWRV4JUJC1faDWzL7D6TFVySijMhMJauncFkC9vgMk2suwFtDrZhNgcW3NazKIwrwdoZZgQDj8sZGbCHklQ4mGRw9XvHSGQkRWBwposr4oR91rNg7MqWg8kWxgAZIxgHaw5fsQcszj1xl3agDCMICAKCgCAgCAgCgoAgIAhkbASEsMjY6yPeCQKCgCAgCAgCgoAgIAhkLQSQqcAlof7LTMhVg8iKP+NUYFi8ylmN9RgQKNdLL+lkAaPCwXqQFGiPp/YRrEcwHNkHrvQZOJvBVdaFfp/95DHN+uq6Dlz6yNiOiQkE/nURbp6vbp/9NhIe+m7ge8jgADkAbDF3nOjPZaaMO0j/DWQkKnQiB/1gg8kPd8tqsV+BqrGDhch14kXPSMFegN9yCAKCgCAgCAgCgoAgIAgIAoKA8z/yAoQgIAgIAoKAIJDlELDZ7fbAHDml1EaWW1mZUEoRCKAvRLmQylVKla0Qgu9HSu1k9H6Yp7e3D5cgyoju4u8Sgtd4wh7Bal8VVM+iglv5qMBqVmUL5KwDPWCvz4OD5nr5JZAVCKrjGvrhcwHnZ/TlEk26HU9KIhlxhD0mHfDeaAu+IMuCMyB0kXC2hSwDZIUwucHXMT+2z4QNf2ZyxugPZ6PAFvY2n0aixawf48PzMcuiYPLDjDAy2tQJD/jhpUIn8XrDDuYCIglrj7XGPfm3yoiifBYEBAFBQBAQBAQBQUAQyLYISIZFtl16mbggIAhkZAQQTPz+5zVRjVs90DEj+2nmW9dHn3h2wKDPR6e3390ff+bFX6IO/Z0nb7786e2LjC8IpCcCIO4+HD5u8sqdR89MX7J2+6wVm/as2nns7DOvvv2h3e5lVt8/Pd1N9diD/zdh2mfjp85OtaE0NEAlfxIOeuVgPGszRCtfKgVV+Bkv5VOcaIaT15V3fgS0OasiKVKBg+cIeqMdkzQI8iMYzsF7kBdMKnhCUuht9dJPsMVlrZgQ4N8U7DeXhMK0OasC5ASIDPTHifcI6LOguF7uiu1zf56Lnm2irxDmrJdjMmZ4ACPjoRMLTOgwWQHfdAFxYAj/dRxdYWksp+WvCvbwU5V/YPFx2IWuBezh+4e9EOfcG7xHTNyVS4KAICAICAKCgCAgCAgCgkD2QEAIi+yxzjJLQUAQyGQIlCpTvmKF0CoRQcF582Uy11WvZ196g2Kg6R4EDatavRaCsVevXL6c2TAUfwWBtELAQsewsd/NbNCs9QOff/jWK52b1qnyyAON68ya+u24Xn37vz541ITv02qsjGKnSrWadfwCAljHIKO4xVkRuZ1B6iv0ioB3nMrbNkA5ou3KntOicoQZSxVxmSXMw1XpIiZB0AbBcATGoR2hkww6ocCYcGA9qcC73lYnJ9AHQf0LzjH1duwH6z5weST4hfe4jsA/Slbh3wrOomCSgrMyuLSTrlNhhgOusU20BQliLN1k9m8Szx+YQVsCGR84mNxgYgWvnC3CPulZIGb46cQK/IlRfqViVLEXYQfEEgglJj+wF+Bfbo3YAnEhhyAgCAgCgoAgIAgIAoKAIJAtEciy5QCy5WrKpAUBQSDLIBBRs049TObIwf17M9Ok8hUoVBjn9s0b1qa33yh9c/jA3t3Xr13Dk6xyCALZEoFGLdq2r1mvQePX+j7aZcn8WdMZhJ1bN60/cujAvnc+GTmuVfvODy+cPX1KVgCoUNFiJXLmyh10YM+u7RllPhR4Tnj63xmARrCaA+rxyiuvtwqsTFdyW0igOV7Z8uDvFcgWDrhzqSNMRy8Fpd/nEkMIuIOowJP7OBB4x2cjEaBD464mA/dh8oCD+ZiLTqpwO7aL+XLwHnNhkgABeviJ+1zmydiOP3PGCQf4dV0P3X8zP5LaBkzosF8gt4Po5NJQICfgp078wB7GwT0mLdgf41jsG/D3UoGRFpXzUJwKbu2lzi5gPQsmmDhDhomVeEsT0zJeSc1H7gkCgoAgIAgIAoKAICAICAJZAgHJsMgSyyiTEAQEgayGQHhkzToOOvbv3rEtM82tUpWq1eHvDgqGpqfffv7+AUVLlCqzZ+e2Lenph4wtCKQ3Aq06dOn+x4ljR5b+NHuG0ZfZ0yaOj9q0bk33Ps/1T28/02r88iFh4bC1Z8fWzWllMw3sJAasE4kDZBUgSJ0YqPcuZCPSIp7KQjko/E2khRfICjyFj4MD4UZNBZ244PJMsI2n9rk0EogE6CJgXIzF1830GTCWu6WiOJjPZajQ15XmA/zkeesC2PpYTN7ov0l07Y6LZEMnnXEPxIKreXiyXCzMretegERhHRD4hnESdSgSyR8maJhMSe63FN/3VVbbdRV7XqmSr1qVVx6MgzVhogLjYG/wXvGUSPJk3tJWEBAEBAFBQBAQBAQBQUAQyNAIJPef7AztvDgnCAgCgkBWRaAylTM6cfT3Q5cvXUS5jUxzhEZE1rhCTh89fGBfejpdvlJYuJWO3du2bkpPP2RsQSC9EQgNj6xxaN/unSBAzXwBkVE+JLSKj68fgqWZ/ihXMTQMk8hg331oFOSgMy+dCHrjTHx6P6ACFSM6alXXjxNh4Y014if6WUCbswt4bfRAvZ7twOWacB+ZFrCjZ2egP2cS6OtsJoad1D7gbA3WfKAIfMJcjH4Zx2BfEYjnDJCkSAe0+5dOzkjBnPRSUUwspGbPAiPO+MC8UBYKRAwTJky2YAz+zWTES18DM194TaGBEaCsvnHq2iEHCawzcYUxgB/vC+wR7JUs8X1MzeJIX0FAEBAEBAFBQBAQBASB7IuAEBbZd+1l5oKAIJBBEQgghdwSpcuW37098wXbQ6tEVt+7c9vWeDrSE96QyuGRGD+DPWWdnpDI2NkUgaA8wXnj6HA1fWRZdGt1X7UbVDstK0BUITQs4uqVK5fTmzQ1YMklWFm3AFgnZjz4l6M8iBoW5VfGonxLc/YCuqMPZwDoZBMLWCfqXyS24/foh4A7Z1pwpoauAWF8cp/t6WLSyREJ7BeLUOOVA//wwTgG/97gjBGQEPATrxhLnx9s4x5s8tz0LA34ibJN6JvU7xjGBPZcHZxJwdknwU7fOYuC8WWhcF4XnUTitWWSQx8L/fSMjVhVoOt1ZfGJp3V3kGYJE0oYH3sCdrF2PE4SrsstQUAQEAQEAUFAEBAEBAFBIOsiIIRF1l1bmZkgIAhkUgRCwiIiIZS7a9vmjZltCniae8+OqHQvxVKRMIyJiY4+uHf3jsyGofgrCKQlAhcvnP83X/6ChVzZhMbLwb27ssz3BNlVe3dGbUlv0pTxJt0KJh5AHnDg/b+n8v1KW1X0+Thlz4Vretkm1kgwZsaw3gOXKtLJCAS8OZDP5AcLXptl2LAt/B5g/QddLNps23DGALJGOHME43KZJjNyzKhFAUIC/vEcdT0OXANml+iEXzwfJhF0giCprwqTEUm1YZKFRbb5M8gD+IfruMbED2yxXcYV11jLQh8L7dAf/iI7BG1syuLlrfwrOFQO0rPwL4/5MfnBdrFHMF6sU/skKf/lniAgCAgCgoAgIAgIAoKAIJAlERDCIksuq0xKEBAEMjMCnB2wa9uWTEVYFC1esnQuepx7z/b0JywqhUVUO7Rv767o6BsIFMkhCGRbBA7v37u7LJVJQom0rA4CstOKlSxdNoNlpyHwnZtO1ifAMiAgnRikv7jNoaxeFhV31UoaB1wGinUNdHFpXj4u/cSZEeiDoD7b5Cf9dYFrJi9YR4Kf/DdmHzBxkJR+ApMPTICgfBF0N0Be4DDuM6NeBe6jLQL5wIRJEyZeuEQSXtGG54tXznTg+ZiWOXP6wX5ylobZ9uf+wI4JpZz0HnNCP2Q7cBvOBOGSWEZ7TKTo17m8F+NuU1Y7rXOAt3IQl5GrFvfRSRG0BS7YM3IIAoKAICAICAKCgCAgCAgC2RKBLP/jNVuuqkxaEBAEMjUCFSqHV42NjYnZt2tHVGaaCHQ34O8eero5Pf329vH1LV2uYqXd27eIfkV6LoSMnSEQ2Lj21+UQoY+oXrtuhnDoDjpRqUrVashOy0iEhaXJTdFm1kZAkDoxUO0VZFNB9Swq9lIslQfCFQ5s60/+6wLbaIMn8vnkYD6IWZQeQlCdyzlxtoau0cDocz9u48mqMMEAuyxGzUF8HksvKeWK/OCyUDrBwoQNrkHTASQC+8r4cKYFkzm4bkZc6OMmR8Dw7yH2hbMe9BJdGMe4FjpuxjJa3BeZJ+xrop9WKgmlbPEqZ12yZ+XMFt4X8CEhM4P2jstSbp4smLQVBAQBQUAQEAQEAUFAEBAEMhsCQlhkthUTfwUBQSDLI1CxcpWqKGUUfeM6RDozzREaXq0GRMJPHjty2FOnkZnRuOX9HfwDAvCkbqoO4Gez2+0ZKWiZkgmlJSYpGf9O96HgcvXgvPkLpOU41WrXqw+7aWkzs9v6demi+ZhDI/p+Zfa5JOc/r/2uqAxXTg9/yxGgR3CaSzlZVHALu7Llsqjov0lwOzcLUaMNZz4giK1rQwACPeuC9RG49NCtgfHEsbiNHvzmckap+R2gZ3pgXJxcBikpggBtuNwSZ4Vwe9jQ56zrQuglmIyB/KTGS2rbGLFlfDnzIVEYPZE0YRFztDEbT8+84PVDO6w7EypYpzjllfuq8i1iV1556X48rxnGBC74jD6Z6t//5L6bcl8QEAQEAUFAEBAEBAFBQBDwBIHU/FDxZBxpKwgIAoKAIOAGAjly5spdqmyFEAq2p7sOhBvu3tIkNCKyxv7dO7Y56PCkL8iFKQtWbRo69ruZbTs93NOTvmZtUQ4K13ensKRWybLlK3p7+yBglG5HWmOSbhNxMTCe+J84d9na+b/tONz1sSefSwv/2nV9pPf4GQtX/m/yrEWu7JULqVwlLcbKTDYO7d+zC2ejFm3be+p3RvgueOJzGGV5nTtz+tSfJ48f9aTfXWjLT9GzyHJi8D1HDauK/TdeBTf3VjZvBMQ5OM6BfNZ5YI0FuMpP8nMJJQTHWWMBdvEZbZB1gcA+kyToa6a/oE/fnb/dXGoJ/Thwr2cXYFz4wH4Y4WWtjv/KYiW20LM98PtEzxDRiQX0Z1IjLZYuqawJrId+8DomNa6OsY7Pf1kxFu+r6safsQnoFX9Znydn2DAeaTG/NLGBf9adp8XwHp/5RBu8t2rXEu6liRNiRBAQBAQBQUAQEAQEAUEg2yAghEW2WWqZqCAgCGQGBKpUq1kHteYzgnC1J3ghwB5SOSJy787tWz3ph7Z2u5cX8TRBIDqO/n5wv6f9je2R6QEh4cMH9+3x1BZ0OGYsXbcjokb6ls9Ja0w8xeFOt7929eqVF3t3a3f50oULr73/6Yi+r7z1QWrHzJM3X37YOHL4wD4zW607dOn+/c9rooBtasfKbP0Xzp4+pVDRYiWq17m3gbu+Z5Tvgrv+ol1YZI3aO6M2b/Ckz11qC8JBD3ZTUNsSr3yKkFpCuE3ZcziUjbQNEg8EthH01p/S1wPZeoCdszH4lbMp8Bl2sNf5CX7WYOApG8kJLvWkQ6LrSyQFFWc/YAzoL+DQy0Pptnku+vh6QNsVacJEiY6Fq7ngunG+yS21WVBdv+aqPJOZv7yW8AGZElfoxLXEsl32wBwqsIpVeRWwKKsfZ5zodrBmOkmVnO+pvp8ECQHCgfeQXkqM9UUYI319OOOG74HA0EkMJj9uvqZ6AmJAEBAEBAFBQBAQBAQBQSBLISCERZZaTpmMICAIZHYEqtaoUw9z2Ldre6bSryhboVJlXz8//327tnlMWNwgdqF9/WoVW9aqVHzD6hXLUruGoeGRNfYYaJIDAAAgAElEQVSSH/FxcR7X/252f8cuNmJf9u/ZuT21fqSmf1pjkhpf7lTfNcuXLOzYqGbotk3rf+v97MtvhlevdU9qxprwv88Gd2pcq/KTXdo2NrPTumO3HocP7N0NfZjUjJMZ+8774bsJmHfnRx7v667/GeW74K6/+QsWLoKTykG5RVjoT4BjDOdns6fIE66l8mAB7P9ICa9cVnV6roOetI9X1pzXyD7/veLSShgSAV9dk4Kv4TrICATAORDOWQkgOq7SyVkXnGWBPjppYgzQ65kTPF2+ltwT8noGBDQbEKTHqZMrTCCwloer3yB6ANwIO2Nh5rvZEiXnt6tlZbLISCK4M4YxGwQEDgt/w/9E7Q57cLRyOJNgfEoAC15/Li1l1MRI5Ra8tTtnPfD3wLlWTDzBB13wHPtGJ7+wtzjLRW/LwuUYTO/Dpb70El9pOh8xJggIAoKAICAICAKCgCCQtRAQwiJrrafMRhAQBDI5AlVr1qmHQPvh/Xt3ZaapgCSAvykVCj975tQ///z1x8nUzjkgMDBHiTLlKuxKYTmo2vc2bHrk0P69F/49dza1vqS2f1phklo/7mR/kjw5/8azvbohmP5w774vpGYsZOiAkIiJiWYtgJvmkFVRrXbd+lEb165OzRiZtS/20i+L5s1q2KJNu7z5CxZyZx4Z6bvgjr/ITkO73Tu2btSDsbhmVqaGtLm5pJJNK1mj6xDo/0fWy97cLInDfrlBaARR21ttB4Q4VHBLi/IKtipboC/d59JNetkoDpjrgXcO/DMRwSWWsO8v0gmygsfi8kn4zASGKzgZD76vB8x1MW9X/eEjgtj+Tj/QDr7AL0TmmfzgDCdPWCBuy2uSUiIiYTu4sZ9YwyIl4zCOvAacMYNXXEvUG7H50xhkPri5RQXVhkv63PAee+aOHM79rmdOMKHAr1gj7BfsS2ABkgXEC175hN4UTlzndvicS2uLe1z6SxcVZ/LMXULsjuAgRgUBQUAQEAQEAUFAEBAEMi4CQlhk3LURzwQBQSCbIeDl5e2NwP/xo78fio6+gQBPmh658wTnRVCvYJGixdPUMBmD3yjD5KocT1LjQbMjKDhvPnd8oiCjJSl9CZSDQkmt3VFbNrpjz9gGmSIpJTs8HS+p0kSeYOLpuHr7jFAe6e8/T55Y8fP82fc1adEG6+tqPriH0mNm9/HdQTkgV32LlypTDvvG07VNDp+AwBw5U4J/UnNJiT13+syY9PVozKd9t56Pu9Pe3e8C1sSH0qvcsWlskxy+enuMY7XZXGoI4G8bSKtz//wJ/R+um59QTx+f6cTeuSlw7LyuPx1uP3nypM/AgQMRkNWfNOcyOGyH73mSecEBfzy5n/h/b79Qi4q7YFHx0VQWyMbkAI+F4DZrQDABp5MXTFrwfPDvBfpiPyJ4DNKAn5DHaO4E6dGORbo5OwL9ML67gXu0Z7FoLoOEuaA/fGRdDbMMBldbiIPaZiWrXPUxK3fFOOhzcRcXd7e3MauPMycwX8wdwfvEeVisN9T1I3T1H4uy5WH7aM/rniYZFpruBGtLsGYGxgIxwd8L7HvsHc6kwCu+19yGiQm0wQlyAvsNey3A+QqbTGxgTrCNtpgz7mEMts9loxL2qSHDyV28pZ0gIAgIAoKAICAICAKCQBZFQAiLLLqwMi1BQBDI2AiAPOj78oD3v57586/TSTMBNfwhWo3A36F9u3e64z2Cfd16PdVvzPfzf/nwi7GTkgqePvZM/9eXbTn418Q5y9YuWr/nGASuUcLJnXHcaVOpStXqB6iMkqdlmBC4nTx/+fq3h4wYm9Q4wOu9YaO+Wbv/78vrD5269tGI8d+ZBbc502Nn1KabZWEgtPzqwE+Gv/bB0JFlyoeE6uPA7iejJ04fOfHHBZ9/PW0OiBPYGDpm8o+ffjVpxqCRX09p0Kz1A+5g4G4biB9jzTcdORs9c/nG3UYCKTlMChQqUvSDz8dMRBCex0Qw97G+L76GudzToEmLpHxB0Bf7Ycnm/X9sOHz6+mfjp85GwN9d/83a1bjnvoYvvzv4c1c2WjzQqRvWzNX9bZs3rMXex3oY25C8SZ53Phk5bs3ePy+u3f/X5cefe2WAsU3XR594dtLcX9ZVCK0SwfcgwPzlpJkLh0+YPp/31/0PPvwor+3Az0ZPMO4H7pvcGqEd8F++/fdTdRs2bYnPwPWRJ/u9DD++mbV4df2mre5PyVxSsw5J9d2yfs2qo4cP7u9AhAVIPWPblH4XgO246QtWsD1gin34w+Lftr376Zfjzf4uuYMv2ytfKSx8zLR5yzYeOn19Ha0/1troO4KdEdVq3XP00IF9hUuUrjd9ydqoX3efODtoxPhJAwe+j79zCJRyYBZ7nYOzCU+L9+rVu+AHn40ed/yK/XTLHs+cf/blt96l6+inB2k5wMqkQkIg3U1BYS7z9F+5p7hzFKjOSUrG11lrAtNCYJdJDYzDwWUW39YzDfgpdcyBNSvQjoW7dYIlOcKByQDur4t46yRhUkF03ANJAV+C6eTANmeP4BW+8jzx6o5fvNxmJatcbXnWhdD7mo2X3Pi6fVfkRlJlo5gUQEA/Ub/iv8C9RfmWjlfx1xzKv4xeOkvfK67md9t1TYNCL29mJN44y4EJNNzHWuskBouD4xpnSGA8/t7ABq4zAYHreI/1xXvMFQwMyAy0y00nskVAcOA7xfuaReZ5v/L6eLImbuMjDQUBQUAQEAQEAUFAEBAEMhcCQlhkrvUSbwUBQSALIIAnwSHs3PWxp577+4+Tx69duXK5T79X33pr8PAxmN6endu2JDdNlHVBUBSB+Jp16zdq3bFrj9YdunY36xcSFh753GvvDqJqOTtGDf3oHehjNG55f4eHevd9Prlx3LmPJ9fLVqxUOSVC4Xgi+vQ/f/9VtESpMq7Ggljw1AW/bm7WpkPnn2ZOm7x+9Yqlrdp3frjOfY2aGfuERlSree7M6VN/njx+FPe69HzimWkLf93S9bEnn0Og8+sfF62CwDf3g7BwwSLFisfFxcbmCU4Ubaa3sYWLlSyF0lIly5SvGPB/9s4CXqqqa+OHS6hgdyPSXQIWdisGNioGBgYqmFgYiIEdKIIC+oqEiYQoAgIiSLd0S3dd4Ma3/3Pnwc1hZu4M8JHrvL/znplzdqz97H1G7nr2Ws8BW7eLPtZ47rj/0SffbvX198x5hzYtP2Tc9zVsjHN005EbJldcd3NdzprnX3w5lSA4nGP264cbv/T6hVdcc/37bTp2OeKoY46N1T8k1zuuf9bDiL//GvBbtx86n3vxFVdfdGXtG5OZ63hlIHVuufuBRwufXKxErDK1rqtT99Krr68TL0KC1FDUCzu30ST46uc+gy+56vqbu37X/suJY0ePuN8RfawJv5+FC+b/y3fmU/chL2iPFFGHH3nU0aSdghQB88jcnly8pINjCwHuZOaIPoqXKluetc98Qf598vWPvzZ8rmnzQ5z4d1lH4F1/W736vo3JjmVb5iG3ut+3b9sKgkwki19+a98FyEq1A0nTvke/YUTLFDrgwAOvuvG2uxzMpf1+ksWXOpBvjtAcfGKRYsW//uKT9/+dPWvGI8+88ob/DkMYFC9eYp9S7ncO4fVnmr3bctTQwQP+GTNyxGW1b7xlwtRZN7umcCorrY0crJGd3nfedfcx19z18B8XXFH7+l5dv+s0edyYMXc9/MRzjzZqxG+SUinhaJVjV3n6tfNcxEAi+JUm6L8ogfz4cTOzg7RCOIblzPZT5OBUlvPYT/9EP+pT6aBwEktTgHHyfGuiB0ROyE7SF0mTASJF6Y3CY1XEhPrGdhHi+ltDUSO0l6zwve/Ip89kxiRSxSdaYtXTPeGsaBKNTc/jXVUu7GAPf8cOaVewdhSxQoRNWpC52kVb5PPH6a+V3F7pWM+1hvwIBpF1PgkmfPyoJUVLkNYJgoH51HoXKXFA9H5OaqscMoLFzJzqmcgJESGKwFCqKb5rjYp4823cmnFbHUPAEDAEDAFDwBAwBAwBQ8AQMAQMAUPAENgaBEqVq1iZKIH23fsNVRokHM4ff/V9jxGzV2ZznnJazXMStc0O+y79R06mLFEDRx97/Anf9Og//PveQ8ZffOV1N4XrQmpQVk7s/QoWLPRGi7YdcSpuzRjCdYhIoP3La98YkzDJrQ+iDV5v0aZDrHI4gr/9ffDYPqOmLyJFDWW4N2jygrWtO3fvG65D1MB7X3Tswn1202PXax990Z7d43Xq3f8I36+/7e77Y/UFaTR81oqsrU3zk9s4cerTP9ER2uFOpIvbDb6FwHciTN77osNPtFO6fKWq9HnrPQ825Hv9Ro1fhLTgc7y0P0RB+M9Ze31Hz1jMGsnN/kTPa11f53bavahW7RvC5Qrss+++f01asIbnrN1Y7UAs8RyHs55DrkBWEFnBe8N9SALKsUPfbwcCjvsnFStRKlb77NDnncttjKnM0RMvvvHe39MWr0c3hTkZNmNZBqQNmPKO+WmSUhlLbjZuy3Peg6HTl26ENEvUTrLvwkGHHHrYsJnLMyHAIGKJGmrfvf+wYx37QfvhVG+p4Hty8VJlWDdfduk9yPFOOFADfhu11vkuwWCnT3Im93/sO2xizbPOPsbdL1DjtDMKc+/F5h994b4f7M5j3XmUO/dzZyF3Hti1a9dDvu7ad5hbY6vq3Vv/AnfvhAcbPHIe9ereXf929/2QaNkj3fUg2qWeOwu6E+2L/O7MJzviYZrdKyjuzvLurOjOypFzdO3K2dNfq5ydPq+Sq1/SnVw5K7izrDsrurO8O0+OPuc7zypHn3HVqXpV3D2dPPO/J/pMf/RVzqujNmlHNpWOfuaZ+qZdPpdxJ8+xt6g7S0THg93hsqpDO8nYqHLYkVsdxkA5ztywoAx2Fo+O/fgoDowFm/1x6nMse2Nhrfr0UcSdrEuuJ7mT+S6avbRPuezFvapkz/6syqZ1kbNGWCubIuiSeedde0r5xHqESGWNcu7vTtY/J2uXNc3nI9x5mDsPj36WXdjIiY1gw1wWjl5LuSunMGaMVd0JJmBIOdZR9Wjd49wVTE+InryDJ0Zt4F3ixD69U9i+6X1ynyNp1zjtMAQMAUPAEDAEDAFDwBDYuxCwCIu9a75ttIaAIbATEcBxC1GAPsUjd9545bIlixdFnW7ZXTp93ZbP7O4fO3JoXP0FnPXOOdrlOLeT/PmG993+xvOPN0ADAP2IIm4nc6VTapweHuKxJxQuQruLFsyL7EJft3btmqceuOPGfr1+6bo94HCO8yq0k6o+AHUYz8lOw2LcyOFDYtnySOOXXyfFzLOP3HPblInjI0LkjLVp40frf/XZR+/4ddg5Dinj0kENgtx49vX3Pv3lp2+/eaZBvVuWL12y2O26Hkj58O58tVG6QqWqM6dNmbRm9SqEa7fr4fytB5M6Z+K40SNffrLBPVnuoAM3/IIZGZnanRzpMzdMnPO+CnM+wUXiMOYHHn/+lQ5tP/vo03dee7HzV60/oY1YERYV3dqAtOn0ZasWP3zTrrXWHv05EzazIdXBT3bRO9RBeyNct8aZZ5+v9GNHHHV0zMgPIjPWu4llnlS/bv2HHy/nImZeeuLBekQFCRuuRMT4/UDeMG8zXcqjWLaXcmt03KjhCQmLVOaIPmrUPOcC1tQV19ape9YFl9ZijX7dusV7zrmWzTvGeLZmLKliT3nIEVLMxSNs1Cb4/j2wX+8zz7voMsYbr69k3wVSgUG+jRjy14DXP27zzaTxY0fdc8Ol5yjCSb9x9JMKvqTXavZh66+JjmlY7+ar3dSuoI3hg//sxzr/reuPnT3b0ypXP+0svn/+/muP9PujL9E6+QsXPjESSeWSXymFk9LgsOs7Ihb8x+CRT5epWKXKd20+eq51y09YOxl50tLYJR6kOXUJd1E0Bp/93Py+rgW7xiM75N3Ux0tnI60Jogxy7Fg+LDvI73iYzMgy0XPtrlfUBeXZ5S7NCj/NE/X8NEnhf9Mnm1pHKakUTeIvC6Un4n3j1Fj93fGKxuCe0gUJty0jS3JaVxSEojf8PmN9ph2JVif624VyijTxIyzUj5/6SnMhTQXZJf2o/6Jhcuz1tTTCNoYjQTQ3apOIAmmjqG7eIIP/1DgzslapnKI9FHWQGy5y6Cv1U6yoH82L5ow5JX0TERJaX9hHXcbMfc03z6WhIlF4X4OC8girU04po7CZ77wvvEvc5zN98E5SX6mxVFbrwV9LuY7dChgChoAhYAgYAoaAIWAI7LkIGGGx586tjcwQMAR2MQRIhULe+9YfvNlU5IFMXLVqRcQhR1olHPLxTH/p7U/asNu86dOP3Nf122++pBxtIjjL5z/7/vZLuO7K5cuWkoonXpqgbYUJB/qKZUuX4OxPta0y5StXxTZIhnBdSIcb6t79QG8nyDywb6/NxsXY//iteySSQkf5ytVq8HncyGFDXn7307ZzZ86Y5pzdd+NA5r6TaYjkZZfzM9wfzvExw7e0I9UxxSp/e/1HniB64FVHtOCEpQzjdqm0yk/+Z2zE2a8jESbsWCdK4c8+v/Wg/KPPvPzG0iWLFr736vNP8j2RiPGjz7zyJg7k95u98JT6wsGNs3vyhM1tSHXMM6dNjsy9y9yzRYTD+Zddda3ai7cG2Z2PvoKIHHQr7nrwscaM87euP2xyTpeMRlo4gmQznRfqjx0x9G/NtW8/7wcphHKb21TmiEgFiLRpk/8Z3+DpJs3afvLem5BjsXBLdSypYk9aqg/adPyZFG9pztueW33wpA6kRbyyyb4LVU8982x+r04/+4KLC7nQpEZ317lmzerVEe9r+EgF32vr3HkvKb0+efvVJktczji1xfpo+e5rL011+e2i9yJO5IpVapwxbdKECV2+79yPV8udafsddPjZlJk3azop9uRsxWmM07TAl19+ddRVde568O/+ffq+88ar+n3Zp0ChAyM6KMWLFJ5OOXfiaFV+flLmSItBBIbvEI6IB8fB1XempwUb5jnLXfMbF8hZ6zttRYjQltIwKaWS33xYrDu36Y/1XGsGR73SPokgEeEgsoKrUgj5JIAc5iISlXpIzu9wWiXsEAnA59y20Ps2JirrazaEx+qn26INjYXPIhchsvis/jSXmgfajDW/sinWM+FFm0qjRLmsYL9ieYP1c7ODfBHuUGQUREtuePhjC4+ZdpTKibZETPDZ141gHfMuQCpQh3GzxsCAZ/x3inbQo6AM/dCW1jt6JRJnV7oo5pQyGrNSYYm44D520C6DFrElXEWIpTJ+Hwv7bAgYAoaAIWAIGAKGgCGwhyCQ6x+2e8g4bRiGgCFgCOxUBEgbc9u9DzVi53HHtq0+DhtDfnvuDXXCuPEMRdCXlDv/a/Xxu9ohT9m7HnqsMbuciaJAWDdcf/CAPr24J82D7Q0Ezs2RQwf9uTXtQrSgLTB+9Ja6Hfc++tQLtPnuK88+nkzbOK1xaOLoLFmmfCUiUHzyh6gU2pk1ferkcHvoGuBMHzUsJwpjex4QAjfcfs8D/X/v2W3MiKGbxMBJWcW8i3hSn4kwQYCYckMG9u8DoXOh0/V468WnG2o3/zFOj4PnEEj+GGizUrVTz2j36fvN1zr9DD0j9Q+RCX17dvtpW8ZMRAGO5ROLFN9MwwIxb9I3zZk5fSrthwXGuYfzHx2E4YMH4myOHNfeetd9vDMt3moaWQMc4Fj33gaPscteO/i5z278cpVOqT56+N9/xRqD82VHdt8nmttU54g1T5tEVji+aMGnbzdrEg+/VMayNXPQ5K2PPy/nyLr7bqp1AQRKbm389cfvPSlT/cxzzo9VNpV3AWHz1Y5shVh8t+lzTyyYN3dOrDZTwZc1U6/BY8/MnjFtSqcvW7fIbTydO3dOq1jt1NMH9Pmtmysb0YJo9Njjx99+f8NnHQk26cF77mJt4ySVg5rPaROmz6nr1lih4QN+ezPaR55Ro0YdfN7lte8aM2zQ0GcaP00EnMS6tfOd9kUc4Jj1IwXkcM7N5JznBQ51+hWu+bSC/s59HLW0ox3uvgMYh7KiBlQn1X/HyxEsbQwRE1iEMxmyXJEo3BMpATmjiBONz48qwF5pM/hRDL7jGVtFUkiTQ33kFmmh8eLgTiZyJIcQiH1gp4gV7fSHiIKwke5DuCblRHrFcqbHs0lRDbQnwWs+5zj10wrkcWRFniA/GuWpH1EuXoQFDWjMIieYNwlkK7ICDBkvp8bEfMg+EQr+fNEu5IQILfoCR07aV9SFiD1fc0VROsJaWhf075Mo9MczvXOpvU+pw2c1DAFDwBAwBAwBQ8AQMAR2YQRS/UNnFx6KmWYIGAKGwK6LQC3nnCYPO6K32mHvW1uqXIVIjv5YhAP3yQlPyhdS43zwWpOnVRfn4hW1b7qN76RMwnEcRuH3Hl2+R9T4OucE3t4I4YjEcT56KyMTcKRPGDNq+Ib16ThDNh048tElcE7IHo7jmZaM3eVdPqy5rizEUKevPv/EpQDaLM1UidLlKtDOpPFjttCMqFL99Jo8Q4g6mb5SKXPuxZdfTTqcDm0+/VD1EBN+uulbH/3cuX27IQP79fHbi4cJZSBiuI4ePvivux9+/NkRfw/s3/fX/8iGwk7hmOezZ0yd4rcJOQLGPtGF2Dfi5c2bPPWoRK9TGVe47OwZ06eeWOTkYv59pR76uPkrz3P/mONPLByud+Hl11wP4Tagd8/ueoa9RERIyJ2UUm+1/Orbw1xOqdefe/whvw3WX0G3vX9kNOVXuH3mFiH2RBFAqc6RiCP0Yz5846VnSPMWD7tUxpIq/oisM4ekGQuv93htkU5s3pzZM0u7yKhYZZJ9F5gzlwGs3OFHHn3MtCkTJ3Tp/HXbeH2mgi8EF1FEnb/6/FNI2Nwwefu9D8vyfk2dOG44ZW+6+ZZjzqp104/uY1rXrz+rV7ZsGdrAMYozddPO+dPPu7T2uJFDh3768YekG8s3fPjwwwZPmPneIYcdefjogb2fc/fUt1Ll4HDV7neJZEsoOLcUPnK+/ufM369YWpCxKivIg392UxojOYm5R6SKiBJs4RmO4FSPsINdURO0A3nJ2uX3VzvnRVgoPZDGJkFt6om08UkBtSsHtZz4tC9iRMSEMNVYfOIk3vg0d8nuvg//jaM+/IgY+mLscqZjO450iY1r3jQmyidak+H5UbsiPBi3omeyguwNjrTKnxWsn0m74aiWZP5G84krjUskBGOAnCC6wY+sEMHBVeuYqApO6lJPkSCaX9rh/aEdxs99dGUOjK4FRQH5At2MSVFIYbJE7w1ryk+XpnaSneN4a8XuGwKGgCFgCBgChoAhYAjs5ggk84/h3XyIZr4hYAgYAjsfAZxwpKvp9n2H/8WypnK1087MyszMHOlywcd6/uTLb77PTvLGDerV8QkPxG4pz70JY0dFHHbhgyiDDm1bfkSe/xo1z71ge6IB0RJJ6bS1hIWLipC2hG8XAt6M97uvv2iZjL3YULp8xSrHOb2OvO5Li6iD3K9b3BEWEDra7e8/I/qAqITpzvGaTH+plDnt7PMvWrJ44YJBA/r2wrHa6IVmb3/Y7ttuQ/7s1xtHc7itCnEwoRzRI9IFuOCyq6/74PUXG/v1i5YsVZbvOJD9+9iAZgnExAknnVwMkXdEuls0b/r8T53+1yaV8cQrO3f2zOkIlvtCy8wj2iaQKqz/Y90EhesjEC58eIbGCJoW3b7vGHlXqp9x9nkdew4cWe30muc+dk+d2pP/2TwdFAQPbY8eFjvCgrlFYyHRGFOdI8S/aY80Vr93/+m7eG2nOpZU5+G+hk83IT1Szy7fxhStj9cekRgnuvxdsZ4n+y6wjiQs/sVHb78WKx2X2k8F3ytvcOSaI4B+/rZ9u2TwKFa6fIRsXLls8fizL7z0vLufeHFAmvsN6Nmx9bWtP/v0H/cIpzzOWZynkZQ0zV57/dgTihQtMrD3rxHx8QcfaVRh7tq831U85dQa7T9pXr/5G6+Rcsp3Vkt/QBoNpLPBEawUN762QzyzQ05Y5/PNcJItq0fIQax6cmhHhMbdgXNYUQFc5UyP1U+83f8+CUEZIilIQ+inK1JUh7+LXuNSZIT61Lhln1ImEQUiGyEClAZLfap+rBRR4fHEGov/d0sip3a8uooU8IkWnOwikrTLX0552eQ7+cGEwx+DX19tK1pGGKlN8KHPDUH6zMwg0y3PVcNjkUrx1lE8nGgzkg7NndgrLQ+RGtIAUX3Ki2DQ+EQk0IbeF8rTrnQoIC4oR1314c81bUFSMU7Nl0/G8D6y9riyDlkzilbyoyqMtEh2BVg5Q8AQMAQMAUPAEDAE9kAEjLDYAyfVhmQIGAK7FgLsDneisGe6HPuD58+dMyts3WGHH3kUzvRJTkcgVv53dqmffeFlV5JKasaUSTjgIgeORVJE9er+47ekUZkScuT6/XzV8sO3Sf1z1wMNN0VnbA+UTjmt5jkQLeNGDYspmp2oD6JG2DEfK53UuY7gwd4/Q9oV8dpzcgIVcJ5Ccnzi0vPEihigDBhJJ8Fvi3RS7NBP5HTdWrxISTR2xLC/Sb/UY/D4mTffeV+Dlu++/tLDd95Qi3RYfruJMKFccTeGiePHjLz5zvoNBvXv81vYSX9y8VJlGLu/zogCoF0iDF55t2W7H/sO+4cUTOgNtHJ6Kls7rnC9OTOnRdI+4cjmim5EzQsuuQJCBNJswb9zZystl7+GIZo6tWvdgnXEfaVwWudyV33+3S/9Wnb4+XdSXt1y+TnVGHO43wqVq52K0z6WNslBhxx6GPaMGpI4ZVkqc0T/RV1kAdeOjghMtGZSHUsqc0FkCToaP3X46otU6lF2sUvf5fTeC8XSPEn2XaB/2oJs+q3bZiLYW5iTLL4QXtWdSDtkni/Anmh8zt7TIDjOuujKh977ouMvQ/78o8+GBVMuer3Zq5B2OEpxFJMijTPi7F+wdEVE8yctyNrw5U+9utzzxEvtXXVulXoAACAASURBVATS+g6fNL/8o/fe7h/tT05oHKo4ZHGwck9OfO7xTI5opROK6FhE0/XIdDmx/9sRv2Z0VrBPkbTgoGpKc+Q7unkXsNVPsyTtDKWFCkc30Fes1EQiK/RM5A0OaPpRqh/6g5jRbnzZmgPV5ocfEaH0UtinXfpyjks/Adzoj6sfhSCbwo7teGPxrUiUGioeDtzHTu3ql2OfdjUmruiWiMzxHedqVwSOokp0349eoU2RFiICFMERre/0TjauTAvyH6FyPub+/Ibg3+wrdRWJo/VJP6xLviu6QRE6kAlK2aSIIZ988aM2aIM1rneBujz3CTCNSXPIVdE4It9Yx0R/EjUESUF7Sq+mqBuRLdQJ45ho/PbMEDAEDAFDwBAwBAwBQ2APREB/9OyBQ7MhGQKGgCGwayCAExnH4DCXez+WRYgS53GHc5jH1IF44PHnXsYZ2/rD5q+qPo75J196833u9+/9a/eLr7zupumT40cH4MTu1K5VizsfbPQ05Mi2iizLjmqn1TyXVFS+LkKyqFc8pcbplB0ZciajXVC2YpVqaD4kkxKGNspVyhHcJu/9d+3bfBa2gV3/kCN9Ymg10B9z1D26oz9Z+5MpR5+OKziZ88xzL7z0ly7fdfjUCQnHS3MVDxP6gpQq4kSyiUi5+qa69R68rfalYRtwYIdTXrld42dQrl6Dx59hvXz+0VvN2n36wVsQQsmMIdkyGhMEAUTKJVddfzN1e/6Us/ufXf2yRW3We+jxZ1g7OP51r1LU3pfe+aQNbTZpdP+dXb/v8JUIjbA9YPb3n3/0jmUn0SqRNZZAYyXVOeJdZh6IaurxY+f2ifBJdSzJYp2z5nN0NMaNHjE0lXqUhUSFuMtyoPp1U3kXikWjTHhvEr2nqeBbpcbpNcF3cP8c3Z0kjmxH3J6JiDiROm881+iub9q26urq+Smb5CjfFDlwbOGiEezqNXrurX9nz5zd+p2mjz9cv167a99uTj0dOGpxbuNQpS7Od6X+EnmhHeE4aOU4juUs33K3eOa6PMHKodnBPkdnBvsVlYaA70gWIUI0Bw5ipeNRn36KJDl9w30rJZGc0LJDTmXGxz2fdJGjPNGmJjmVKcvfEiJYuM89SBgc1FwZh8SVfRw0Vt92pe+K57BORFIkWi6yT2ST+qGOyBSluZITX+3F6tMnf/zokzBmGptIKfqSEHnBYL8SacHq8S4t1H7JrZnYI/SjIxQ1gR30I8JCa0aklMgCEQdcieiBNBBJJk0LETeKqgAnRZlgkR+5IcFtrS+RQLTBOuCq9FOUJdKCd0rkHHbY36aJVrI9MwQMAUPAEDAEDAFDYC9BwCIs9pKJtmEaAobAzkMA5ya9x0v3VLvO7ZG0QONHD9/C8Vj11DPPJpUTZIMvpFzvwccac/+D115szA566pOSJ9Eo23/x6Qc4fa++8ba7tgcaOAmdA/r0rdevqHEaDmnEmn17SpevXJX8+MP+6t83WTvLVc5x3hIxEMt5Ks0BpwGyRdqssk6wmf5IXZRsf8mWczrex1O223cdvrrizApFn3vkntsSaXJUqBobE9o4ya0jnLkVI7ofI4eH03AhXn3o4UcciSaIb59seMeJl19creTxLd569YXtTVbQn1JtuaxcRfle6/o6tyPmrWiXqY6wwCGOA5vnONyJHiLt14rly5bKZvQL2F3/+L23XntVzUrF0UaIR1Yw5hOLFC0ej5AgWgBiYeK4MSPjzVmqc3RyiRwCcnD/vr18u2O1n8pYkl1TKneIm2s+L3URDqnWPfGkosUWLZj3bzjaKJV3oWTZHD2Vnl2+65io/1TwhaikraGDknv33dSfBMaOrI1EnrmAJRyeEA3aBc5tCAty7eOQ5XO+gw894ki3xpa2eO25e04pemS1j95548sSJSJ68ZRRqhv+jYzzViQFTlo5hNE5kDiwdAlw3MZzqIsw0K53p1/gihcs5u5ny4nPM8rJmYw9h7jT3/nvkxSC3Xeecy8cESAiRbv4KSMnt+ySRkE41Y/60A57XbkvwkF2KzqDtrgXEedwhyI21JauIj30XeSH7AuX96MAwtEHvl3hempPjnec4/4ufj+Fkp8iK17/sezDHjndFTXnEzF+RIaEpjcEaydkRnQs1kdeYc2z8EyGnAlHRviRDyIjRLYp9ZhILOaPtc37QtSDoidY27LHF8wWMSFyS0QX5J2IPkVUCCPuQ1T4KZ9EXiiyx7eHPvQ91jzaPUPAEDAEDAFDwBAwBAyBvQQBIyz2kom2YRoChsDOQwCnKr3PmbmleDSaEugS8HzS+LFbiEHj9OXZd1//FzUAUXFvw6deQBeg81etP3HBAeVJS4OQbqJRLl44fx4pdc5yaXq2BxqV3W5odmqPHh5bOyC3PnC8x0rVgwOaurkRMH77CG4TPdDzp+9i5vIvUapsRHAbR3/YLlJFxXuW2xhye36wS0lEmR4/df4mVjqwcP14mFCOeY5cXYRM2xbvvhGuS3QF9/4Zu/kYZUOnL1u32JpImNzGqOezpk+dzGe0ESBXICR8IeZpEyegCxCcVDRHGPzRZ195E+Kk3SfvN/f7wF5IHcTiY6Xv8ssqgiJeyieE1qe6fhOJYqc6R24pVcaG3r/8/ENu2KQyltzaCj9Pd4Is3Dv0sBziItkDUsvhUjGW5kcq70KpshUrL5g3d05uYt+p4CtdjbmzEpOvGmuZilUiUVq9uv/UeerE8ePPu/yaW9xX7QBHY4IIgnD0wEanJXMgvy+fffx+lyOPPBKHOlEM/E5DbPDOHupOyAIIDE5SBMkBT5dyBssp7TuHs1zAXDiiQmLCftobF4MwLjtI/xcHrRzlik6gD+zCuS0tADnWRXrEE3/20xYJKqVAku26v2XkR+yFJGJDVznGFbmgSB3tsIe04AAzTj33Iyc0HpEPimSJRT6ESRgRDj6REh6bPxJFfijiQGXpU2mxuOf/XRTGJkwgyAmvufV1HNS36vj2Rt5bd2QFhcrmDfY9KU+wYaH6ppxIgs2in2JPS+SuMPCJLX9+WD+KXBAJx3fmhXli7bPeeaY1xboT8SISgTqK+lEEE+ODBNR8h0ko2hBhwTNIEU6ib7j69mjsPlYJhm2PDAFDwBAwBAwBQ8AQMAT2ZASMsNiTZ9fGZggYArsEAgULHYDjLJI33jcIoejHnn/1be65/OnpOFbDBrMDfeK40SP/dR5cnrE7/d3Pv/nRbaqe/+JjD0QiJXDyIcScyCmrdkm/dLzbAS+x3G0B6LSzzruI+vHEjhO1DdGB03TksMEDw+Uk2rzIESzJ2Efeexzkf/b5tUc8DHDys0t/6qR/tsCYdFAL5/87N5YGQjL9JypzoPPW8txt8tcu7bjFE2FCJaXgIQXXX/16/xpuSISF09se6z/7z4b1udqwLeNdunjRQpd5bBmExJXX1bmdHfy+nRLLRvsAEXqih1q81fQFNBDC9iazlqlTsWqN06kfL2qFuZ02eeL47TVHtFOqXMUIYTEwCX0VsE92LKlirxRwZ7hUY6nUvemOex/it0ei5n7dZN8F9EkQFE8Wg2TfAd598GIdJTMmBNcpN27EkP6OkPvA/SZdUOua6yAxcKRKGFqOWJELG/c/6OCDNm5Yj9PVF8uWw1epcBTtQDl2oWsnOZ/D6YwUFRHPyRzebZ/jDM9YlR3sVxgbaJN+/VRLkC0cECY88x2/fjRCPKh8ksEvo+gTnzxIBm6VEcGgyA0RK9JK4Dm2Q/Lwmd+dcOSCHxWiv0WEkZ+WS31qLOFx8F0OdT2LR8IoQkC2+DoPIoaESaz+aN9vm3GLbOKK3SIHwngq5ZeiTXK+Z67IE6Q53mB5f5908NdKwnlxxJiPj0gKrrSv6CCJqcsG8NYa1phE6LDGmC8RF/64tLaVmoxy6lNrkzK8J2hVKKJDKZ98QkR2i7RSdBLffYIkWUItIU720BAwBAwBQ8AQMAQMAUNg90PACIvdb87MYkPAENjNEICMwGTno1eqhcgIbqn3wKM4oREUdhvKp4QFmEn1hCD3GCfWTXkc8++36djFbUA//Mn6da9XOhqXEuWEWM52yI3CJxeL5DnRkcelPoqmrk9292ZctCFT5v/rwjqcmHOqU1KmQpVTcJrGIjvyBDlemDBe3Ctf+ZQaBfbZV468SLcujcwpaIAM6relILPsQqwapzZYh21FkHqJY0c2YeTaQtA81THFKr/WhRBw35nMLtSERyJMqCiR485ffv5JrIaKlixVlrmd7gmzUy4VG3KzMbfn0yb9M/7k4iXLXH7tTbf92PGrL/xUTghjYx9pfx5v8vq7EBgd27X6ONwm9jq4csUrsh5cyqdEhBlOdT/lGO+Q0oOp31TxIRUS0SREF+SGRypjya2t8PO/B/brjQ03OQF2CLtk6hPNdfv9jz5J2rD+v/+C1sNmR7LvgqLChgzs1ye3flPB1734eUi3xW+D3y73Yr2TFapUj6T8mjF10p9rlsxrO3n8mNF3N3z2k1pXXonDFY0WOWDT77mv/mHdu3dnd/uydWtWr3a/LzjUyaevnd84R5UeB0csddkJzsnha2GI1JAuhnajRwoiuu05k7nlO6H/26m/2mUqS59DXXao+79N/o516ot8EUmQWwokv8/wFPnpoFQut2n0Uw/x3w4/YiJMtPBdjnwwhnCJd6hdOb6Xu4KxCIsIrF4j+ixiSo5vEQ1+WUWBiKhhDTBvvpMdLQVpS+SW2svHns9yyDNuzXN4vH5qJeY2J9Jj/YKMYO0/2UH2Ji7Ztz8c0ZEIQ41RJIEflSMxeK0j/h0C6YANIi9EgMl+1VFkjp/SSSmtREBQF0H7xdG5o45IDaI4WAN8Z5DYBf4S4RaJJMxFtoRTfiVYQvbIEDAEDAFDwBAwBAwBQ2BPRMAIiz1xVm1MhoAhsEshgKMWg8664NJaMqxytdPOfOipF17964/fe+KMi5UuSKmklrvwCXY0t+zwc68yFSqf8kKjB+4UiUF7TkpiH+d/izjG/eOZZu+0aPvDb3+SAob7hx959DHoZYxyUQ04+bYFpOpnnH0eO/r/7PNbj61pp0r102u6jDZriBYI10c4m3tOgPcs/9nt9R954ssuvQeVKpeTkkcHmPB5aBzNC5yf6A5IYyHcH8+d7xLHZeR47vX3W7bu1L0vzu2tGZtfR2mSFB2hZ8c5oQdE0/3d8YkwoV7RkqXLQrh0/6Hj17HsYj5WOi0IEWQqI0IpbANr8JV3W7Y7+rjjT9zWcar+FEdCEL1zuCPLvm/ftpXfrjN97VxHGl1x3c11IRLeeP6JBrH0RrCXtGBopKg+GiOX177x1iZvffy57iFCXr5ytRr+u+D3R500x9BpbpnPVp269X7hzQ83syuVOaJ9cJwwZsSwZDBLdizJtBUuAxn08hMP3b2vY3dad+7et9rpZ52bqB2Iohb/+6FnZkZmxktPPFgvVrqtZN8FCED6cinWcsUhFXx595k21qbGwu/jm5+269Tymy69eKb7rI9iLk3auJHDh8ycMX1tt27d1r/yVIO6Rx973PHX3PHgT680bUp0E79zG+vVq5fnjoZNev/4S5873fcC/86eMeO4wkWKTJjwD85XCInFS5cuTa/foNEVr3/0eTP3Hacqv6nKsy/nsQgNrpxywvoO/VjTIIes7wzPCtZNzxOkz1KaqPBvsogFkRQ4urX7nKtSQyWa9lhO77DDPZnlp3Zkix9NINJGpIHai+dw953Rwo26nJBCEjAPExR+e+G2w6mc/OcSkta49btCHeaf5yKvlCaJMcTb3S9SgXGI5GC9cF/kTSxM1R945UR35DvElXdrOnO1nxbLXyu5zk2UGJOjX+vCj+jwI0pEqmCDooIkmi6SiXH7hA420J7WvAgrRWkwbv5bqY0Efn2ljgInMOJ9EjmkFFMiWbjSdm7vUq6YWAFDwBAwBAwBQ8AQMAQMgd0fgc12sO3+w7ERGAKGgCGw6yHAzn92eTd8rmlzlx3qQMcv7Fv3vkceR3fivVeff7KNIxWcT44diJsdpH2izA1173mg9s133APx8M7LzzzWs8u3m+k0IHp9as1zL7yvYeMmLd997SU1gsYFqXdwvs9weXFOOa3mOTh5n3DRGduK0n0Nn25CG6edff5Fr7do0wFHI6SLi1RYgC6BE7/dyJhcUEmh/fYrVGj/Aw88yPElxw3o/Wt3HMzFSpUut2L50qV3uN3e51x42ZV1rzo/ktqFo3/vX7ohusyzNatWrYTUuKhW7RuuvqluvWGDBvwRFpuGsCDCJF5aoMJO9Rzn5jon4BBr3DiVSU/04JPPNyUlDpgxL9tDmHrG1MkT2c1++30PPz5/7uxZOO3PvuiyKy+75oZb0JMgCkE2JcKEdFEukKbwT658vNRVEBbgFh6jy+//3VOvNP/w6Vfe+vDTd5q9SJqiK669+TbWzKTxY0atSjL9TjJrZnzUgd33t+5dYpFwpEU74aSTi/3ubGIuY7X5i9P7uOSq626GWICcKexSTF1/a736RYqXLO3jddyJhYuAi9MjOLh99/7DPn3n1Sb9ev0XNYBD3skUTD33kiuudpFAsy68/OrrIa7uu7HW+X6/qcwR5A7k4cihW6Yy25axJINtrDIDHeH58J031Gr63mdfftaxa28iHn7v3uW7CU7HhBRdjovLRwq4Cy6/+rpa195cNz09fd3TD95xE2nmtuVdIEplxbKlS5KJrkoF3y7ftm933W316r/0zidtPn7z5ecgYuvWf/hxyLxW77/xik+yEFHE79mIIX8N0FicRM2ohnfXuerd1u1/coFTf9V/9MmPFs+fO+H08y+7DcH3FUsXTXdl8436e8C351561VXdu/7+ylvvfdA5Ky3/sVfdeNs99Z96qWT37zu0d2XY6a9d/3LAaue4hITlJKecyIOIszWGhoUc8nIO5zjUs9Y68e2NGUFWZnaQllcOX9/ZTtuqi0OX+qRQw0FMqsGk0wdFxyONCV8nQA7tZJahH8kg5zgkA3ZotzzthNv07fTJBY2VKxhK+Fl/nyQaH1iLPKDP8Hd/PNjo20c9OcilnSBnuZz6ifCQU53/bovU8nVCYtWVg55naW7ONwYZKzOD9f/6ZRXpABZJbypjvblDBAr9SAheAvSsLWGsdFH895D72C3ixV9rPjmFjYrKUKQK9bT2hSdYKNWaUqxBAtE+ZaQpA3mh9RMpF+OdSYS/PTMEDAFDwBAwBAwBQ8AQMAQMAUPAEDAEDIFtRQAn+N/TFq8fMXtlNmf3v8bNkAbEB207d+V7rD4aPNWk2YAJ/67s0n/kZHamxyrDbnSef9Oj/2aC0uQkeerl5h8Mn7Uia8j0JRvYoVzc7Q7f1rFQv3OvQWMGT1m4TuNJ5sr4z7/sqmup/3Djl16nzh9jZy3FOR22iXJ++4wBp2xBx32Ey3b67a/RP/4xfGK8cZFKib6efe29T2OVcY7Nk3uNmDKfMoMmL1hbr8Hjz2wPjNRGlRpnnDVw4vzVwoj5fMqRB6Ts8vtJhAmpwXoMHj+LlD2xbMNxO2zm8sxmH34eM/ritnsbPObPEW0RseJHMWyPMZOiaej0pRtJ3RWrPdZ675HTFiaK6mDdvvdFh598e//Xte/fWjtq1wVMHDR46qJ0yn38vx9+gbiIuY6iZX4bNunfeHoPyc5RzfMvvpzxJRuVkuxYthV7xl6/UeMX+R2J9S6yrt/8pF0nInsS9ZXsu/B1tz+GEImUrN3J4kt7ELv+GP6atGDNnQ80fCrc18VXXncT5ZgT/xnpmFywyekde/45ym/niSavveueFXTnwUuWLDnwgzYdu4bW2JAbbrvzVvd8/2i5fdy1gDsLRc8Do8/2ddd87szvzrz0Fz7Dtmb3Co5wZzl3VnZnRXdWcGelyHVqk9LZG5cXc20Ud2dpd1ZwZ5XoWdldK7qzUvRaNtrvCdHvKpfoSl3aLOLO4915YrSfMu5Ke8m0QRls4SwfbY82i7qzVPQ7dvI8UXvh56qjKxiABW2rvzAesiVZu/1yjJe+uDL+k6N9MSaw5wpenLmNBbvKRds42l0L54InbTIHJd1ZInvjyuLZ//6vXPaAIqyHnLWQszZYI6yVI5J9vyjn2oykInNnmjtZm6x11u4h7jzGnce5EzuPcufB7mQ9Hxm9d2z0OeuDz5RjnfCZ8tTlu07GyueT3MlnntPHEe48IFqHunw/zJ2Hu/Mgd/JuYRPvj96diN2pjNXKGgKGgCFgCBgChoAhYAjs+QjYPxD3/Dm2ERoChsAuggApmUqXr1iFyAknsD1WYrzsVkao+Nefv++0LaaSziVWih12FjuHQDY7+relfb8ujlja5Mou931dKEXkui9X9z93JcKC1FNEFSAKzo5vpaKibKVTTj2D9FSkhopl1xFHHXMsjk68GaNH/D1onpPLiFUukgrJRQkg8hxvfOTcnzV9yuR4faXlzZv30MOOODKSUsmJ/m4vnNTOQU54hJQ86W6s7H6PZUcymCSyCyf6WrcjPZ5gMTvtnb5EaadlPnfShLGjfX2J7TleUi/Fi05hTjPdImUt5NZn6fKVqjqe5mh26CtNWLgOYurZbtt9rNRiKovmCQ79ZS78J1YapFTmCMKI1Fz9f+/ZLTf7/efJjCWV9hKVhZQgkiQi+L1+ffriBfPnTRw/emSy738y7wIRQkRLJSuOjb3JvAMaF8RqCacVsnrlyhXDB//Zj0UdHjORLtXPPOf83r/8/IO/lj3nZ9opNU4re8jhRxZZsWzJ1L8HDiDVHLu6lYJpY6VTalRyr/3R61avnDKw/x8z3DPt2FfaG+04125z7RoPp1WK/Hs63i5x53w+yj0+3J2KHJC4cHZQ5LmM4Ojb0oKCJbQLnWfaEe+nx5EAMil1GAMpr5KJlNYueNqfGx0jv3EQfJxEHyjiItaufkUuyBZFnkjDQHW0sz/ZqA/NhaZW45OmB+1orpL5e0VzQln+m0KaJ9ms+kQcgK1SKIED4/d1NzTeRK8ZzxTRwNqkP+YYfYh4tjJeyuVEJqydXCBY+WcQTH89b7A2wrcrYoHPRFgsznNBJJom6cOtfcrSv9JPhTHUelG0CeUUxaMIDM0fERXMBVETipgRxnovNFZFp0irQ6m2qA/Gen/89wZbN30Pab4kPWYraAgYAoaAIWAIGAKGgCGwZyKQzB8Ae+bIbVSGgCFgCBgChoAhYAgYAnsEAlFnrT8WOW65p8/SB/Ad837aJTlRfWJCbcYSAt6kc5DI4eoIi+NdI0SHST9Bzuns4JBz1wXFmhUI9q+W5dJCqQ8JfCvVkpzIPId4xqENAZJM2iBpDSxzNi6KDNDtbneXE6I2+aLMPn5y3EtzQc8kwIwjmv4lIi2c5ayOta6EdfgZfZEmyCeGwACnuZ/2KVabm+Yg+lApi1RW9SknRz12cF9jULqvWO3HG4d0IMADO5lbpZdSHd82+kMI3qWDysgOlv9RIFg+IDuY/qLGKBKLuti12hEWc5I1aFOH/5EWGrf/HtCXyBqtHT0X9hJUF4mj9FQiI0ROiOSia6XD8udXeKs9fx58XJRGLdWhWnlDwBAwBAwBQ8AQMAQMgT0YgWR2Zu3Bw7ehGQKGgCFgCBgChoAhYAjsgQjIAauhyXHK9zD5QFnpUIgcoNym3fbbmGNffftRCTk2rBzkXNMTs4KCpTYGaZGsZtIz8h3O3NcmIxzjaFgkQ1YwJogAogpIb0Ub1IU8UXo9iS2HNR7oMyyCLIc8u+6pR7uyQ5oQECRENyTSgghHPoggoi2JbtNOPDIlvFx9kgKbEUw/KGq/nOn+Ji1FHhARsTWHiCTGiL0SuQ5vBNNa4go+kDDpQdY6J7Ttgi3WjFGEgdaZNCyEfcq2RYkzAiD9SBERNFr3+u63L1upxzxgL4dPIvnj86MlWGcqGy6jPvxoiqh5KQ/PKhgChoAhYAgYAoaAIWAI7CUIGGGxl0y0DdMQMAQMAUPAEDAEDIE9FYE4EQ7h3fe+83QTFFFHfrisvsdrIxUoceyza55oBJEW1M8KMtdlB/mcf3/FwDzBYZepTZEHfnSBnMxhIiaRHfSFODfOZ67HuVPRANSTiDafFfWhnfNhgW7dF4nhi4RzD8c9JINSCfnC23Ji+7vyZTe4KL0S93B+07aPQaIx+o52bCaKAcIE8WeRH9QHt+31dw99Mk4fM5Em4YgQ2fdfuqT0yXmC9XMzg4Xf+amZFMnAPTARvonGHveZiItogU1rOJrJcbPvMRrxyT1hl6wdIiY2I2/ChJ+lgEoWTitnCBgChoAhYAgYAobA3olAMruz9k5kbNSGgCFgCBgChoAhYAgYAns8AjhTcaBGTz773yP3t/Zw6aBEUCgdD45p7UjP0XGY9pJzrueXo9/f0a7IDz+tTyRaIgV7qEt5nPXUxYmvtE3SMKA5pfPxd/2rf55jM4QAdaTVIAJGUQyKNuB+rF38cpQrLZFSdFEfm4j+gGygD0VIJEMYCR8iPyAquIJnOGokmbaSgdaPXvDTQPkEkNqR858r404P1s0OgkU/+pEtwheMuY/tGW7t+KRPMnblWiYGcaD1vj2vET0X/8zVMCtgCBgChoAhYAgYAoaAIWAIeAgYYWHLwRAwBAwBQ8AQMAQMAUPAEPj/QYB/ayPMTPSBUvLgVP/Peb9mbFawrPeqICuTezzzdQUUFaBUPck63VVe/9anHRzh+u7vhBdxAALSqFBKJ0UGiNBQmiYJg1NHhAV1SDVFhIBYnnAqJsrTN3honNKBoA8/0oAyfuqheDOkMtKigDDxU3up3tYwT/HwjjU+jc230ycdmOP8Qdo+G4Olv4qcUB3mnQMMGPcWQvPxBm/3DQFDwBAwBAwBQ8AQMAQMgT0NASMs9rQZtfEYAoaAIWAIGAKGgCFgCOwSCDjhZBzTOPJxSIsM8NMEYWfeIH1q/iDbiTHnEAoiN3ySQv9mF4GQ2/jCznkRAdgS1pf4TwQ82guP2gAAIABJREFUh3zw00IpGsInF+hbjnxfvJn7iuiIFx2gdiA80JoAlxXRPqUtQdtobyiSIxmiQWmlqAN+wj03nBI99yMpwuViRVPEKi+SimeOSMlYH0x91hcy13wqpRRrBEzyubUTTs20LWOxuoaAIWAIGAKGgCFgCBgChsBug4ARFrvNVJmhhoAhYAgYAoaAIWAIGAK7IQJKAYUTHgc14stKEcS/xfMFCzpnB4s6EwGBs53UShKiVoooRV7EEzWOB4vSLSkyAltoS450kShy8itaQamOlD7KF8amr1iRE9Jv8KNCYtlF24wVcoGriBlFekh8WxglmnI/AiNKCmzCbluXSqwoDV9vg/b9CAxhImyxn/RUiibJCma9mSdYNZxyYKSUXJRjTTBHrBEOrZltHYPVNwQMAUPAEDAEDAFDwBAwBHY7BIyw2O2mzAw2BAwBQ8AQMAQMAUPAENiNEMBhTTTBYneuiZ44rKUJAYGQGSzvJ8c9wtHawS+HvC+6HS8dUTxIfHJB2gnaya+d/UqjpLLSr5DzXRETYVHpRNMQy+Gv8hor7R4RxQKbOMBLUSCJogxEFlAPXKlDefQvYkVAbM2SCRNEtCsNkXjpokREKNqE8hAQC4OpL3DFRuacctiO3VoXrBHWChjYYQgYAoaAIWAIGAKGgCFgCOyVCBhhsVdOuw3aEDAEDAFDwBAwBAwBQ2AHIYBj249k4N/f0nnAeY1De99g6R/pQVaGdt/nkBg5O/hx6hN1weELZSdjvlI6KcJCTn36kdOcfvwd/YqmEGkg0kJkRW4pmmJFX/i2KnWSyikNFXag3QBWctgn+ltF9oAf+HAq5VQyf+P4hAOfhXfYVn0XueN/jxfxItuUCiw9GFtndbQPCacrooS14KcCY/zJapUkswasjCFgCBgChoAhYAgYAoaAIbBbIZDMP+Z3qwGZsYaAIWAIGAKGgCFgCBgChsCugkBUiyDDXXFE45xWWibtsM8hIdZN2jeY+ymO+oiGQdSJzTDk2M6NKAgP2U/v5DvAsYM2ScckJ72uSkGllFA+ASDhbfpRe6k41v30TYo0oK2ctFg5xIxSZhWK3ve1MBL1BWnBeHT1xcVjLQVFrOiZxhkuG8Y81t9OPqGj+hor9oPtimDBN6TA4hSOfoQNeLA2uBfBJrtXLLPtniFgCBgChoAhYAgYAoaAIbDnI2CExZ4/xzZCQ8AQMAQMAUPAEDAEDIFdAwFFEOCQl8g0ugU4q4NgUgP+H4e1IiPk1I61k1+Oco2Meorm8KMY/LqQITj1caRzhShQPbWndFUiCBTV4ZMAflqqZEiLcJSGdCz8WZFDn3s4+cPpoMIY+DofGm84FVQ8kidWuqpk012FxxsmRyRwLtKCFE8IizM+DuZaeib0yVpgnpc7UitycNVnHyD7bAgYAoaAIWAIGAKGgCFgCOwNCBhhsTfMso3REDAEDAFDwBAwBAwBQ2CnIeCczxEnd/QKWYAYM05qSAMc2fybnHPfYNrz0jhQyqZwlAHlpAGhVEbSpuC7L3od/re+xJ0pI3IDO5ROCTNFJnD1xb7j/d0QJgXiERgiIEReaAwibrgSJeETJ4kIB18rIpyGKhYhoVRLseyLZ3Os+7HG65MrSrvFHHMGwe95mGNSQWme+c7cYxNl8obWyE5bq9axIWAIGAKGgCFgCBgChoAhsLMRMMJiZ8+A9W8IGAKGgCFgCBgChoAhsDchwG57kQLstI84rN2Joz5/ML0pjmx25UtDQqSEMOI7RIIOOefDEQi+s92PHqAvaVZQBpJAqYhoU5ELfMbJrkgB2RFPt8G3R+3QrlJQ0S52c8o2vy9fkyL8N0o8QoGx+MSHbPNTVtEHpyJHlHrJJxliERyMIbc0XH4UitI6iXDyx35AFGcRS8w5cw/2jJU1YYchYAgYAoaAIWAIGAKGgCFgCET/gWxAGAKGgCFgCBgChoAhYAgYAobAjkEAMgJntUScpaeg9E8HBn3yyxEu57eiLKS1AKlBGdX1SQUJfMdytitlEhEV1BWZoKtIAz/dlPrEyY494WdCLUwSSBdDZABEBW34JIWfwkn1FXEhMoL2ExEHIjd80kHjoE2l3MIe+scOEUX+jOdGToRXh6+DIeIHXKVDkqMRMvIyiJID3SnNkvC8Ywtrwg5DwBAwBAwBQ8AQMAQMAUPAEIj+w9mAMAQMAUPAEDAEDAFDwBAwBAyBHYCAS/0jhz2ObZzaSsdEuqacZ1kZaUFmOo5snOyxhKdxusthLs0EX5wbpzgkRPiQU14RHvQtgW1fzyKs58D3sKB1IrTCUSES1pZ+hk8u+EQFbfp9p0oi+OVFrIAf95e6898Ivjlj5ogXuREeW6xyfhvMB5Eb9JETKQNxkbk2T7Ckh+abK3OMLeCeU8bZEF0TifC0Z4aAIWAIGAKGgCFgCBgChsBeg4ClhNprptoGaggYAoaAIWAIGAKGgCGwiyBACiCIBjnnRSAoRVDBYPY7a6IObUz2Bab5TrlwhIXa8iMTKBvPKU+0AXWktbA6+p060sEQXGo7nHIpFpwqi42KJggTFooIoX4iUsKP2kg0lnA5tct9yAHIH/BGO0KpmnzdjtyWRaxxMydKLwVejFHC2jnppuZ/CZEhjRLw0PwKI2yydFC5oW/PDQFDwBAwBAwBQ8AQMAT2KgSMsNirptsGawgYAoaAIWAIGAKGgCGwsxFwO+qVEkrpm5RqSY789cHcT/IF2Vk4thVNIae86jAMaVHgPA9HDShtVDxCAOc55EahaF3aVfqnWBBJ7JtnIkt8IW2RE6orvQZpcejqR4wobVRuU6IxxBtLrOcai0gDxgl5AFFBpEOyfwfFIle4B1khHERc/DdHWZlZwT/3Y4PK+ZgpHVee6FrIbfz23BAwBAwBQ8AQMAQMAUPAENhrEEj2H+p7DSA2UEPAEDAEDAFDwBAwBAwBQ2AHILDc9YHjGvICZ75SOvHv832DDYvzB8t/J8rCJyL8dEaKulDqJ8gLX0jad7THG47EtnHgIwzta0rEq0M/tK3+YkVBSOSaNvy/N/yIEr/9eFEgyaaEilVf9xQtwhghS5SGC7tE+CSa7nB6LMYmPQ9pfwgPkUsZwcJvmDvIEYTLhSvzgz3MOe2wBuwwBAwBQ8AQMAQMAUPAEDAEDAEPASMsbDkYAoaAIWAIGAKGgCFgCBgCOxgBt7PeF98WESHHd/4gK71AMOPN/YLMdTjH9VyOb98B7hMd0mvguTQuuCqSQboO2u1PFAZOderJoS8kYpEAIkloD2c/9RTd4WtR0L/sor0w8aDoB/9vkWQIFtqKl/4pPIN+GifpgSgFlp9OK5mZV5+MlXEvdqdIB6XzgojIwTf93w3BuNsgKqT7IZJHUSrYsTa6BpLp38oYAoaAIWAIGAKGgCFgCBgCew0CRljsNVNtAzUEDAFDwBAwBAwBQ8AQ2MUQQDcCZzjObzns/4uiWNprv2DNSEzmnp8+Sc54HOI+OcEOf0VZ6L4ICxELXPVZEQaxUkGFSQbZR1SBH+lBP4rykEMeG9R/LMj9sfJcKbFEiMSbJr9ePPvCRAtEwkHuJLICEoFIkkQppsL1+U55sEIkG7ICckcY8EyRFsxHZrC0O33RD4cwke2aa+beDkPAEDAEDAFDwBAwBAwBQ8AQCCFghIUtCUPAEDAEDIGdisAhhx1+RB537FQjdoPODzr4kEMNp22fqPz5CxQ4+tjjT9j2lvbeFpLB8EC3YDn3XpSSG7nbYU/0hLQjqITeAb+HOPCJXsgMpjyTJ8jcKIHusKNfYtY+iaAoC9qTU11pkfwIC0UGUE5i0IkMl0aF9BewXe0pbZKc+3LSx/tbQ8+xG5IljEPYDkVEcF92hIkF2eD/90SfRahAKPjRHSKB/LZiERbUh6zATiJS+A5pocgJ4ZARrJ+zOpjUEDz/m8OcPplb2b8xOvfJLRQrZQgYAoaAIWAIGAKGgCFgCOxFCBhhsRdNtg3VEDAEDIFdDYG8+fLl+3nAqCm313/kiV3Ntl3Jnnz58ufvOnDMtEbPN3t7V7CLeevwy4AR51921bW7gj2p2HDrPQ827PTbX6NTqWNlN0cgGQxf++iL9i++3eILwy4pBJa6Uji3cdwrQgLnNv9OTw+W9c0O1k5w1IATcc455IRX2iXu4USXyDV1lQ5KRIXqSXfCb4syOOJzO3Dk0zaECI5/6ol48Ov6Dv94ZLQiRqjPmDlE3FAnFhmhv1sUISL9DerGIhx8kgN7Ofw2wEJC4GE71YfGRVsigg6M4k2kBPeUGistyMrICub/b/8gc3XO3OX0B2bh+WXO7TAEDAFDwBAwBAwBQ8AQMAQMgRgIGGFhy8IQMAQMAUNgpyFQtETpsoX2P+DAgoUK7b/TjNgNOj6paPGSDqaDNm5Yrx26O9XqIkVLlCpZtkIlomN2qiFb0XnVU888e/XKlSu2oqpViSKQG4Zp7qhU7bQzDefklozbaY/DXpoU/BZK9wAnN7v48wULvskKsiM+eUVS8Nl3visNFFEAcs4rGkNtUwcHu6IuuCpCgDqJogw0mIIRe3JSWMlZzzM/XZU+y75EKZZEzFDWt0EpmHwQFb3h63Rgv8gFjYU6PuGg6Ap/7Iou8YkK2akUWrTjEzwigSjHnPnRGpAT64MN8zcE01+nTTBi7sCCaAvKMreR6I7onPtjs8+GgCFgCBgChoAhYAgYAoaAIRBFwAgLWwqGgCFgCBgCOw2BkmXLV6LziePHjtppRuwGHRcvXbYCZo4dOezvXcHcStVPOxM7pk+e6LZ9715HuUpVq48ZMWTw7mX1rmVtbhhCREJCjhkx1HBOfurmuKI41iECFMWgdE9BsPKvPEH69AwXZSFhZ0UP4AxHC0G7+OXAjxXZQPtyumMZZeTExwGvunoWtl4pl6iDHfStCA4iPBQZoasIAKVwUnt+BIWf4or21nhjCffvEx8iaOhf0Q8aC+PQeMJRFIm0K/SMdkTyKD0X2HG/kDvpm/EqSgTs93VRFU5o++aNQeYKynEoAoXvlGFuaYe5tsMQMAQMAUPAEDAEDAFDwBAwBOIgYISFLQ1DwBAwBAyBnYZAidLlK9L5+NHDh+40I3aDjkuUieI0ZsSwXcHcilWqn5btjonjRkfUgHeX4/jCRYoedMihh401R/pWT1kyGJZ1pBAdjB1pxFCyQLsd9zi/IR4QhcbRTaSEhKizg/S5jk5YkhWsm5LtSAuaFXmgNFDcxDnvC20rIkFmxCMO1JbKiQyIZb6fAkqkidJYKfJARIjq+yQJ90Q8iBgg+gACgH5x6CvVlRz/1FEKK33W3zB+9AjP+O6f0qvIbSpEnNC/IjI0LvoW+eCLg2uc+VwqqJXB7HcLBcsH0I+IE0VqMJfUZ25XR+c6N3vsuSFgCBgChoAhYAgYAoaAIbDXImCExV479TZwQ8AQMAR2PgLFS5Upv2zJ4kXz5syeufOt2XUtKFWuYuWlixctnD93zqxdwcpylU+pMXvGtCmrV+1eqZWIDAC/MSNt5//WrqNkMKTM+vR16yZNGGdaIakBvdwVZyc+DnMc+HLYZwd598sTrP/XRSBkOZ2E9WlBZqYc7PRAqiGc4SIoRCqEtSCIYMB5LqFrfaYNnvlEQjzLVQaSgX6wEVtFlOCYVyQHbeC0D5MKilqgDVJM0TdkC9EVpFEKEx6046eX0jj9FE0QCSJaNG5FgVA/npYGz9Se+qUvjUGC4JoLbOazRModWZGZN1g1rGAw9QX6PyAKnI+lRLqZW+bYDkPAEDAEDAFDwBAwBAwBQ8AQSICAERa2PAwBQ8AQMAR2GgJEDowbNXzITjNgN+m4VNkKlcePHrFLRKGgOVL45GIldsd5q1Cl+qmZGRkZE8aMGr6bTP0uZ2YyGFaoUu1UMAbrXW4Au7BBbuc9Dvhl7gwLb+cJVo/JDtZN3RisGp4VZK5yLvYIYSEnPPUgHxRhwSjDaZk0csgNHOeUl9C2L15NW2HNiTBqioyQDdLCoE9sp20ORUUoEkPt8B0ywY/MkM6DNDr8v1F8bQm1ATlAGz5JIVKBe9KXSGbGfRylWUFbDugIjqSB8kkSpYeizDqXqmtDMPYa3fOFw8OC28uic5yMTVbGEDAEDAFDwBAwBAwBQ8AQ2GsRMMJir516G7ghYAgYAjsXgSOOOuZYRJvHjRpmhEWCqTj6uONPPPjQww7fVdJmlS5fqUoed4wdOXSX0NNIZRUTGcKuf3b/p1LPyv6HQG4Yol2BhoVFsWzdqnEObaIMRCb4ehR5g2X98wZ5CmQHGUud+3xlniAj3ReTxqkuPQcc9n5qKIgDEQG0yY5/HPq6D3GhVEi5kRVhnQoG6kc6YL8iLrBBQtjhvznox48ikdZEjsj4f4cEvP0rqbMUUaEoDz+tlUS5k5kEER6yM5wayo+U8MeSk/Zp3ezMYEbTzCB9nrRFsF/9gwt1wHdddG6TscnKGAKGgCFgCBgChoAhYAgYAns1AkZY7NXTb4M3BAwBQ2DnIVCmQqWq9L477tTfkaiVKV85gtOuEmFRulzFKtizqwiAJzsXBQrss0+pchUqm65CsohtWS4ZDMtWrFotLW/evKYTsvU449x2pxzyEuDOE+xzlHPlF3LpoFZlBxsXZAVZq6SroFRGEnemc5zlipYQgcGVMpxKxyRxapEfSteUiLjwUzZJF8MXrPYjKrDRT8ekqAvu4czXMyIsdOqebOCqFE1gg+2cSsvEeP0+Uvn7RmWlnaFICnA/zJ2QKsJZURvYjYD2SieGXjCY185PKSXyRnOheTSSdJteCatsCBgChoAhYAgYAoaAIbA3IZDKP+j3JlxsrIaAIWAIGAL/zwiUqVD5FLowwiIx0KWjxM7YkbtG6qySTk8jI2Pjxn/Gjh7x/7xEtmvzpcpXrJI/f4ECY0xwe6txTQbD8i4dFB2MGWGC21sLtNuJj3Mbhzi79TlxkK8OVgxMDzYscp/TMoPMjDyBi3QKNqzIE2RlSdyZcr4jXwSAIi8wSVEVK6Ofccgr0oE+aUORHT5hEGs4tM+hiALID+lV0IaiOhQdQVn/bw9FUkgY2ycdfBKAetKOUFlfkDtMrsQiWxQ54Wt/0K6+g4EIHq6kzhJRQTnGxnjAyNXKyhNMb3JQMPZGoicox1XC50SAMH7N39ronMbC0O4ZAoaAIWAIGAKGgCFgCBgChkAIASMsbEkYAoaAIWAI7BQEylSocgpi24hJ7xQDdpNO2bG+YN7cOUsWLZi/K5hMlMJkl1Zpw/p05b/fFczK1QZ0FSg0dsSw3S6VVa6Di1HguBMKFznZqdpvTd14dZLBkDJLFi9cwLsdq528+fLlO/fiK64++tjjT9ietu1pbTkHN4QCjm9pIhQI1ox3BMVC50x3vvDsDXmD9fMygyxXLHOdi7rIwGnui1/L+e4LcYsg4N//pJDyNSYgABDuVrooP61SPMFqP5KCVFCyVZEPkAwc4RRN4fZitS/iIyzADQnA4dcJi4vHak8po/zUUf6yIaICvCEmGIvIB+HIGHJ+8zKWZQcrh+QJZr+rNFAIh6tP7FYkBnisjs7lnrZEbTyGgCFgCBgChoAhYAgYAobA/xsCRlj8v0FrDRsChoAhsHsiUN7l+f+h77B/7m7wxLPhEVxw+dXXterUrc/2cISWq1S1uu3Czn2NlClfqequkn7pgAMPOrhIsZKlXVTMLiEAnjt6/5VAe2HN6lUrZ0yd9E8q9XbXss0+/Pzrb38fPLZJ849aF9hnXxzR23wkgyFlEpFCL739SZt3Wrf/4bEXmr2zzQbt4Q04Rzdk7nKc3u7EkZ4nWP57WrB+kXOeOz96VqaLrlidHWS7x1nr8wSZkaxOiraQNoNQEmmAk12RFzj/IShwuONk1zqR/kVuCPskAPUhQTg51EYyehLxIiJoxydFRL740RWyMR6pkmgM0pgAKz7TLpgcFMWIMWkcEBoFgsz0PMGKv9KCKU9lBhtXSfibvoWlhMeZs+XROcwNR3tuCBgChoAhYAgYAoaAIWAIGAIeAkZY2HIwBAwBQ8AQ2AyBex556vmTihYvWa/B48/4DxDSfaNF246nnFbznBJlylXcFthOOOnkYghJW577xCiyS/6gQw49bFdJm1WhavXT0tyxq+hppLIGy1U6pfq4kcOGZLsjlXq7a9kXGtW/A6Lr6pvq1vv4q+96oCuxrWPJDUME4g87/MijHM5xo1gOPfyII7Fj+l5CHG0r5q4+kRbSbMgMFvdMDxZ9u9FFWjiiYo37d7wT4V47NU+Qvcy53FfiQIeMkFaFIg/8Ne+LVCvlEc8V0YDJOO/1N4KiMDSU8Pvj98EzXyicNsIpmGJB4rep8opsUHlFWsjWeO9xovRQ4WfqQ2mwJJhNn9LmUDqrHCJi3eSMYP7/HHH0B2VhiJgbtQupRHnNF3NnhyFgCBgChoAhYAgYAoaAIWAIpIiAERYpAmbFDQFDwBDY0xFgFzpj7Njus4/9se67334FXcr0PPPnzpnV//ee3bYFB6I4qD9m5NDB29LOnl63bKWq1RjjrkJYVK522pnY88/YUbuVfgWkD+TPrhKpsiPW7cxpUybdcc2FZ3zzxacfQDLeXv+RJ7al32QwJH0ZfYwdOTQuYfHYPXVqX3NO1VItmjd9flvs2Vvquh36OMUXuVNkRFqweqRLBzU3OyhwRHaQ6TQs8hXMCtYvJU3UvsHGJdr170cPKIKAKAGfgPAFsH1I/b8Pwn8rxItkgCjJ0Xf4Lz2SojzCdWKRHurfT60k8oN2wIHvStXk62L4tidKNxV+xthkIwSEH8EhQXCeg9uaIH1G3mDqc/mC+d9QjntEp3DlUDSGCKNF0bnbW5aqjdMQMAQMAUPAEDAEDAFDwBDYbggYYbHdoLSGDAFDwBDYMxD47L03Xnn24btvfe/V55/0R4TT/MaLz6h082U1q4rU2NoRs1M/MyMjY8KYUcO3to29oV7ZilWqEREwfhdJwVS5+mlnZmVmZk6dOGHs7oQ/OGLv3kRYMF7m6q2XGzea/M+4MXXuqv/wtkRZJIOh1msigm3d2rVrZkydPHF3Wj8721bn+EZTYYk7EePOCFZPcOmIljodhZHMsouuyEgLstdmB+mznHN9Y4EgY13eIGODBK8xX9ETvnB1LNFqRUT4+hfJDJ96EtkmyoD6vpB2IoIiVvtKAyVCYZUrpMgL7CYyhDMWeZKMAHfk9XAntqo87cpu3UOzYq1LA5UdrBqeN1jWNztY3IVxSqdCuh+yl2fM0ZLonCWDnZUxBAwBQ8AQMAQMAUPAEDAEDIEQAkZY2JIwBAwBQ2APR6DQ/gccmMoQp0+ZOKH7D52+jlVn8oSxo5cvXbI4t/YKFNhnH6Ix4pWrUKXGaZOccPP69HU4d/baIzec0AOY6Zy7Luhlxc4GKX/+AgVwSM+aMW3Khg3rtat4u5lFijCILNIKbbdGow2VdQLvfBwzYu+L6IG06NSu1ceHH3n0MWUrVI7gEO/Ily8/u8NjHslgSPuzpk+dvHLFcpefaMuDdFAnFStRanvPr9pLZP//V587ql3nAOc3AMd9ZpC9cUOwfOC6YJ9j04N1szOcQz0ryHuoSxHlNC3WTssOstZkBxlO5yJHiJtDaZtwwPuaEDjcFS0AwcFzEQ25DU1OfT+FExEH0seQvoWiFuK15z9XW9RVVAW/NRABKqf/rviC4bHajhc9orK07wtkq31FpnBNDzJW5QnW/ZMWLP09CMbfqegVcMImbHOhLZGr0kGtis5VbvjZc0PAEDAEDAFDwBAwBAwBQ8AQiIOAERa2NAwBQ8AQ2AEI7OPyKb33RYef2v3Ya2DLb7r0avH1jz0//ur7Hh+07dz1vS86dnn3829+fLvV19+jEVH11DPP9k2qdvpZ5z772nufJjKzYKFC+8ciCK647ua6fUZPXyTS4qCDDzn0qZebf/BNj/7D6RcBZbV76z0PNrzutnr1E/VTaP/9D0j0HFFuhH4HT12U3mv4lPkVT6lxerj8fgULFnJyGBXGjx4+lDQ1PQaPn/Xr0Ilz69738OM7YCridlGsZJlyr7zbsl3rzt37Mo54BXcUTuyGL12uUhXfyQ5pcEPdex54+Z1P2950x70PJSKFtgVLyIMHHn/25c+/+6Vfp9/+Gv3AE8+9UrZSlWqs4ylut34ybeM8vtnt6m/Z4effm7732ZeJiLM7H2z0dK9hk+fxfvQYNH7mW5/97ztSkCXTTzJlsH3BvLlzFi+cPy+Z8pRJdj0wT0+98taHZ11wyRV+2+dfemVtxgEGyfQJWfN+m04/9x09Y3HvkdMWvv7xF99cf9vd91P3iKOOOfbVD1r/z2meHxKrLd7jNt//OiDe81FDBw+k3tHHnRCTDDrvklrXMM9Dpi/Z8F3vv8fFIo1yw5C1WKZilVMSRbG88OZHrdt817N/3nz55EiPCU0iLMIVwJ/1w28IvzsIevOeJIP57lbGOcIR4IYM2hAscVn5Vo8s4OiFvEGWE4Je3seJbjtNi+z17rsT4E6f5a6rHJmxEUe8oi0gE/gsIWk+c/qi2z4BAUQ47imj1EkiPPxycvyTVsmPfBBpEdaj8KH3iW0/UkFkCnWZT/rnhOTWZ64iYyinCAnaj/c3jggJniuiRGXVLmTEmiBj9cZg/fQ0lwIqTzDlSQgJxidxccbJ54Pdia08Xxado91taZm9hoAhYAgYAoaAIWAIGAKGwC6FgBEWu9R0mDGGgCGwJyPgMiBl7OeIhf2c13/jhg0bVq1aEdk1v/8BBxx41DHHHY/DEydn2Al9x/2PPnlMHEcj9UuVq1j516GT5p553kWXhfFjV3Re5x3MctusEbru0PPPkTc6R/e+jjWgv7MvvLQWdXAu12/07EuOj4gbjXHNzbff3X/83BWQI7HmqX6jxi82//TLzmvXrFn9VauP3nFBFvs89nyzt7ewyeW5x2GJk/Tya2+6rWejptYuAAAgAElEQVSX7zpQ59FnX3kTnYGdsQYgatr36DcMggfCqHHTtzfT75BNOxKnosVLlYHcEWFx2BFHHf1ll98HNX717Y+xEyc5AunbG6/yVaqd2tk5r2+6s34D9ErWubm55+Enn3vu9fdb0tf4MSOH5dYnu/m/+L5n/ydfevP96mecfR7zfHntm26NVa90+YpVGjzVpBkRNy3eevUF9DF4D+rUe+CR3PpJ9jmRIamkg0p2PdA/eiyQR7wfsgdSCbKCcYDBhVdcc30iWymPI/+4EwsX+fyjt19Dd+KsCy6rVafe/REMylWqWv2ya264JV4751x02ZWVqp16RqnylarE6scF6ODoDmKRRvy+QJYyzx3atPzw+MJFit7XsHGTLd/bxBieWKRocffzcVAi/YpFC+b9CxmW6HcmNyx8u3gf33G2s35G/P3XgN+6/dD53IuvuPqiK2vfmOza2N3KOYf4amczOkPLg4kN0oP0ORsdQZEV7Ot+OtOcAPfGpVnBhlmOxtgvT7B+ZprTtFAkBI56IgH4tz8RAhw4+yExSDlFu3LY+8SBCIVwqidf70HRCiIBBKuvl6E2pT0RjvbwIy2UCor6EAPY6JML1BWJoj58AiJWWij/nsgNiAbaVt/09R85s2JAgWDmW2nBzDcZe6EoPr6uhlJK8X6tjM7N7rakzF5DwBAwBAwBQ8AQMAQMAUPAEDAEDAFDwBAwBLZE4OJa1944YvbK7HCUAQ65gRPnr463SzvNHeyMHjZzeebRxx5/Qrjljo6gYNc6kRXd/xo3o8+o6YtwIFMOEV2RI0RC0H/x0uUqxJqfY44/ofCgyQvWduk/cnKs57Wur3M79Z9p9k4LtQmBwT0Ef/06dzd44lnuE02inPo4Y7l38ZXX3bSj1we7s+n75z9HT4X0uahW7Rv4zo728C7/HYnTtbfceS924NAnsqVzr0Fj+o6ZuaTm+Rdfzvdf/p4w+/cRUxdsT7wgv1hv7bv3G3rIYYcfQdvMJ9FA2BJrPsP9Q76xTigLqcK6JKLn+95DxseaXxz6lCWKgLYgaVgb4YiFrR3nkUcfexzt3/lAw6eSaSOV9UB7RNzQ/m33NniM75AjQ6cv3chO/0uvvr7O8FkrslhL8fqG1KBM0/dbfaXIgAL77Lvv4CkL14kk4v3T+xWrHaJYeH557RtjkkJFXUgTz1nbfv1zLrr8Ku4TWcRvCc8gWjr9OnCUXy4ZDPUOQ+DEGyvRXb1GTJm/LVj4dR9v8vq72C+yiLVKhAprKpm53l3LZPcK8rrzCHce484i2f9+USp74Y/lsxf/XDZ7xcAK2ct6V8peNaxC9qKuFbJXjS6fvX5FBSeFU9qdZdxZ3p0nuLNi9DP3+EyZ4u4sFv1eNnqtFK2nupXd9yrRU5/9K+V1Uo7PtF8u2jb9l4ze47nfnr7LHsrSL+VPcmcJd5ZyZ9Holbrh+rIt3pU2NXau2MfY6QeMirizcPbcNidk9zvmRIdvCXee7M6y7izqzpPcWcydPCsSnQPmwtcE2V2XltltCBgChoAhYAgYAoaAIWAI7BIIWITFLjENZoQhYAjszQic7HbSN3nr488H9u31y1effbhZREKZipVPieyyHz5kUCyMLrnqupuLlypb/q8/fu85/985s/0yOJwhIAa6Zzg+Czon993XX3bO33/+0ZtyK5YtXeIcM5Fdp0QVEOUwdeL4mGLK7LAnHdD37du2CttB+pjGTd/5eOSQQX++/vwTDdRm5y8//+QLt1ucHfN+nco1Tq/Jju9Xnnr4XvLr84y2uWY6Je4duRbA7+GnX3yNKIZbLz+72oDev3Z36ffJSR7gbCYSxbdnR+JEpAMaH0QePPva+58ef2KRk++vc9VF/X/v2W3N6tWrJrv7aALg3N4emNEORAH6FI/ceeOVy5YsXkS7zGeXTl+3jcyPixJKtIMegselPuty3Iknnfx8w/tuf+P5xxuwLt0w1hYpXrJ0pRgpwo51UTW0y+57+kCU+akH7rixX69fum6PcZWJ6jYkEoJWP6muB+qVcmm7uPbp2fVHCLjn3/jgM+bsqfvvuLHHj53bz5s7e6YLjomQMeGD+ePdHD74z34vNKp/x0YXekWZKtVPq8l8/PFb9y58nzdn9kyE7v0UbmrLBTUcXMW9U3wX6RPup/DJxUpwz/+NoB62Thw3euTLTza4J8sdlHFTWDAjI3Oz9zAZDMu4aK6MjI0b3U/IZmSHb0vp8pWqjhs5fMi2YKG6kIdEoHT6slWLH75p15r7rFXWoDN/h/6ObI91mkobbic/v5uR3yl3ZAXj71kTrJ+bGaxFdDvb6Vkc4vQsNqYFBY50T11KqA1z04INC/YJsjKIlmCeSe0nzQWiFdDGkE4OUQZr3akoB/4bQeoj6inKgXtgrOgL/6pIB6Vq4qqUVER4kNIqt/mRnbRFBAT/fSCyT4LbaGXwWSmnwvCFIywiyyNaiPFpLNySVkZO6qssJ2D+72cFg0mP7hNsmCdhbmwAp8j7Ga3va4Esjc5J2A77bggYAoaAIWAIGAKGgCFgCBgCW4GAERZbAZpVMQQMAUNgeyFAeqW3Wn717ZrVK1c+9+i9deXsV/sVq9Y4Hac+DtBwnzhHlRLou6/bfBZ+XqXGGWex49hlZtoXTYZnH7771qmuoVi208+k8WNGyWnplyFNExEUOCO7dP66bbh+w2ebNne+1f3eeOGJBiIgKLNk8cIFH77x0jO+YDS7uCu6XP3df+j4tX+/Rs1zLqDv0cP+/mt7YZtbOzhPX3RE0RTnYX3w1msuEVFR69qb61J3/OgRQ8MC4zsKJ/pnpzrpl2qed/HlkCevPdvowQleOqb8bjs+Du4N69OV3iW3ISd8Tmog0vq0/uDNpiIPVEHpy8AE8iFeQy+9/UkbojSaPv3IfV2//eZLytEmmgR8/rPvb7+E6650BBEpwuI527dpUK4y2gu8V872hKmstmY9YFupchUqz5w2ZdKcmdOn1nZpodC+aOKRD25ocYWsST0GKfbi4w/W89+d08+98BK+Q2Ro/DOc+HqRGILVZ7t0UBKbjoch5BcYTJ88cYLaQz8GwuTVxo/WF1HCPBQrVab85H/GbvZ7kwyGRJZMnjB+TLz1iI1EC8UjX1PBgjE8+swrb0Kqvd/shU2RMwh6Q35OnrC5/du6hnbF+lEHORFWjgzIzAqmPrs+WD9tY7Bh0UaXBsoxf87Znu+gNEdkZAXp/7j7CzcG6dOcy301Tn4/FRKEJ8QsKY90SOOCq4gHyvFZAtjhvyGkaaE2RCZwpS59QpTQD/2FNSfC9USOcF86FtImkbB3vKnxdTH8dvks3QsRFbqucxilBQu/yQ4m3Lc8yFzBOH2c+KyyIlQgYhZsT7KCPQTuzBM99TnNfdepZ3zX53hX6kfa2BXXsNlkCBgChoAhYAgYAoaAIWAIxEPACAtbG4aAIWAI7EQEnn/jw8/Y/dz4oXp1tKPdNwfnPs7QWE5A0r+cVLR4SRz/7LoPDwOHN05P9A5wHv/Z57ce8YZawTk0w05Klb234dMv4Gwc3L9vr6WLFy302yDVDHn1u373zZfhSIpYfZUoU74iefR9e0+tee6FpMSCDFk4/9+5O2I6ECdG6Bx3/8N3XH+Fcvwf7yID2GWPDX8P6Pt72JYdhRNaAOymnzh29IgnXnrjvT9+6/FzmCw6rnCRk2dNnxozRVeqGJJi6rZ7H2r075xZMzq2bbWFfgcpgWhz6KABf8Rrm3RmpBz6X6uP39WOd8re9dBjjSGqiKIYFqP+4AF9elGOVFep2p1MeXb+g5NPkIXrbe16IAqiSNESpYYM7NengBNtqdfg8Wc7tP3so8lRYXJSPB3uwiuIZgr3WbJshUoQiZ+9/8YrkB3+8zPOueCSSc7pTiSN7s+ZOW0qOiZh4ftLXBo11Y8llk192kMsXescp/4Nt9/zAO+hL+p+5fW33MFci2xS37lhCHkKUTV+9PCh8eYEYge8Rg/fkpRMFQsIMDQ72n36fnMiw9QnkWBEovTt2e2nZNbGjizjOaJ9x/M2meAc5VnuJDJpVZCxPD2Y+fbGYJEb+oYFjqw4IE+QgTSF81hnumiL9bPSgoxl+YLMf/MFGxenES7lHurvAOky+ILauicbcdZL1BoHuC/CLQ2IsGPc162gHfojwkHXWOP324Ik8Mvqs+4ni59PpijiQwLe6UHm6jUuqiJfMOGutGBcXfqAVMFOX5uDvkS8RKJSwJ45SNaIROU8YgH7sIExKs2UvmOTTj33ywljzesmTZEoucHay+udEB1hIiRMfkRIDzsMAUPAEDAEDAFDwBAwBAyBHYmAERY7Em3ryxAwBAwBDwHEZXGOf/J2syZD/+rfNxY4OArl/PSf54g/P/Mi9wb16/0b0Q/h+pADOBLRr/jozZefjQf+sc5LjxAuu6PDZSBErqh9023cj0WKIDZMFIcT6/0omcl1TsYzKaf0PJWrnXbmW599/R1O0+ZNntxuIsu52fLQUy+8itYCaalIt6Py9zz61PPsMuf76FAarh2JU9lKVauBa0nn5D30sCOOfP35xx7yx0RkDpEvkxKk38kNA/95LeeohiQh5Zd22/vPcTbzPRbhwH2weeDxZ1+GtPrgtSZPqy4Czlo/RLKQ7ils1+89unyPI/26W++6LxWbky1b1qWEIjIkUfmtWQ+05zilcrxjOOGvvOGWOxwZd8Bn773+sj9+ns+eMW1KuH90aXC2d/6y9Sf+M/QqSBPnUqwN8O/PjpIaRKzoPmnfIPwgiYgQOsapdof7gfgiNRzpzvTs3Isvv5qUUB3afPqh7p3uSI2nm7710c+d27eDgPHbyQ1DBOJJxZQIZ0gGCNRYKcVSxQJiBRLXJ8YQCkdHo3mTpx4VMZPsGvn/Kufvlnd9KJ2Rn8po0076bbHBOc0R4V7nzszg3zbpwerRLj3UJCe+/e/6YL+T8gX7FcnryIvsIE8+lx5qeVaQsSozyJyfP8hM953emKCoBhzypG/ivyu0y2df3JrPEs2WiHbYce8TD3wmnZIc6NQV+eEPXXVo08dJhIOc+cnCRT3fPj5DxGALZ0aw9h+HWauDgklPrgkWd2O8ImpEihBRpv4lSr4uinmydsQtFyIqNB8aJ5EkPg58Jx0W/43SehKBQfSJCB1FoChChvYoRxmfBFJ/IpH8qJjNPnsRH0ZgbPOsWwOGgCFgCBgChoAhYAgYArkhYIRFbgjZc0PAEDAE/h8QIP3MY02avYO+xOcfvdUsVhc4pdkxPWXihC10Ja668dY7cRJTb9SwwQNj1Xc+xPLc/9lFVyyYN3dOvGEULVm6LM9i6VfgBJQwdrgfdo9fcvX1N5OmyE9VlAiuKtVPr0mqKHac46Rs2fHn3yFr7q9z5YX+Tun/B8g3NQn2195yVyRl0W9df+isB6TywbmulEfO+T7ct2NH4lTeiT3Qd0UnZoAOyPy5c2b5thRzuiUQGqTx2h5YnXdJrWtIGdTt+w4xxaEhlnA2jxzy12ZOdPX95Mtvvs86adygXh2f8GjwVJPI2ubehBCeqgveHdq2/Ih5qVHz3Au2x3jUBu8I4vKJdv5v7XqgDyIDuE4YPXLYLXc/2LDtJ++96bgXcvRHDq2Zae4l9seFTZc6srJLp/+1CUd+nHHuRZdSduTQzd/rubNmTuf+8YVPLqq2Lq5V+8ZMNzE9fuzUnigSp2++BWFxTZ3b76Z8t+87bprb084+/yLew0ED+vaCuGj0QrO3P2z3bbchf/brjZ6Fb2uyGFInN8KCqJHwe741WGA/GicQEyecdHIxROHrN2r8YovmTZ//yWG6PdfQdmjLjyrYtOPdtatd8/F0GFLtGk0LCMH1wcw31garhmYEG50sxZoJGcHyPzOCDS6qImNZnmCD0zzf4ALlNqzME6yfnR1sXJ3mZC98RzdObKVtwpGNg1wpoiAupD/BfQ4986MzRF74JAc6FHxXmiU+q44+056iGkQSiMQQHqls9/cjQqhPXSJyNrgxrwsW/ZAWjL8rTzCpkSNwVsiZTxSFNDsoz/iUCorxg7H0Q1Kdo3jl/agKyvBd5AS4iXgBe2l66DnptbBXJAWfpdMh/RHGxD2utKc5UMQIY6R+hKyP9ucTbJuRbJECOemolHJqe+Fg7RgChoAhYAgYAoaAIWAIGAIRBIywsIVgCBgChsAORgAHYfOWX3UmBRS6EmHdCpnDLmuc0jOnTZ7om0h0BWl2lAYmHAlAWaIqDj/y6GP43NGlqEk0RNI68XxGqB/ywbsUPzfSD05lnI1+O9XOOOs8duX/+vP3nZKFsHL1085cumjhgladuvV59JmX3/jwtRcbN6x301V+6ptk29qacuD5TLN3Wzhd6fT3vUgA2nqsyWvv4Fgf1L/3bziRwyLmOxKnci6dFzYtdELUX4aE2Llfwu2Y57o9CAt2xjMvY12US5gYoY/DDj/yKHboh1MUCf8zz7vosrMvvOxKUknNmDLpH90nZQ8ponp1//FbyC1SEsWbs69afvg2qXzueqDhpuiMrZnfcB1HRkQEsSeM2Zx8UrltWQ+aB4TRiSThnfMjFnjOO5wzT5sLUUMQkR7p+6hYtG83miV8HzVs0GZEpN53HPQqf8V1deoi9g1JMtNpXOD8J+Wanjt5jEJX33jbXURM+Po16NuMHTHsb1Io9Rg8fubNd97XoOW7r7/08J031ApHa+WGIX1Rhndnyj/jtyBXZUuFytVPdSTMn+E5ShWLox0rA4lCqrxX3m3Z7se+w/5BFLzR3XWuaeX0V7bHutmaNnznrbQFXDthIoCmteudz3IEb3IAb03f1HE7/jm8SIsv1gYT6qYHa8ZmBAdWyQ72L5URpBV0ERaLnRM7My3YOC/bRRdkBSv6bHRlshxx4W5vFFngEw6KUMARjoMbx3Y4xZIiM6RvoWHovsYsxz+kQY7I9X9i2NRRminpW6g93Y8MNQ5GPukhB79SV9EO54pg/Zy1weKfMoN+h+YJRtd24/9LpISc9diEfUSBiEjgnlJIrYxivbVTFa6nPhQ1IeIAYgFSCEKCk8/S8BA+inzhOaLkIh6oywnxdLA7D49+57kiNGiDPkUAKVJDBBp2iMQRwSHs/cgN08fYXivB2jEEDAFDwBAwBAwBQ8AQ2ISA/nFukBgChoAhYAjsIARefvfTtkcfc9wJ9a6/9OywqLNvwnEnnFSE72Gdgqtvuu2ug10umJ+//bpd7Tp33PNPDGcsO/CpS+RDrJRSm/dTuAjO4rA+Rf2GTzfJEVleuxZtCV8UmPo1zjznfK7SIMgNPpy6kCicpAa67oJTy8dKlZNbO9vyHJ2EcpWqVm/9YfNXFy+cP09tnXvxFVeTWof7p9Y870JfnFhlSMG0I3CiP/RHuH7y1qsv4BAPj7lEmXIVueeyLG1zhAVOdUiwYZ7As9/f+ZdddS2O/VjOZso98PhzL0PwgJ3qEW3x5Etvvh/RV3GpiC52OguxMFV5dsp3ateqxZ0PNnoacmR7iSaXLFu+EoRgPH2VbVkP2M48OJ5vPKnRvmr10Tvh6AEnb1EWR3547Gece+Gl6IWExwnhcPo551/M+xYmj+bMmu4Uk/+PvfOAk6JY/vhe4MgYyElyhiNHQVDMiPoMPEygfx/mhCgGEDMmRDEgGEBAEBFUEAQREQVBcs4555y59K/vsoXDsHt3e3d7XKh5rz+7O9Pd0/3t3sWr31SVx6OCBetGouu+vd7owfl1q1cs45WQUerxRNg5BFK8dJQ1eTDI1UJpLuOYMGbU8H7vv/myDMfbv/tIiqGXg3Bes2L5En+h6bjOd55QVxLm6hzBIlgWtRs0uZQ+JV/Ii+wvPNQG9fuoF99Nf+M/j+f8hddRQy8GYAzGfMYofCaHhGzXePm6pWjY5FNImOQVLeg7rydBhIn1b8R5jq9P8FzQMpcn/qCEhRLNIWb/Kc/JHVGeqGJhnuMrEzzhOeM98SfCPRH5wz3hueIlhJSOB4M4hm9NMu18ZYzOMFDqMYJh32kId05GvQWYM/UIt+Ssr4muNXeDhi/yFz7KzYj7IyzQJ8Z7FTBUcDnsWXD9Sc/e8U7BSD0p6AuBgqTgjF3zXGDMV1EAz4ojwjgYD49E19GXG8LpaaPCjObPYEwIDBq6iTBWfHaKSOq1w3n4MXaECooz1wfj598SFSyop94zui70r3Nn7DpX+uG99ufMZ+KdoyPPhbdNSvdwosDsohEwAkbACBgBI2AEjEC2IWAeFtlmqW2iRsAIZAQCJCZudXWbmz56+5UXFrpCvrjHJzY+b6Lj7Vs3nwkHxFPZnZ7s+hJPcvOk8cqlixdI3mgMKmcdGBk58euYUd8lNe/CkmTXeQ/qYzS+WhJhfybGUMLe+PPiwFiKwXCFJIZO6h5cJxwUrxhvefJbQtCfY4hPTj+pqXPPA493wVtksBg4tR/yd3R7+8N+GGwHfdbnPUJpbZWEAe77pBcnDLsXFypchCfqx/4wfIi/+VaSpBIILnt375T4Lqk7yoknDT0ECvd0y50dvSGC/IVVqt+keUtCKiE2OBNL3/9olxc4/5F40LBPae+PqXPkwwb0+whRDI+A1M3o39aVq0fX4b6BjNmp2Q/cBWFQtJ6oatF1hcHn5yQrJyTU2pXLl7rzgtSWfA5zZ5ybwJwE2jBY7Mqfwr12bd+2hX5EN/OGhGp7+50d2QP/TP3jNz7/K1hU9Oa4IKQcvzeIF1qH80WLlyjF67hRw4fc0Dy6QvcnO90TSKygXlIMvblWJF/OymWLFgRat9oNGjfj2sI55woWwbLQ8fd+vdsz1zSsUqqviHoZSKxwixQYzTXvgXoXYFRXzwoNr6Qhfc54XKT0O4BBXQrJ2vdIOT2eHUNjPBtePuGJORAjOS1ElMgd6YnMF+aJyBnuyVlawkTtyeE5OEuSce/P4YnZF+7Z+X2U5+gyScx9IpcvXBRhzpxGajWS6zlneCcVY1SocKsvTkZqfMeYTl881e/0ylBBRIUSNxb1pNCcGvxbSJ+INoc98XGHJKH2cc/hBXGeNV3yiFiBEIAocYEUDPoaoko9E3jFaK+Geh3rHpimpVjhm4iyUaFC584Y8PJQAUc9JtRjhFfOFfTNRcNCcY6DduwB1g3Rg8/MHU8LPC4u9rWFFTz4fJGv8B7vTGXEdby2uBdt8bJhnNxLPW40DJUKGmdys1jCbt+K2IsRMAJGwAgYASNgBIxAUARMsAgKl1U2AkbACKScAEa7J55/5S1irw9xhfkhrI4z1At3ubhwkaJxsbGxTkPw3Z0e7UxiX8IEVRFjbCAPhao1anuTJE+e8POPSY1YcjoX3bvrbMN35+5vvIeggncHT2j7uw9Pcm/fsmljoJBW7vuq0ZLQM8yrza2nk3mn14EQgIF94tgfRjiT8nZ/u09/wvm88Oh9d0j0o2I5JUbSts0bN7jHlV6catVt6PWuIAG226tFx1SpWo1agcIcBcsTwYY2Wzae+4Q9OSU0T4O/BN8YzWk7aujAz/W+CBUPdH6ux5SJ40Z/P+TLzxCA2CPO5Ob+xqjG98uuvPaGYOcQqD6G9EChqFK7H4qI0CdfjYsqiWgxcshX/dxhzfBaKVO+YmV3LhS8KPA4cHtXhMtxxbU3/CdOklL4Ewjj5diyYf1avnd4sLS55b93jxXRQfcIwggcylaoVIXXjg89+SzC1yfvvtbdyUe2OoZHz/jR33/rLwSYm2ViDKlLeCbCUCUW8gtRghBr7jBrKWGh4x8x+Mu+6ZX3Jsj96Azxo4ZczQWhxnwN6aMGeX2C3RueKC2MvGJcx0gtySq8xvs4z8ntsZ4Nb57wrHv+hOfgX7Ge2INxnhPr40TOiBSjfpwnX804T+yBBEnIncMTVTiHZ/coETGm5vAcl5/Ck9swXmNE53B6VagnhCJy55two9OcFXpevQswfHONMasYoteoq2GbnMKIMywV86QgWJw+f3JbTplnpGfD21GeXcNyerZ7U7ho2CQEEu7FfelT7+sMQYWIALtdPpZBboOgqrNnnN4QmsMCUUW94VXMQuh3ckcA0yTinEdUQMBgzTR3BYNBdOAaBbGBOrzSP/OmHz6roKOhqOiDc4xFw1Kp0ME5FXucCb11fF7BJy32c1A0rbIRMAJGwAgYASNgBIxApidggkWmX0KbgBEwApmBAEbhd/p+/d1ueSK6R+cHOzqN/Bgq3//8m1FvfzrwW+dceEJaIifxlKX3wMj5f/Lk+pcfvffmKXFPICF3oGTa8gB+XUSG5IRcct+HMDmER+r9RrdnylWqUo17+7uPRKUqLOkozoRVSmodECx4QnzKb7+MIQzNPZ0ee9oZbz+p9qm93vzya67nafA/Joz9Sfvq9ORzL7W+7sZbPnnntW5LFsydhTGYaxKRZ7P7funFiZBV3JvcBP7mrAbitAqblCdvfoxRnj0ub42IyMjILi+9+T7X2G9qEHeOCaFt5dJFCwhvxHnCDX3w1bc/ST7nHa90ecTrKXFJuYqVyNfizxPIPT9CBhE6DNEoteutSev9jZu+U7sfKvqS2hMG6duB/T92j5e9hGixRuJ2Oa9pYuydYr13nr9JPEti5AuC9xH5RPzNf/3aVSsKi4sBeR94dSaYxpMEA37FKtVqFi1estQ9DzzRhT00fcqkCc6+CojFn8/yVTzHM8vfnud3JhBD6pevfDpPR2J1atdv3Gzh3LOTiNMmJSz+Hf+5nmWp3TOpbK9P46vRXoULuuU9Bl19Kl3fawJkfaLf2TaVw/HmtcAIjdF9r5TTgsPhpXGerV8e8uz6Mc5z4J94z7HVCBVhnth9kZ6Tm8I9x5cmeOKOh3ny1iI8VLgn/likJO4O9xxdId4Xh8MkzwVzUS8EDU3kFDFUXHCPX+fm9KDQnAqaq0GFG/UkUDHB7WHBZxUsJLO4zwAfF5PbE7M7zHNoVk7PyQ3hIlrgMeLxbP7ilCQa514qHEmPgQUAACAASURBVKkQwPhVCMATQdeB+cGMfBUwDNXhZMJY1OMGTxOniKP5LVRg0fwfjIu5UP90GLDTogL1ECgQaHhP0WvcUxNwq4ihggT1aAMTFSrYqyqA8EqbYlLwyOC+HLqvde1VKNG/M894XIQKpPVrBIyAETACRsAIGAEjkLUImGCRtdbTZmMEjEAGJIAg8dYnA4YVEmPu84/e117y44oF5d+DJ6d/G/vT9ySOxZtBrxD+yZm/4Pk3en2yTyzBQ7/s+6Hmt/AnJJDgGKGBRLvJwXH6PqfDM+XNly//82+8/8kvP3z3DWFpyNvAecLR+OuLhM3u84gzmqBaryFMlBNLKqIAcyLUFEbpl97p099fvxWrVK+ZnLEHU6d67boNqL/YZwy+7ubb73y4y4uv/j5+zA+D+58OEVVUHrvn9cjhgxjBzjrSgxM3rCGCBU++b5Akyv7mR7guzrsN4cGwcNZFjOCzLOVZa3nX/Y88Rcgj1kuiZa1x5ycg1BMJuZUna9xn4HdjcCDo+lCH23Wfi/G8NKHD3OND3MADwXk+TL4rfB8CeZYEM8ciYrSn/sb1a1b5a5fa/aB7FAHMmQ9F70U4KN6vW3U6t4QeKhCJznHGEMr3ngTYiD9wXiq5Y6iPJ4WzrYZ9wlNr/uwZ05xJzhFBSazNuLr06Nk7PDwsvNcrz3d2z100UELFeORrn6QolBRD+inqC/kViDO/R1Vr1a63aO6sGe6xpIRFMOMPZr+kpK4v0bbXGMtySdFcAxhyNXmyhv3RvBAqbFBX8yVgrNbzDCXNnkoXg3ucFH7fd0rheyjeFltzeA7POubZPynOs33wMc+WfrGejb1jPPGSdPvUvgRPzM7ThvSEU2GeXaMSTosWiyTA0DhJUv33SU/snkhP7JEIT1ysM0wU+xmjOcZ+9YRw5ntQkcE7P0dx5pTQnAoqLmjIJxUn9H78ZnGf4yKuJHiOLInyHF9XwHN0nsdzdE2E5OwI9xxbF+45NDvSs3+yzFgEmX8P9aJwCi/0p3k1YLQTZrBLyb5Ibhtfngf1OlEhgT2hLJUTPBgLIiPnqKMhrfgMN2c4KNioFwl1ucb8VDijPgf19HdIxQfO857+aYcHntbHawMPLcQKRA7EDQQM9rIz14a259xZIcHM28JH3l6MgBEwAkbACBgBI2AEEiVggoVtECNgBIxAiAk88NRzPfBY+Kx3z5cD5a0gRBFG2lOOp55PiHuFDo2kvngCvP/ai13wUlBhw5+QgFjBk92aeDep6R2Xx7Kpg7Dy8nuffnWRxJHp89bLz3Muf4ELvQKKP2GE8DSEpULk0HvgBTJ49O8zurz8Vm/nfUWMqU//c/85Hbefp8F7vfp8Z5IxP/vKOx86DbOEbfp+0j+LEXDwiMAontQcknMdQzr1Dsjj/jfcdkeHNz78fDDheojhrx4vUTmjvIYZNYo6+00PTjCqVrNOPeXkb16VJcwR58lxkZx5J1UHIzd1LrvyurZat27Dps0fe67HmzP+/P1X9pK/0EEaSgqehEbqP/znSaxZj6cfuU9FDPqLypkzpztcEudf7Nm779c//vY3YYv4zN4hXwZP4rtzPiQ1B3/XZVtiSPPg3eHvemr3gwoSP3476Et//ZNwm/PiVLXVef2QT7AsUfqSspyHL4LmBAnRVKxk6UvIS8P8SVo+ef5ajMxnjjXLly3mA+HjCEPlvi9hmcpISKirbvjP7QM+/eBt9Xxx1iPMG58Ro5znESe5J0mw9XxSDKmXVJ0adeo1jJJN4NwT2n9KWGxcd1qAco+fPfv6B/0H4RGSkv0SbBuH4VXFCjUkY6zVp/Y1XA7X9Ol5DNMYyPndxQCtRnjNdeE19qd10mKf8f2A9I1B/rh4HpzynNh03HNs5TEJDRUrQsQpz6onjnvW9Yj1LLvvlGfloyc9a7omeA5Oj/McnBHrOTCdnBYJnqMLIj0HZpz0xEiKjBjxYDi1M8oT69U8VVTQ5NdqDFfxgjpO47UmHXeKF1pHxQ36UkO7tj2dd+Lk9mMyrhyeA3/l9hxfFe45Mv+UJBmP8sQfFg+RIyKoHIj37BkfJ/OjvbNf1oECbwbOGmC0R9SBzYFQCxWuveYMC6Yhw3Q8On83Q82HokIX7OGNGKn7kHkhQqt3huu23o+0wxuCQ8NC+aun584SH3z9F5ZXRAz10nAK3/Tt/C5YiKjE6No1I2AEjIARMAJGwAgYgTMENC6qITECRsAIGIEQEGh62RVXE3aIrv/3+LPd6jW+9LK/fhv/M0bZI4cOHiSsEmF1br/n/ocJleT0qJBH7NdgxO0l4aIIAfPz98MG/Sl16Isn0Xk9Io+uu4dduXpNr0E7qaTe2o6wUQgqYnD+vUHTFq1efvrh+3bv3L5N74MxXyLNeJ/Kdh5jRg4bxJPevb8Y9uOwAZ/1uUAs2A936fYqycJ7vtj5EWfdqjWivTk15s+aMU3PY+hFjHi060tvEC7qO0laTL6Ox6VPOGDo7Tds9G+NmrdqPfzrzz9556VnHk/NEu3ecXpOo36ftZRwPcz78Q63tSEJt/aruQM6d3+zl0TfWeYUBdKDU1mxchMSaPmSBfKosP+DnBBcOe4QtFLD5Z+//viN5N3kLZHoUAVEX8jV4cEnn2HdP3zzpa4DRVQQm7rz6Vvv7Qj7RJ12HTo9cssd93ZCeOgtgtqvY0YOd44HpuyvBzu/8HL/D956Va+R44J9/eWIX6ZsWLd6JXuPp/GfFe+M1MxH24ouQEgXz6133feA6IH7m7S44qp2He5/uOtDHdvNmzV9amr3Ax5DGP+dCa2d41YvowP79pL8+MyB58wuiTlGwm+8LK5qe0s7cXbI/dn7PV/+Ycqc5fNnTp/aZ8B3Y/iteK3r496E53osWzx/Lu/3Cny8stycCOuFyIfAOKhfn/f8ceT+5D/pKAm5d2zdvIn93/Lq62+8/j/t7iKk1E/fDRmQXIbUU87smXkz//6Lflpedf2N1zWpUQbvHfVEqV6rbv1e/YeMbHdV02j1vkkJi0m/jB713Ovvffz8670+7te75yuEiLrh1jvuYY+tWrZ44WHpPC32T1J9ICj4PCswwmooI22m4gOf+W9tigoV+rCQhgPimua0UIOw0zMhqaEk+7ovabTXwy9hkteYreF+1LitBvBYCadEHgjGcdKzbyLjwviMIV3FlzhPgUbhnmJ3RHlyV4j35CwTLwm9T3nC8+YQ1yDmiAHc6TXiznfhDOvkZMLwnB4n/4bLiosVTuLNcmK1eIOczO+JOxom3h/SVnTmqAtzikghynseES+WJHj2/XpKhAz60cTe3E9/x7gfv/u88m/bKWFz5t+BZANNm4rqYaEeOOwF3VOsC9w0P4R68LB2mutDOWoYJ/VSwftBPXjcQgPCFffFi0IPf54Weo0xae4M3c9cY1wUhB/OI14QxpIxqBDDOLmu4b28Ap0791VaC3RpszTWixEwAkbACBgBI2AEjIARMAJGwAgYgSxIYPCYyf/8/Peitf/t+MCjJJnmqf4Zq3Yenb/5UIKzfDrkh/E8pe5EQIz6KYs37qXe+18M/cEZ158nrDmPAdCNDcPzj1PmrsBwmRykPFE9b9PB+LkbD8T932NdXnC2+c8dHf/HffDwcPdFOKivRo7/0zmPX2ev2OJ8QlvbdHvrw36z1+894xni7Atvh0nzVm/XfuBzZZubb8PQqefGTF3gfSo8NQfhh0ZNnrV02vJth97rN/h7QhL56++xrj3eZKwYXZ3X04MTXjTM+dqbbrsj0FxZc9aKpM+p4eFsi3Awa92ek8r7lxlLNyC2Ueejr78fy2d/93r8uZd7wpP1YR391UEc4vq346eeJcKwP5977b2P2Hvw7v/tmEkksE6rOdHPq70/G+jcn9xDvZNSux+GjvtztnuPOMc+8IeJ0ybOWXmWd4Veb9bqymvhxti++/XvBYg9jIvPczfsj+WcO1wWbRF0aIfY4Y9TBxEhaN/yqn+9ZfzVQwyZvnLHEWVDn8+JAODvO5EYQ/omV8iI32Ys0r5YSzw1nHPl2pz1+2Ke7tHTmxPFeaSEBfN3ruv4mcs2kWQcT4603D9J9SVGVxJk55CSW0pOKVFS8ki5UEo+3/uC8lpYSiHHeepTLnLU0/aRCCHpFTpHhIuLpFwspYqUolIqSakspazvtarvtZy8VpRSQQrvqVcm4c+CVRMWt6+csKl3tYRdo6okHJpTOeHkrkoJcbHlZQ6VpVSTUt33Gi2vlNpS6kqp5yh8ptTxXdfXmglxcdEJMYerJxxaWCXh+MbohCMLoxP2T66VsGd87YQD02om7P4lOmHrF9UTFt1WJWHhLTLeMMbHHHTsOhfGzByZK3M+69/cpNY7VNd9681eyuXYD+wj9sgFUopKuUTKxVJKSKkopYqDLe9hrczhW9XHtr6PayN5pfC5tK8+n2v6eOt1Xhv46uo51on+arnO63XWirXjM2ut68r5Sr7x833g+0Hx7m9nCRVb69cIGAEjYASMgBEwAkYgcxJIljErc07NRm0EjIAROP8E8CDgaWJn/H8M/XUaNLm0cLHiJXi6WcISzQ+UHJuwO/ShYXucM+rx7sdfLJNY9yO/GXBWHgieVOep7mByHCCAnDp58oQ79BP3f/X9zwYO7Nv7bRIiu4kSwogQTkVLlCxNeKp58nS4O9cBbcpKmBoEmEB5NQiLUy26Tn25XeEl8+fO4glywkTVF8Pq6x/2H0zfHW5q3TS9VpSE03GxsRrC5cxtQ80J7wqEmqUL580mlYO/+SJs4Xmj+QzSigl9VpNcA3hOSALlJZokmxBUrN/En38YkZp7BWJKSDExXCXwdH9q+g/UlrGzj7du2rhePYeCvU+gsSfWzwUScwrPCX/h1GhHzg/GtmrZkoVxstmeeOHVtzG6/zR88FdvdevyaKAk5bQTh6dzPKvok98WhCwN+5TU+GrUrteQ0HN49CTmsZMUQ76/lapVr8WrOMssd4+P3yRCOQXinxIWJGcvL+Hv8MRatXzJorTIe5LcfYHBVeo6PSvUW0K74KlznubnCXnNP8BT8eqdoCGJqMM5Z34C+vB6XCRTc07usAPWE8M9YyCkDzkLGJMmxuapeUIN6RP+6u3A+DRUE0/Pn/aeyCd6Y6knIj0Jx8I8+cTRL1IeuI/IHSMlzBNVTL0o6FPzfejcnWG1TnscnNp3Urw1cnkSDsZ5TuyI9yQcCvdEFgzzHF0V74mQZODh0mfc0XjPiS0kBxd/jj0xng3vxXhObde1gKmOXb09NFk13gKHfR4nqeaXFh349pR6LOge0HBK7B3Whd9I1gh+nNMcH04PCEQY9RyhLl4UmvODHBQc6hERyNP+tGfNv+GiaAOzxPLeqAcFzNUDhHaEPtslhd8sTcqtSdvPeBKl115Pi7WyPoyAETACRsAIGAEjYARCT8AEi9AztjsYASNgBIxACglE12/UdNBPk6Z/8u5r3b76uFfPFHZjzYxAhiWAV0PPj78c2ujSllcwyNZ1KxTdt2c3Br5sd2QGFg6xQo3umsRZjbGsmxqUMfpSODBGa54HfY9RXcP2YMTl8IbMEQNuSMJCJbapRLhgLIxNk17zSi4YDT9Ecw0f5UywrXkQuC7jjozwXHzFSU/Bq6Mkn0SEJ2cpMX2XSvAcW3PCU+Q/EjIqfw7JQSFhpIrl9MQfiRNhQvqPkHmHh3lOSRiq8JwRnliJ7BV7SBJ+n5LrOcM8x5ZHeHJVFDJi/w73DTPuWKznyOI4z6G/wzx7xsKLsE7qZaNhtjCUqzHdO2YRKs4Ro8/3lw1vAx9nzbnhFIUQLhALEBpYC+YIc+ahydvZN9ThGp0R6orrKmAgdqhgARPNb+GcOnUIJeXv0JwkmpciOcgYg45DvyfsH9bpLEHeBIvk4LQ6RsAIGAEjYASMgBHIPgRMsMg+a20zNQJGwAhkOgKE8Kleu16DG5rVKq9x7zPdJGzARiAAgYbNLrv8rU++GiapJ7Zvl0z0JC2/tlG10tkRWGZg4RArWCLNiYChmEPzC+hnFSIwAvN0vD4Rj9FZE3M7n/zXp/9DknQ7JXtKBAwOfUofQ7Xmg2D8zA/jM0/eI2qoAVpfuR7nCYvIKd4VYSIyxHkiLhRm4fKaR+rER4hQEeYp2DrCc2SliBcXxXsKt8/pOblFJAXxkjgs+eWjColZvnS8J2Z/mCe3CB6nDiRI23BPziJhngNT4z3bBuzznNqj49Kk0awD49LE5sdFoMgUh0+0UK8KOMJeE2rjKUGeCc6zDggLKiwhcmjeFE2yTTvdk5rXQjng9eDMXxEMH02Wnpw21NVE4Igk3JdxIlioeOftxwSL5OC0OkbACBgBI2AEjIARyD4ELOl29llrm6kRMAJGIFMRIGcECbff7v7MYyZWZKqls8EmQYD8HeSLeaRLt9cmjBk1nOTafYf++Csh3rIbvEzIAqHCKypIUcGB/57WpNS816fceSpdhQ2M/GrMV8Mzy639aPLlDLMFfIb+4yJcIABouCKnEZ2xYjTXRNHMSz00TnsIJMRJ8u6tvjBNG52hn04n5t4/Sb1MJGjQglhJ4B3hyVtLQkpVEclhc4Ln6HLJbh4TLx4Z4Z5TEhpq/+Sjnpg9msRcQ0ppwmxECgQUuONJ4TesXoYB7BqIL5G7stRk2rzqfFWY0KTW8GbOiA8w4DPiEXuRNuzPg1I0cbfuUxUruKZeF8nFoqG9EquvYbmoy1gQLdhDuj+ciebPEi6SOwirZwSMgBEwAkbACBgBI5C1CZhgkbXX12ZnBIyAEciUBCRNw8Xd3+rTb/7sGdNGDP6ib6achA3aCPghQJLqNz/68psWV1zTpvcb3Z4Z+mXfDzHaV5FcIV/3/fDd7AQtE7LQvBVqeFfDL0Z3Pcd/W6s4ocZnjLX6tDv1MKirod4bAkrX/XyEgkpqz/kM/xjGKYdEwGAu5LzA2I3nCIZonT/X1DDNvE7nt/g3V8eZqcobNX6f9vje/4cIEn+IATtc2sRrSCz4UE89U6hL/1zn3rDE8E5OCvVuSWpKGfY66+/ztFDPCs2XwpidQoCGuVJhQvOQUI/9xnWYIRZoaC/9u4/zEnPL2x/nUuptEYij04NfPYc0D4rmPkFY0nXMsOthAzMCRsAIGAEjYASMgBE4PwRMsDg/3O2uRsAIGAEjkAiBtrff2TEqZ85czz9yX3u13hgwI5DZCWCg/3TIjxNIbv7U/e1vmjZ54i/MiUTrJJ5etmhetvGwyOgsfEZjlkcNxvqk++lQR6cP3mN45Ul2nnp3JtHGKMzBOa5TDwM7Hgr6xLzG9adepnnS3CcMHBDhgjA/zEeya58ZP0/6YyDHGK3Ju53eI2rMRmhQwYL3KmwQLkrDDqmXAX3B3NknzLbBNbN5Uvj2RcAXh2ihYg112T/q3cNn2HFO84eo146y15Bk9KEhyHivQgi8OQ979q7+TahCUWrCBnMf+tfk3Rf67qN7g3uy9zOVB0xS62bXjYARMAJGwAgYASNgBNKOgAkWacfSejICRsAIGIE0IvD9kAH9Rn/3zcDDhw4eSKMurRsjcN4J9Hj34y9IJN/ZIVYwqLqNmrVAmFs0b/Y/532Q6TSATMLC6TUAGYzBTi8Lzml4KDW4q7eBGokxKPPEuybVpg11MTaf5V2RTujT8jb69PxOHxfmjIDBU/QYpzU0kXpc6Dllo6GcEHI4YITQw2f4qNjDOfrkuvPJ/MzOL+Ba+MJDOYUeFXE4Ry4I2DB/Fcw0/BjeErynjgocugc1h4RTpODfWGei7cSECtppUvDE9hHj0j2v+5x74+2BOKICVGJ92DUjYASMgBEwAkbACBiBbEzABItsvPg2dSNgBIxARiVw8sTx45SMOj4blxEIlkCDpi1aXXPjbe2/+eLTD/6aNGGss32zVldeu271imVHRKELtt/MWD8jsnB4VChS9axApDg7dNG/nhT8dzShkUisjUFWwxRRX58w57yGhNIny/Ua9/KG+cmIoaCS2lu+HBdnhBjxuIAZexguFMQLNVDTHXU1ZwfX1fiNAVuTZmPUdnqnaGJvrntzhsh91QsgqSFm6uu+RNTeufoSvqtHAudUGNPQUCo0aJgl9ph6AmmIKA2nxf7kmooc7FHNu4K4oZ4t7nwV7POLA0BVrwoua74T+qHNXikaHkxFKvUycs4pU6+XDd4IGAEjYASMgBEwAkYg7QiYYJF2LK0nI2AEjIARMAJGwAj4JdDm1vb34EUxqF+f95wVCI3UWJLLf//NV/2yC7pMwEKNvypWqBEXo6yG2NGQO9TBIwDDrIbwwQirXgRqpGd51biv/WtOgky/9I68C8wlVoztiAte4cEnZOQUocGbU0E+e70DNJSTfPYKPPIZYzv1vR4BAYSJbCFW+NkQznk7Q0OpuKBNECec4cVUuFDPIPXIUK8XFYTUY4PwTbpXtQ17nXwlvAZK1K0eRs6he5Of+05oUnrqqQeN0+so038HbAJGwAgYASNgBIyAETACaUfABIu0Y2k9GQEjYASMgBEwAkbAL4Ey5StWPrBv7549u3Zsd1a47uZ2d+bKnTvPlAljf8ou6DI4C3fOCgysaiD2PuEvRYUL3mMA1lwNmlgYQyyiRQGHcZbl1bbupc7wRng/Hig6H6f4ovPyph7yeQh4fMKDek3w2StM6OETLv5NPH5a2LDDySjsrEhNzv2iHhi6Hv7yQji9KXQv0w7OmtMCDwsNu0V98pMgLLD/ERvY57xXDxrOqUihHkS8InxoSDBn2DNNDs591MPIvCtslxsBI2AEjIARMAJGwAj4JWCChW0MI2AEjIARMAJGwAiEmMDxo0eP5M2XL39EZGRkXGwshm8Pibb/9/iz3davXrl8/uwZ00I8hAzTfSZgoaFweMX4yqsmCcbYqqGdiP3PdYywGGv572reUzAMaxJuDYOjn/WpeG/SbTXsZ5gF8jMQ5xh94Yk0vwe14aO5PM4Y032iRYYXYzIy9yDH5vbCoLk/AUM9h3Qf8qohtzSxuYaWYl+zfxEqCPGFCEHYrkJSCrJ/pez3vWrYJ/a5hkjjHP3zneC+9KUin+6bIKdp1Y2AETACRsAIGAEjYASyOgF3bNKsPl+bnxEwAkbACBgBI2AE0p3A1N8njIvKmSvXnf/38JN4VFSqWqPWx4NHjitWstQln/d553XvI+nZ5MigLJw5K/Rxdk10zH8vOxNK83Q5uSsQLC6SQqJjirbjCXVnYmH1rFARg5X2GpIzg1jh3JY+sUIN3pqEXOfD/DR/BbzCqZ+NtvZ5+wazj1wFIeyc4hsge89ZdL8iTmjOFaoiLKhgwStFRQ7q7fEVvDH4zJ5XgQIhj72AlxHfE/VUoo8smyz9vG0Au7ERMAJGwAgYASNgBLIYgbP8i7PY3Gw6RsAIGAEjYASMgBHIEAQiI3Pk+HDA8NGXXn7Vdc4B/fTdkAGvPvPo/RlikOk0iIzIwmeIh4B6Veh/I6s3siY3RqjQhNHU1cTFPKGOgVefLsdAq0+ka+gdzqmh2JtnIDMJFj7hQcUKxq/ihBqgNW+HflavlPjMmFQ8nb4OGeI2DlFJPWecD7Vp3hYNeabiqnoS4TWBWKFhpdj3mtibtl6PMjlUGFEPJT57+8pM34MMsWA2CCNgBIyAETACRsAIZHECJlhk8QW26RkBI2AEjIARMAIZg0B4RETEtTfe2r5xi8uvxKPir9/G/zx5ws8/ZozRpe8oMhILV4gjp2CBQZX/VtaEwYgNvMfIivhAXcLjYKDVhNtqqMW4y4FYQVHjPeecSZG9lTK6wdZn0HYas5k/goUmdWZ+mstD53dGnJH5+QtNlL6bzu4WkIBLsPBXT4UqZ/4JvIr0M+vPd0C/Fxoeis+ak0TDTDlFO+/3IaPvf9s6RsAIGAEjYASMgBEwAulLwASL9OVtdzMCRsAIGAEjYASMgBHIIAQcIY6cORkYHd4CGORJPIz4oB4WCBSEtcGAq9ecsfg1bA5Pm+sT5WrMdYaJOisEWEY32Lq8K5xeFrDRpM5uAUPzWiDIZJuQZxlka6dqGK4wXvr3ovvvRvWw4V7qSeHcG7zXnC8acu0sDyO5bh4WqVopa2wEjIARMAJGwAgYgaxJwJJuZ811tVkZASNgBIyAETACRsAIBEfA6SWhxnfC3WBkxTCPcRXDK2GheI8o4XziXA24CBOEh+JVExqroTYzG++dooN6myDsqBCjT9c7OdAmzpejhdBQwa2I1T4vBFzrpCl2dP11EXXd+aweNGfCPMk5b1J53wQ034l635zjZXReJmo3NQJGwAgYASNgBIyAEciQBEywyJDLYoMyAkbACBgBI2AEjIARCDUBnvx3JDzXUE8aix8D/BEpmoOC2Pv8tzOhcFTcYIh4VXCedhwqbGiYJM6pITczexpgmNZQUMzXm1hbCsZq5q6flaMasc94WoR6Pa3/dCHgFq70pipk6P5XrwpniDBvXfO4SZd1spsYASNgBIyAETACRiDTEjDBItMunQ3cCBgBI2AEjIARMAJGIDUERKzQsDXup8R5ely9JzC44mGh/92sYoUm0dZkxLQhZJTWdyYbzsxChdfG7OAMM+ZGgYkyZI6ax0LFCtpRB2YclssiNRv2PLVNxDPGu69dIaTcnhj6ObN/B84TfbutETACRsAIGAEjYASyHwETLLLfmtuMjYARMAJGwAgYASOQ7Qk4km2r54B6CWhOBvUM0GTB/Hcz7wkThZcF9dUIi/cFnhbqXaAx/Z2hb7JCcmHmo/k81KMC4UJDZjFvOKmIo/k78FLBnSXDJxjP9l+MFADwCRpuQcIEihSwtCZGwAgYASNgBIyAETAC/z4pZiyMgBEwAkbACBgBI2AEjEC2IOATK5irN8eCFDwDMLIjSGjsfUQIrpNcG5ECjwrqUFfbcp2wUUd959Tr4kzOCs5nkRA4mpic+eeWgmDBwWfeM2dY8qrhgODhzGXA+TQ37v1EzwAAIABJREFUZAdIEu1F77xfFlkHH3Z7MQJGwAgYASNgBIyAETACWZOA/sGVNWdnszICRsAIGAEj4CIQERkZmS9/gQsMjBFISwJFipUoWbJ0mXLB9kmbuzs92jnYdtmpfo4cUVHFSpQqHcI5q3GdW2jCaPUQwIuCJNu8YojHAI+AgREerwHNTcE1TSyM0MF1Z0z/EA4/3bpWIYJX5qhhnpy5ChB81AND2fDqZBzKAet9nOKKrgMeHt4SygFY30bACBgBI2AEjIARMAJGwAikjoAJFqnjZ62NgBEwAkYgmQTa3/vAY916fvBZMquHrNrd/3u08+/z1+y4uFDhIiG7STbqGAFo+IRp81tff9Ot2Wja50z1kyGjxt/78FNdg2Vw7yOdn+v40JPPBtsuO9VH0Bnx24xFIZiz07itRuxcch8ECfWmUA8M9ZzA04L/ftZ8FRjnNQSSJqCmruZySHNvghBwCKZL9RxBsNB8FDBBoGHeKlLAkxBZHOkVglZFCsaBx4eugzNZuHedTbgIZsmtrhEwAkbACBgBI2AEjIARSF8CJlikL2+7mxEwAkYg2xL4v8e6vBCZI4eGEDlvHGrVbdA4UgZy7OgRwrjYkUoC5SpUrlqlRnSdiwoWKpzKrjJt8/CIiIjyFatU279vz+5gJ1GhSrUaWzdtXB9su+xUv36T5i2PHDp0MARzVkO25mXQ3BUY49VLAkP8cSlqDEeooKgHhuaooJ7mvGCoXmM+sf0TSVgcgimFrEtNnq3iDDk8lIH+rvOZ88ydc3zmUOHAySetB6rikzMBOOvpTJCuHjC67uEiXESYx0VaL4X1ZwSMgBEwAkbACBgBI2AEUkfABIvU8bPWRsAIGAEjkAwChYsWL0FZOGfm9GRUD2mVStVqRq9dtXzpiePHeSrYjlQSqNOoaXO6WL965fJUdpVpm8vWLoWnya4d27cGMwmEjqo1atddNG/WjGDaZbe6NevUb7R4/uyZIZo3goPmOcAjgN8FzmFsV68BwkHpU/v8t7Mm16aOJtdWg7kayb3GeVduhRBNId26VXHGGd6JecJBPVQQKshvoaG1VMhhkN526cBEx6IeIOr5oQnB8aJxiucaKooF8xY7jIARMAJGwAgYASNgBIyAETh/BEywOH/s7c5GwAgYgWxDoHp03QZMdtG82f+cz0nnzpMnb6ky5SosW7xg7vkcR1a6d+16jZpilV25dNGCrDSvYOZSsnRZb+6KHdu2bA6mXbWateuxJ2dOm/J7MO2yU12+rxdcdHHBJfPnhEKwUM8KNcSDVp/CV08CPC32SdGwR3hmHZJywPGKxwXtNK+DGsqzineFbjnlhccJ+Ts4OIcowfw5R4EVog7v1TNDRaFQ5Y9QEUXzbKjAxDpqeK988h5xxRnCSwUrXffTk/IJFyZgZKdfG5urETACRsAIGAEjYASMQEYhkF4xZTPKfG0cRsAIGAEjcB4I1KhTr+HRI4cPbVi7asV5uP2ZW1auXqt2uBxLF8ybfT7HkZXuXVNCbG3esG6NLG8oQvZkClTFS5Uuw0C3b9m8MZgB16rXsAn1ly60/RiIG94VXFu8ICSChfu2mjhbjfGat4J6iBEabkgTS/NZc1XouTOP52eRUFBORjpfNfirlwKcOPBgQMzgVb0aEC7wUEHUUHEgmK9JMHVVFKGNvtcxI1QwXh0jXiDkKtHE4YxPvWV0DZ39BTMOq2sEjIARMAJGwAgYASNgBIxAKgiYh0Uq4FlTI2AEjIARSB6BGtH1GixfvGBevBzJaxGaWjzRTs/LFs2bE5o7ZK9e8+bLX6BM+YqVs7vBvWixkqVY+W1bNm4IZgdUqFytxv69e3Yf2Ld3TzDtslPd6HqNmsTFxsYuX7xwXlrOW8QEp1eFGtL5fUKYQHzglfMqWmDM1hwM6jWg1zQR9ZkhZkGxQhlh+EeA0HwfatyHhYoACAGIAwWkUJ86KhykiYeFywNC+9R1ceaqYKz6gJauJyGhdKwqQjF+8m9wjfqasyRNxpuWe9f6MgJGwAgYASNgBIyAETACWZ2ACRZZfYVtfkbACBiBDECgRu16DZctmn/eRYKqterUi4k5dWr18qWLMgCWTD+EasJTDLNhSxbMmZXpJ5OKCZDDQvJt7zp+7NjRYLq5pFyFShvXrVkVTJvsVhcPHkk5s+ikJJ0JwdyduQ6cybN5r0ZrDSnEOYz0TqGDp/L1yfzskPgAYYb5EvIJLxTlgShB4e8K5QVbRAuEAGfYJZYx1SKAJjP3veqaaP4QvDp4j1jBNb6XjJsDMQVhQkNIaaJwziNW5PddV6FD90EItp91aQSMgBEwAkbACBgBI2AEjIA/AiZY2L4wAkbACBiBkBIodUnZ8sSgX7bw/AsW1WvVqb9mxfIlp06dxKBlRyoJqMfKkgVzs7VgUbzUJWW2bFy/NlicCBaE0wq2XXapHxWVM2fVmtF1lywIacJtFRo0NJCGAeIznha86jk+q7eA06tC+8jKooWKDmrox8CvQoV6MCBO8F5ZKisNB6UeKqHYwipaOL05uB/iiq6lzoHxIIBxHU8LFVsYF3NgjggWmpw7Qjw6zkrMHYoJWJ9GwAgYASNgBIyAETACRsAInCZggoXtBCNgBIyAEQgpAZ6Q5gbLFs8/r4muo3LmylW+UtXqSxfOtfwVabTiVWrWrhsbGxOzYsmi+WnUZabshhwWwQoPOXJERRUpVqJksO0yJaAUDrpqrdr14LQ4NAm3SYjt9JZglBiqnfkYNIk29TRUlBrdNUSUV7igL+dT/ymccoZp5ifkkjMZOYZ8/TtC/5ZQMQcxmKKhlvBmQBTg8xmRJ4RJrXU8uo54eXB/DhWgECO4zjg5h4DB+qrXCNdUfEGA0aJiTYZZJxuIETACRsAIGAEjYASMgBHIigRMsMiKq2pzMgJGwAhkIAI1atdvSELmlDyBjmdG6+tuvCVP3rz5UjslntSOiIyMzKz5FiRdxAV1GzZtnhQH5nj5NTfcXKxEqdJJ1U3tdZgSXuvUyROapDi1XXrKVqhUpUXra9qkuqN06oCQWMVLXlJGHCxWB3PLEqUvKUsC+C2b1q8L1C491zKYsadX3WhfUvIl80PnweMTLZiSGtOdngT638lOzwkVORAp4qSE0msgvVCfcx8/IZeUj+b3QLBRPrzHk4GiooAKGOqt4MwzEep5sUa6LnhPqMCCUKG5NPg3hfBPCBoUhBXqqlcGr5pcHG8SFTkYO94WHmcJ9YSsfyNgBIyAETACRsAIGAEjkJ0ImGCRnVbb5moEjEC2IlCpWs3ojDDhGnXqNVy5dNECMe4EFS4FY+3QcX/O7vX5N6Pa3nZXx9TOhXBQ9LE0heGLylasXJUQNakdR0rb3/dI5+cG/PDr1K9//O3vxMSIV9//bGDvL4f92KVHz94pvVdy2ol+cmG5ilWqiQCUZrlJ8ID5buL0hR99/f1YElInZxznuw5eErnz5Mm7KUjBoqSESmPsWzZtCChYpNdanm+Gge6Pd9ZRUTs3rF21IpRjdIgWTkO3M1SUM+E2nhlej4pQjikD9q1JqDHk8zuoXhMMVUUJvBL0bwv1sOA64gViQHrkg2B8HIyFcSJGcF/Gq54Sep3P6jlCPR2zhrSiDUKGhr/S8ZunRQbcoDYkI2AEjIARMAJGwAgYgaxDwASLrLOWNhMjYASMwBkCbW75793DJ0ybHxmZAyPMeTsQHarVrFNv+eKF84IdBGMXm/hFCB0b1q1eGWx7d308PSRv77G1q1csC7Yv8nB8/9uMRXUaNrk02LZpVX/Ap73fHjvy28G1GzRuNuTnyTOLFi9Zyl/fFxcqXITz60Ns5I2u36gpHgJpmUw9/wUXXEgIIDxy9uzasT2t2IWyH/JQ0P+m9auDSp5dsnTZcrTbmohgkV5rGUo+qem7Zp0GjURgnB2s2JnCezpzIKg3gSaVpktCPnmLu3+8EbLBoeGy1KhPGCUNocQ1mBFiCT6IBQgUemgybmeuiFAhcwpNCCV4fRDuibGRt4L3vGoSdT6TlPuI75wm3ta1Z+zqVeLMj6GeGtli8UO1WNavETACRsAIGAEjYASMgBEwAkbACBgBI5BNCPQd+tOvI8TAfr6nW6VGdJ35mw8lIKCkZCwFCxUpGsgwH2x/P0yevQwPhWDbUf//HuvywrxNB+MJUZWS9mnZ5uq2t7RjLJ9+8+MEf/3ytD9hldLynv76eqxrjzdZ22o+z5W0ul+pMuUq4L2RVv2Fup/b7/nfw3AINmzZU91ef3f6yh0YSQMe6bWWoWaUkv75rsH18ede7pmS9sG2cYf48X0+E/on2P6yWn1f0ukoec0r5UIphaUUl1JUShlf0c+5fOdLyGsRKbwWlMJ5TWCdpiGVXOsXLp8jfffifoybz9yfcZSUUklKBSmFpFziK+V853lFLGfcpX3XmFs+KXl8fWn/3j1ihxEwAkbACBgBI2AEjIARMAJpRwDXZjuMgBEwAkYgCxHAM6F+k0tb/jR88Ffne1o1atdryBhSmpR5755dO9NiDnnz5ctfRoz4077q+2FK+mvS4vKr1q9Zufzg/n17U9I+LdtM/PmHEaxvuw6dHiGE0jqXx8jxY8eOblibeo+UpMZct1HT5vFxcXFrVy5fklTdYK6nJNdJMP2ndd3q0XXq79qxbeuxo0fPEh/CIyIiipcodQkhowoXK16icNFiJcRh6OL8BS68EEGmXuNLL4uIjIhERCPUWA5xLcG7JEfOf9/LUh656bK6ldN6zJmhP/3tWJLCEG7BzjGAl4RZos8GiReFhksi/4MmtuaV8xTCMBFCScNr4eGg4ZZonx4eCZq/Qj09eFXPDzwjnEnBOc+Ynbk5NOQV3hcFpBAaCm+Sg745MgdnrhMo2V4J9ktn9Y2AETACRsAIGAEjYASMQAACJljY1jACRsAIpDMBnpqWHMXH4+UIxa0JUYMBNFhDH0JHbGwMRps0OzA6EoYpJeGJyI9wYP/ePfL/3UkNiNBT8pRrAgZ0f3UJB0X4oqUpTN5bsUr1mlMn/zouqXGk1/VvB/T7CMGi5VXXtXUKFoQQKiBG8Q1r/Mf8hxPrfFIWJTVjxbDO2ko0ozWnTp3E+JcmRy1Jsrx80YK5gfYh3jY7t2/dkiY3S6NOqtasXW/7ls0bESBIEg2XcpWqVCtdtnxFd84T5nXk0KGDEvHqQMEiRYrxeurEiRNHDx8+BMcYKaf4n7xGhEeEr1uzckWgPZ0rd+48OXPmynXwwP59aTSVM92Esm/nWBP7zakRXa8BdRfPnzMzredn/SVNwOU1oPkrNB8E4aD03wqM+hTq8HeF5rHQMFB8pmj+h5D8u5fIjPg3QQULqhH+CfGB0E+FpCCucDB+fhcRYhgrSbn5zJydYoTORcPqwiGGf36c9bJJmLCkN5LVMAJGwAgYASNgBIyAETACRsAIGAEjYAQyPoGf/1609okXXn1bR9rq6jY3fTZs9MRhv/w153+PP9vN3wx4MvuRZ7u/Pnj07zNGSFLiJ55/5S2Mxlq3liSn/WTwqF/6DBzx88AfJk4jlMoXI8b90av/kJHv9Rv8/au9PxsYKInxFde2/Q/ho2gzavKspcVKlrokrSh+O37qvEE/TZoebH9i7AmbtnzrQZJHJ9a2cvVatft/O2bS3A37Y2eu2XW8/b0PPOavPgmrmZ888F5Wr5OUvOur7/Z57vVeH7vZXHhxwULvfjZoxMeDRo774Ktvf6LtyN9nLlGePT/+aijrFuy8tD7iSbe3PuynT5G7+0FY6D/859/rNWrWItA9pizeuPeFN9//1Hn9wwHfjflj4frdtPfX7pX3+w4YPGbyP3qNeTPP7379e8HL733yZd58+Xma+KwDFo880+21r0ZN+It9wj4klwdM2FspZeBuV61W7Xr0eef9Dz/pr0/Weu7GA3GIGnqd8T7do+f7E2Yt3zxp3urtzvWH8S133tuJdYPVjbffdW9ajZV+ChUpVpx9NXv93lOMm8IeZM+zPzo9+dxL1918+531mzRviYiIUKn3P72/tx3q3P2N9wKNKam1JBm9OywYnkCsE98dvv+FixYvof0joLzR54shfy3dvP+rkeP/JD9MoHuHsm/umZzfnA8HDB/NuqblmllfySfgCrFE2CMKwnB+X1iki+W1jJRSUnhPmCjCQxFCibBLvC/vC6dU1veZ9tpXmoaEcs/MN37nuHPKOQ1JRZioAr7xVZZXwkMxxgukECaqppRaUqpLqeL7zHtCRFGHcFiEumKOfD4n1FXySVtNI2AEjIARMAJGwAgYASNgBNwELOm27QkjYASMQDoSQHgggbPeEuEBg3jlajVrFy9Zusy9jzzV1Z0oG6P2D3/MWd7pia7dCTMTGxsXe9+jTz//2HM93tR+yBWB8TYm5tQpSftQjCe5c8pj0uQDIBRS2fKVqsiD9eck4L734ae6vv/F0B+OSzib4QP7f0z9Bzu/8HJaIOHp8opVq9dMSVJmMQAl7N65YzvjCTSWZq2uvJbk05eUq1hp6IDP+mzbvGnDky++/o4/Q2yNOvUb7duze9e2LZs20N9/Oz7w6Le//DW3/X0PPo6R223AZY2KlSx9SVxcbOzFBU8nsZa3sSUkUbKXZ4XKVfPmP9e4n1xuslQX3Hb3/z14d6fHOvtrU13yQjS6tOUVTVpecXWgPnk6P2++AmcJDLt3bt+GwCARsM4RHuinenRd71PrHC2vuv7GYeP/mnvZldfekDd/gQI3/fee/5NtUs15P8QBko23v++hx3ds3bKJfcI+7P52n/7UW7Z4wdzkzjmpert27NhGndJlyvtd85qCBBFCtrjXowNvkkGjJ02/p9NjT8te2ZYrd968z4oAhTcM3zMEn+dee/ejNSuWLj4u8Zpe7Nm7b2qT0CM0NL3siqsRribMXLYJ4ZE++/V+65V72l7e+NKqJQvccV2Lei8+fv9dX/R55/XxP30/bO4/0/7ctH7takJ1KQP5qpcjTNnGdWsCJupOai3x5sAjQ/tkH5O7poKECZOwWusaNG3Rquur7/ThOjlkRkycsVD0qWjGgzcIHjqB1iSUfSf3N4ffvWC9xJLaY3Y9+QTwEHAUd7gj/fsBTwU8Di6QgkcCIjqFf2vwYEA45T1eCNRVr4v0+vtDx433A2Pg+8J7xsxvJOPgM54UeI0wBz0HLNrThnkwr4ulkMeIOdGHJmfXROS0scMIGAEjYASMgBEwAkbACBgBI2AEjIARMAKZh8Dl19xwM09iY/TE0Mr7Nz78fDBPXyNGuI3txUqUKs3T4ZPmr9mBkVFniifF1GVbDvh7kh6PA7w1kqKChwD3f/2D/oMwBFOfJ6vx4EiqbXKuY3BMTcJtnuZ/u+/A4f7uRe6GGat2HsVbAOM/dTDQcr+Hnn7hFXebiXNWbuWJdc7zpD313vpkwDCM+zzRz2eSJ/u7FwZ6klz78z5IDodAdcbNWLKeROB+7ylP5zMmvB4CtceTAiO88/pzr733EXvFXxuSGOOhQBJjhAg8A4b9MnWuep1cVLBQYWc7CXVUl6TQ7CW9hsH+0yE/jFePApinhoGzLSID/d52z/0P+esTbxiukxOC/fr5d2Mn41lz7U233UF9xAOu49mAVwVeIyp44cnANe6RkvFyP/bNmKkLVtMPXgxtb7+zI+vz55JN+/T7k9y+9XcgMQ+axNaS3wnG0ePdj7/gno2at2rN2uJdxTXESq6zRxDG5qzfF9PhwSeeYf34reEa/fsbbyj7Tu5vDmvMGPFgSS5TqxdaAqIhk8gaLwU8E0g8jWcBHgcksMarAk8LXvFQqOh7xWuhjBQ8MGhH+7OSVctnr6dFqA+5h3pb8EoSbrxAKDpuTbzN2KtJwbOC+TDHaCn1pdSRgjcG7UjWjZcFHie5peBlASNLwh3qxbT+jYARMAJGwAgYASNgBLI8gfR6winLg7QJGgEjYASSQ6Bxi1ZXnpIEFkeOHD705IuvvTNyyFf9uj/1QAeeviZWvTw0v1/7QcB48+Mvh+Kp8FD7G6+cN/Pvv/TanBlTp2Co50lt932r1qpTb+nCeYkKFiT9femdjz5fuXTRgte6Pt5J82lIWPw8eHAkZy5J1akm46BOSp6SJoZ+eclhsXTBvNnu+8Clp3DBm6Tz/XfcLChJhOqBD0+6/zb2p7PCFBHiitA4i+fP/oen77u9/WG/CaNHfstT8Af27d2zcM5Mb8iq4qVKl/E3p2qSVJkn4Y/KjZKaczDXVy9fsqh0ufIV/T313+rq62+kL2dIH2ffGJURWyTX81khc4R5fX/MaNuw2WWXY1ifP3vGtLc/HfjtqmVLFnZqd10r9Tpx5gqJktwI7/T9+jtyKTx5339v1GtijEsYM2Lo1/SHx8mSBXNmBTPnxOoydq4vXTD3nDXnfIUq1Wry3dkj7hS33X3/Q8zngze7P8tacl09iDo9+Wx3GfaJ+2+7rqUm8Bbh7xL2S0ryPZStWLnqIAnFRli1datXLr/7hlaN7r/12st+/n7YIIQfvovB5qMhHBljXiV7IBCTxNaSfUw7vIr4riCc7JS98OR97dryGxIpyby5zj55/vVen7zc5eH7Bvf/qBfrV6xEaW/INzj6u3eo+g7mN0c9geR3zO9eSKs9Z/0EJqBCgu9Vk0zzbwNeBfz9gMcEuSs0RwVeBySr1lwOXCPhNmoEeSK4TkmPpNuBJqa5OHjVvBuMX8+T7wJPKC1cY05HpHBNPS40l4cm9eZ+eHCcScSdHiKM7V8jYASMgBEwAkbACBgBI5BVCZhgkVVX1uZlBIxAhiRAPPsFYiDnaXGSyb7d49nHAw2U+Ps8gf3BG92fXbNy2RJnvWNiPeez+4lxYuVjpFw8b/aZPAX++u/40JPPElLnzReeeghDLnXw1pAQTrVWrwhsRA0GKsmID+7ftzexsDeB+qteq259xoPI4K5z6533PUAIrM/ef/PlvQ6jK0bj/h+89eraVcuXOtvUqtuwMZ8xhL/2Qb+vt27csO7VZx/9H8ZbzksqEG8uEBU+3PcjFFFSPIPhonU3rF29ErGiVJl/Q4RxDeFEDbaFixY7k4PgrDn58jisW7XijIcGfZEHItBY2XskQG/W8spr8oq7yNP/u/M/R0U58zd2wvawl7786N03CE3krHP48EGvQESoL/pLydz9talVr1ETkoGvXr7UrxEfQ/rqFcsWM/ZHu770xqy//5w89Mu+H2pfhD3zrqMktX7q/9rf5FzP8pWrVmfdgx3r1W1vaffdhGnz8TB5sH3b1k/9339vVCN6QVkccoDMmvbn78H2K1pcTRJ1B9pzSa1lBZ9gsWLpwvkdHnzyGcLJvdT5wY4qeJbxsUDcG9Svz3vjfvjuGx0jLHi/ZcP6tf7GHaq+g/nNqVGnXkO+n7LH0izkWLBrlN3r+wkJpeGcQEPopAv5+ZSCsR9jPtcRNAihxL8piGYY+/mdxZivxn/qhd6lwrWAMp8EKc6E34yZwngJCcXDAiSwZ6yMm0JYq9y+uXCe+SG+kKyb5Nx4bOGZxiuf4cH8vKKMiRauRbCPRsAIGAEjYASMgBEwAkYgmQT8JuVMZlurZgSMgBEwAkEQyCOWVgyceEZIWoSi7a5qGs1T6v66wNCIgW+9PNE9atjAz911JKoLBiPPSXmS3HlNw0YtnHvaa8DfQbiYdh07PTL191/HIZpoHULeEIpl7MhvBwcxrYBVMfQvmPPP3ynpK7p+o6bk4Vi26OwcCSQav//xLi9u3rBuzYjBX54VDinQfXgKHjEDkaOKJIfocFPrpk5De0lfThHyDLj7IKQQXg6J8UzJ/GijT/+XKV+xMuKF9nNN21v/y9z37Nq5gzwa/vq/tNVV12LQnT9r+lS9XrVmdF08IxbNmzXDXxsSsx8RsaFdh/898vpzTzywc/vWLf7qkVvhngceexrPi+++/uKspN7UZ4/wOkdyIaR07v7a1ZY1XyoiCHN3X8ebBIHtj1/H/tThoSee4bvU88XOD6vohLhFInDa9ez29CO7xPVE+0Bs4Hs3esQ3A4MZ75Vtbr5NwoZ9+4sY+99+qctjbnGncfOWrekP4SSYfqlbqWqNWitlcwdql9RaVqhStQZtySuCtwzfWXJTaH+IU7zHi+fTXm+85LxPw2YtLudzoD0dir6D/c2pHl2vAd/HQIJOsLytfvAEXMZ29UDg7wYVLhAd+PdLvSgw8PMZTzT+faIuAgH/RmneCK6nu1jhmr3ms+B3Rr1AEFMQGxAjECkomstCvUkQNBg74oQKGggdHLRTcQYB5JzfsOBXwFoYASNgBIyAETACRsAIGIHsS8A8LLLv2tvMjYARSGcCFcVISQx58lL8MOzrL5xGavdQrrz+pltJ/Dz484/fJ1SU+3rh4qeNxngwOK/hkUFy6cS8Gi6/ps3NhGcZPrDfx9qWBNbPv9HrE8LczJ7+1x+pRYOBkifiFyXh6RHoPggWyxcvnEcIIGedK65t+5+ixUuW+l5CaQUSe9x91qrToPHWTRvWYYQfMeSrz9xhZiTh+enwPMsWn5O7Q3MMzJ81Y1pqmbjbb954+gn3S8pWqOS8dt3Nt9855ddxoxkn3jIICM7rhHW66oabb18iYpMzxBHM2Cv+wjTRhqf6CxUpVnzdmpXLx3w/9OtA82krwhWiGntUvW+cdTGm89lpIE8tG74XCEsansvdn4Ypwnum/b0PPvb94K8+c+5x1ok9TViwSeN+GulsT74Y+neGVEtqvHg4kFh81NAB/fFc8OeJQt6IPbt2bF8vPJPqz3mdEE54r4gj0/zE9n+gtaQNPPDQaC2/E6LV5Pjk3de6OfvSkGLvvfL8U+7fDzxsEKN2bNtyVjgxbR+KvoP9zakhyeHx4AmGq9UNOQH1SMBojyihXhN4qCFQqBDAQDinIgDv1fuCaxqCKeQD9ncDh6eFhm+iGuIKogPeFBz67w51NMSVhrRyjh9xgvBRKt5P2GaSAAAgAElEQVTwynUVds5n+KvzwtduagSMgBEwAkbACBgBI2AE0oKACRZpQdH6MAJGwAgkgwBPVVMNQ/vXfT98J7EmbW5pfw9G0l9+HDHUXz364ulj55Pk1OMpc3IUJNZ305atr94rj+//M23KJIy8T/fo+f7Hg0aOm/33X5PJZ5GMqSRZBaO2N6RTSgWLAMbrG9vddS95FX4eOWxQkoPAciRjIEwSuT4i5EPf914/62lz+iCfADlE1OPB2S88EYWCNUonZ2wioqynXqmy5SpofYzFlavXqv3Td0MGqMdH8ZKXnJVbo0Xra9ogPDjD/NAewYKcCMeOHiXe+llH6bLlKyIicXLAJ++/pZ4J/saJKMT1cT8MPxNGyFmvbsOmzTGCL0hinyWHgdYpU6FSFcSZQIJF5eo1a1OXvCaICV993Kuns39NvD3g095vu++LUR8Pm2mTJ/6S3DEVLlasBOHW/v5j0oRAbRpf2qr1LPnOJLdPrcf64kFF/phAbRNbS8QXxM9li+bNaX/vA4/haeT8HUDQqyNrRO4Yt/jIXmcv/PXb+J/93TtUfQfzm0MSeBLEM79g2Vr9kBJQ47vms8DAj1DhDaknB94KGO/VI8HpWYG4oaGgnHkkQjrgZHSOCIMgwSueIhRC3iHIMBfGzWeEiLxSCkhh/HhWMD+8KjgHB67zGS4Urxe7hYVKxipYFSNgBIyAETACRsAIGAEj4CJggoVtCSNgBIxAOhHQp8SnTBw3OtDTzQyFsEdNJDn3tMkTxrk9DLhO2J96jZq2IL670/CMkQ9j5MLZiYdhImzUkvlzZ3V6omv38TOXbbzjvgcf7//B268+IQl7/YXjSQmeBk1btMKovXSh/wTKifWJwZL8AO5wUpK6oEAjCcODsEKy7OSMSyIBRWOox0D82fs9XxaN54C7HXXWrFi62F/iZJ76J+dIYgb+5IzDX53tWzdvhFHpshUq6vUbbrujAzkjZvw1eeJGX5goDVmlde6476EnEKvGjvp2iLPf6LqNGKvfEFy69xCqfht3dlJyZx88/V+3kRi7xXuDcEPucRcsVKQoRm+EkUD5L1LCI7puwya0CxSmKFrWgcTfza+45vrvBn3+KfPQ+7C+5JogxNX0KWcLDISOulS8h+jXmVQ8qTHivUDS7qm/Txjrry4eEiRznzVtStD5K6rVPJ2MnvwTgcaR2FoSQgwxpXipS8rkyp0nz8C+H5wlfra5tf09eNT8+O2gL93945nDuT/kN8jfvUPVdzC/OZJs3MsHD6uk1smupzsBDeekSasJ8USoJIz7CBcXSMEjDC8D/sbQvBWEWEIUQADQ5NXpPnjnDfG0kM8UxoPYQkGIYIzMB+9FnRueFJpQnG7Us4JzCBWIE4gWCBXqEcmcvd4lJlqc16W2mxsBI2AEjIARMAJGwAhkQgKWwyITLpoN2QgYgcxJgITWjDyxcDxcr1KjVh1EiUBPbzdo2rwV193GVIy6tE8sbwRCAKGmKM0vv+q6CWNGDe8nyaslQkzQCYkTW4WGTVtcTqJwf0/7J7V6tRs0buadh0t4qde4WQuerp859Y9JSfWh12vWOZ1wm5wX/nKBkN8AJn9ICCZ3n4RiKl+panVyGCT3fsHUw9Nmu8TmQWSiHaJKm1v+e/fPko8AIWOdZJjmPMZx7bdG7XoNG7e4/Eo8DCTvOk8Bew88LkjW7Wam13kin/fMJbFQWswXxnMltJK/ueCtwFP4gYSRYObvrMuaEyItkBAVXa9xU4z0hKga0v/j951tW1/X9hZCWI3+7puBbmHpsiuva4ug8fsvo0cFO7bEQkgRDor+Zv4dvGCB9xGhvPwJQslZy2hRK6lXVeImDR3wWR+3EHNTu7vvY41/Hz/mB/ecr77hlnZ4DAUK5xWKvoP9zeH3j3VcsSSwoBPsWlr94AmQdNtxsCSasJoLvMeTC1ECAz3eWxjvCZuEwR+Dvnou8KreCmcSUsu5853LwqOihe93Q0NEafgqPiM6kLOCv5eYE3NX8UJDXVGPZN0qWOjclZPfPFXBr4i1MAJGwAgYASNgBIyAETAC2YeAeVhkn7W2mRoBI3CeCRAKhif8p0/5/dfEhlK2YuWqXA9ksPtP+w73Y2BxGyTxBsCgu3Lp4oChZiR/dCn6Hjdq+JAbmkdX6P5kp3vSWqyIisqZs3aDJs1Snr+icVPGtHf3zh1OThjr+Tznn6lTkruUNevWb0TdLz569w1/hnrWxMf6nKe5a9Rp0Ign1Qmtk9z7BVtvy4Z1a2VJLiF0FbkWEB7II0I/6yThOq9OweKhp1985aRkDB8mhmrnvVTkWRggyTlGYOr/OmbUd4mNsZxv7wUK93TLnR29IcPSOlwPIZACCW0YvBFjEHQIleX0rmAsGOh59SdKXHPjrf/1XvNjvA92rZz1m7S4/CpCdgUSHRLrm+TviYWDSmot+Z7Tf5yoWm7xhnBd7BcECXd+G+6LBwXeFYFEq1D0HexvTuXq0XXE+Wi9U5BLzVpZ25QRwCvAUfh7ATFCH3TCWK8GeUIi4VXhzAnBTfFYIJzSYd81zRFBH+ddrHBS8QkXmhhcc28gwjBvBAjEGUQJXjVnBwKF5rPQ3BcIHHiZIN7oYXksUrYFrZURMAJGwAgYASNgBIxANiZggkU2XnybuhEwAulHgDBHxOif+vuv45IKu1RYjNaMTKLebHePkJA8ra5pc9Pff/w2nrA1zuskj167cvlScjwEmpk8pF6Qa+NHf/9tSoytySFWVzwhCC20aN6sGcmp765TW4zX/sJaXVKuotfTYOumjd7cD8k5SLhN+KRfR48a7q9+ZXlMnfPLFy84R7AgVFSga8m5d3LqbBK3AsQKcmy0vf3Ojogjmi8Dgy2hwyQndxX6IsxW8yuuvn7YgH4fkVjd2T/MqBso1FjVGrXrEjLJnXDcPcYLLy5YiHNbNp7rcYNnB0Zvrq9atuScBOXJma+/OnhH4NkRKJQZc6MdIbu++eLTD5x9FClWomSDZpddTg4Ht+BBOKhmLVtfQ/LmtNzriFgN5Z7/TJ38W0rmXKZ8pSob1q5aEahtUmupPNjThA9z9kM4KD5PHPvjCHf/V7a56TbOTU5EvAlF38H+5lQREZEQbSlha21CRkDzTmDUJ2wSYoR6S+BRgbcX4ZPIAYEgQaEOhns8FC6SgjFfE3NrIuuQDTgFHSOiMBeKHogtiC4IEvy7TEGc0UO9J7jO/BB1CBHF/Jg/fXp5iPhjoaFSsCjWxAgYASNgBIyAETACRiB7EjDBInuuu83aCBiBdCZQtWbtutzy7z8mjk/q1hLtyfu05nGJp+Su+78nu3YnZM/QLz/90H0No688le8NIxToKCDWQ66JI0ZAUSOp8SV1HU8B6iyaG7xggdAhwkvtBZJzwH0fwjchxoiTCoaxJA9yXuCtAvNAIg75GAi/JPbjpf54YghH8EjyZimssH7NacN1rboNGl9+dZubRo/4ZqCzqzUrli2uIMoJRvIuPXr2RnT4os87r7tvV7t+42aB8j8glOGh4M7v4G/IefLm9xrj9ri8WxBVurz0pjcUE3lVEMZSOOVzmjF35udvzb1sfB4Fs//+c7I7MXorYUbbyeN//sEdDqrpZa2vJnTanwESTKd0/JJjoT5M//nrj6AFC7xFEFI2rluzKtD9E1tL2laQxOy0dYc4I1QXYib7efKEn39099/yqutvxDtn5rQ//ebdCFXfwfzmMAZyg6Tl/krpOlu7swhggMc4r2GhMMpfKAUPA4zyeB6QhBoDP4IGYaKog1eFih2cp6iRP6N5HjAPDWOFaMFn9SxhnsyFVz3491mZOOdCO85rAm71wqBdmOWzsG+WETACRsAIGAEjYASMgBFImoAJFkkzshpGwAgYgVQT0JA8s6dP/SOpzvbu3u1NKHxxocJFnHUxrre75/6HZ4nh9p+p5xpLMUo7wyhhsNeQR9rPMXlsn/cqiiQ1lpRcxwuAJ/0TM8oG6rd6dL0GGMf9iR1iEQpDrOG6sz3n6jRscqm7Twkh1QAjbmKG5UriRUH4KQy57vZ4xezdvetMWCr68neflDDSNiowPdj5hZfj4xPix/84Ypizv9XypDlCzYOdn38Z0av36926HD927CwhiyTtVWvVrhdIIFKviNnT/0py72mSd9GNMM6dOe66/5GnyIMBJ8G1JikvoWCY1KrXqAkilCYZd7etL0niOTdh9Mhv3ddaXnVdW85JIvGR7mvNW1/ThnPTp/w2IZjxJFWX/BWIAsnh6e6rVJmy5TlHThV/90lqLes0aHIpAg0eIwslGbyzj5p16jfCA4v8I+68FsVKlCpdSdZvzoxpU3SN3fcPVd/B/OYUKV7SG7Juoyh5Sa2DXU83AmqM528GDYfEbzCfNbE2nxE7MfjjZaHJtjH875aiOSwYNF4IGf3vD+aBqM84EWbcOf+YF4IMXhUaCkvDXCHW0J42iBaIFxkqBFa67Ry7kREwAkbACBgBI2AEjIARSCGBjP4HQwqnZc2MgBEwAhmLAGIDYoI7hIu/Ua5Ycjo8EU9E63XEh54ffzn05MmTJ9584amH3O0wYoaHhYfnzpOXuNoe6n8xYtzkHu9+/IWzLnH3+axJmPUaIYm6vvpun0slEXdqyDW6tOUVeAQQsiol/dRr1KwFBnkSdrvbY+RlmsTp12uIFe/2GzSi/7djJnHN2aZ6dN0GfJ4zw3/OC4SP8pWrVnc/ta99cF15cq772336fznilymwTcnc/LVZs/x06BsSb4//acQwd9x+DY3T6cnnXsJAPvHnH84J9VOjTr2G5A1ZPH/OTH/3QJThvIS9mpvUuNeuOu05QbJqrQvvx57r8eaMP3//Fd5pGV6Je0gO6RaEwnJ7SHBNdJO8rCMeMu48FAhIkivlUhJ1+8t/UUe8TsjpsmLJovlJzTuY602at7qS8abE8+YiUSG5lzukl94/qbUkLBh1J4wZOdzNq658d7j2x69jf3LPB68NzgXaI1wLVd/B/OZInnvvd8stuASzPlY3JAT0txXxglBHe1kmKepVwTmM9HgHIkjwXr0x+IyAgYGf6xnNs8IJTL0sEBkQJRBf8LBD0HYKxeppoXXog+vkuaAt+1hzYCDyKIOMPPeQbBzr1AgYASNgBIyAETACRsAIpISA+4mhlPRhbYyAETACRiAJAng6LHA9ER2oCUZFDPYPd+n2Kk9DS5j6LQ89/cIr5SpUrtrlgbtvVQOgsz3x/SVP7drLr73hZvFu2HRVm5tvxxj/4H/btnbWk5QJK5cvXjiv44NPPLNj6+ZN8sD8sZZXX3/j9f9pd5dEoDpCUuPULCaeALRv2rL11W/3HTgckQEDt3gq7MQYHxsTEyM27xwYonPnlvgvBQpcICk7Sk6bPPEX5l2xarWaBw/s23fvw091bSWCTYebWnvzF3CMGTls0G333P/Qq70/G/jpu691P3rkyOEODz3xDCIHYZJg4Bw7hm6MyoGSipeRDNMY+v2F3qIfPETqN2ne8tGuL71BuK0rrm37nw/ffKlrWiYDJoE0YafIxTD8688/cbOXVBVeDw+M071efaGzv7Wp6AsRVL1W3fq9+g8Z2e6qptHisIDhzHuw90jAnByPF7xRENY6d3/jPYkOVSBnzpy5Ojz45DPcn7kP/PG3v1m/1OwRd9uKVavXFI1u9psfffnNnl07tn/wRvdntU5NSXyOcDTll3GjSVjvbIvIk1cs3ON+GDcajwd3v4WF6VbJxZGW3iCEmMLLZlC/Pu+lhAH7nXaILClZS03IPW7U8CHu9hp2jjw57mt8xzi3wReCzN+9Q9V3ML85sm0xhHtuveu+B/C6adLiiqvadbj/4a4PdWw3b9b0qSlhbm3ShIB6UvDdVw8JNcLjZYAhnr8pMNbjmYAhnzbqeeHMeaEeCGkysBB0oqKChnZCiMDLQoUYxs81RAtCYfEZ7xIeFmCeCBTMGzFHc3pomxAM17o0AkbACBgBI2AEjIARMAJGwAgYASNgBIxAkAQwqs7bdDD+2ptuuyO5TYnrP2Xxxr3zNx9KoPwyY+kGEv0m1r719TfdOnPt7hPU/23uqm2BvCXqSYid6St3HNG+py3fdui513t9THz95I4vUL3vJ/2zeOaaXce17+S8zlq35yRjp88nXnj1bdr8uWTTPn+8MKQ7+5yxaufR+x7p/Jy/8Yz4bcain/6ctzLQWDH001e3tz7s56+ORIQqP2n+mh3U+Wf1zmP3P/7Mi6nl46/9p9/8OKHPwBE/+7uG6ML9n3zxtXcC3btZqyuvpc6c9ftinu7R05tnwnkMHffnbLxDkjt2hBnWxLn3NC/JR19/P5a9mNy+klNv8JjJ/3Av1sodwqzTE127z92wP5a8Ee6++D7QjvH6u8/Y6YvX9fz4q6HJGUNy65B4nHsikiW3jbMegtu05VsP5pRkLf7aJ7aWiGt8b3t/Oeyc/BT09dXI8X+OmDjdbzL0G267owO/QZrA3X3vUPbNvYL5zUGQdH7H8Z6SvOwYjO1IRwLkWvAV8i5ESckr5UIpxaSUklJWSnlH4XNpKWWklPC9L+mrf5G8XiAlv5QIKfTpzeegJR2n5vdWzrH4xsY4dd7Mq7KvNJDXRlLqSKno48BnSrTvfA3feVgxd9jl8M3dO2c7jIARMAJGwAgYASNgBIyAETACRsAIGAEjcN4IEEbnljvv7UQIm2AGgdDRrGXrazCO0kdy2vIEOMKDOzySu+0FF11cEOMofePtkJy+k1NH58gr/ZJ/gdwa5SpWqVZN8iwQXghDM0+p80R4UYlZT9x+7Zuk201aXH5VYmMiFn+bW9vfQ8isxAyZhKYqXLR4icTGTX6HxO4VHhERUUgeT8egm5z5p6QOc3bn5XD24zbi+7sH4XwCzRXvGZJEBzM25txCckAgFDjnzliubntLu2D6Sqou48ag7W/Pcj9yRvjrg7XBAybQ94r1Z58ndf9grt/1v0eeGv/Pso3J/T66++b7QK6JxO4ZaC3h0/b2OzsG2vOEdStVplwFf33zHdPk5X5ZhrBvvV8wvzkIK/xGJPX9DWbtrG5wBFwGfIz3OaXk8QkPGOGL+kSJwvKKQKHG+eI+YaKAvPK+iM9gT/tcUiKlhLv6D25wIajtGo8KKogMzIM5Mg9EC0SJ2r7XavKKeFNTCgIGok0ZKRV8bGBCu3xS6Iu5W+LtEKyfdWkEjIARMAJGwAgYASOQtQgEZTzLWlO32RgBI2AEjIARMAJGIPkEECpy5sqZi3BkyW9lNY1A5iOAAd938LeCJtwm/BPvCXGEiI7YTEUNMUsoKA6+H4SH0pwVhFXSUFD0R/i+s9wMgtTz0xyoY77OeRP2iTky5zxSCP2kc0bE5vpO3/wRRwkDRWF+MICLvocHhzc81Pmeb5oDtA6NgBEwAkbACBgBI2AEjEAaErAcFmkI07oyAkbACBgBI2AEsi4B8mHEHolRo2zWnajNzAicSwBDu+amIE8FnykY8znP3xSIGAgRJJ3GQI+xXh+O4pVrGTIekltA8AkYjF/zbzBu5lvIz5yhxXXEDOZNLhbNfQEb/c2wB8Xsm2UEjIARMAJGwAgYASNgBJJBwASLZECyKkbACBgBI2AEjIARMAJGIBsSUJEB4z2Gd7wKnCKEihf8TaEeBSSgpj7eBgga9KFiRmbxMFBhRb1BNHE2ibSVg9NT5JCcR9xAsGDeHAd9HJzCTTbcQjZlI2AEjIARMAJGwAgYASMQHAETLILjZbWNgBEwAkbACBgBI2AEjEB2IqDeBYgPiBWEhuJQkQIDPgZ9rqmxXg3+Wof6tMd4z5EhPS1ci8oYVZxRAQbvCeZBSCjKcSlHfEyUD+IM7RAw1LsiM8w3O+1pm6sRMAJGwAgYASNgBIxABiZggkUGXhwbmhEwAkbACBgBI2AEjIARSG8CrhBJEiHJa2/HaI8HwVn5GHyfqYCQgREfg716YnBePQ80TFR6Tyc193MKDeplQm4ODsQZBAn1MiHHBXNnnsyfQhsVc7yNLH9FapbD2hoBI2AEjIARMAJGwAhkBwImWGSHVbY5GgEjYASMgBEwAkbACBiBlBPQZNnqIUFPGOI58CzAOM+BgR+vA4z3GO7J5aAhlLwVMoPB3jFGb0gsR1JuFW00hwefnR4VcEDIIJ+FJizXcFLKJ+WrYC2NgBEwAkbACBgBI2AEjEA2IGCCRTZYZJuiETACRsAIGAEjYASMgBFIBQH1NMAgr3kt+DsCjwoEC4p6GmhoKE3U7cz1kIohZIim6mUBA+arYoV6jygL59wRaSwkVIZYPhuEETACRsAIGAEjYASMQGYgYIJFZlglG6MRMAJGwAgYASNgBIyAETi/BDC6Y7DXXA0IE5poW70teNUwSFxzhkU6v6NPm7srA3rjvQoVzJP58hkGmTH8VdoQsl5SReCCCy+6+NDBA/udbj2p6jAdG+fIERVVsHCRoju2bdmcHrfNTKzy5S9wQaGixYrnzp0n7/FjR4/A6MTx48fSg5PdwwgYASNgBIxAZiSgieQy49htzEbACBgBI2AEjIARMAJGwAikA4HlO46EVS2a13unwyfjIuLiE8LzRkV4c1XkiAjjc0REeBj5KuJi4hIi5BxVvTkvxMPAGUrqnNHO33zIeY6G6pGg7/VvFv181vW6pQuElIAjJBT3cf795AyF5UzQ7fSoSMgMYbBCCtA6TxaByMgcOf5YtH73T8OHDHj/tReeTlajdK7U7a0P+2Fo9ze++x7p/Nx9jz79/GU1Sl8U6mFldFZRUTlztrqmzU33PvxU1zLlK1XJkzdvPicTBKn5s2dMGy1rPXbUt4Pj5Qg1M+vfCBgBI2AEjEBmImAeFplptWysRsAIGAEjYASMgBEwAkYgjQm4BAN373hUeE7ExOdYuOVwTjG+x4SFeXM0FIiKCD+eP1fE8ajI8IiTMfG5TsbGY5RLiE9IiBHx4rAIFwmxcQk5lm47EpsgqSDkM32pYU7fY+hXTwzOoYpo0m7CLlEQAPL4rh2WV/JiEI6JazG+8Qc0+KWxoOEUI9SzxMnMwj+l8f7MLt2VrVCpCk/ix5w6yb7OkMeV199068y/p/zub3D1mzRveeTQoYPpMfCMyiqvLGDHh598tl2HTo/gAQKLKRPHjZ4/a8a0g/v37UWowAslun6jpk1aXHFVvUbNWtx29/892Pn+O27eu2fXzvRgZ/cwAkbACBgBI5AZCJhgkRlWycZoBIyAETACRsAIGAEjYARCS0BDPPH3AWIA+Sk4hziA50RFscSXF3tbuMgHR+TChScT4pefOhq/JyHBU06u5xVR4gLahXnClovGsE/qF5C6UfK6R85rv7znKOzrFy+Mgr73uFrwdHY13+cD8kri7vVSCkmpLgWDKMIIAsU6KWukIKAwZs0twZi93h2+c75bpuwlEQ8JEydShtRa+SFQqVqNaE4vWTB3VkYEVLZi5aoXXlyw0PrVq+T7fe5Rs079RjOn+Rcz0no+GZFVm1vb39PlpZ7vS9SnvBPGjBweFxsbe2O7u+7t/mSne44eOYLQetYBS+rfcNsdHb4YMe6Pe268vLG/emnNzvozAkbACBgBI5AZCJhgkRlWycZoBIyAETACRsAIGAEjYATSmIB4JiBIYOzHowHPhqJS9vleEQ0QIvZLQSRoIOVCKQgEW8VS31zEi1MiEdwkn+tLWeCrU0+Ei+HyfpmU66QgOtC+rJQdvvbMpKKUYlI2SEHooO9fpNSQ0l7KPClzpNSRMlfKEilXS5kmpaSvPX1Th/YIHQgbGFN5Upmnm3k9KvPEE+KUeFqYwAB5OzIkgcrVa9VmYMsWz2e/Z7ijdr1GTRnUiiUL57sHV6pMuQoXXHRxwSXz58xMj4FnRFY33n7XvX/8Ovanvr3e7LF3984d/YaN/m3OjGlTAokQB/bt3fNS5wc77tu7e1eHB5945qlub7z35gtPPZQe/OweRsAIGAEjYAQyOgETLDL6Ctn4jIARMAJGwAgYASNgBIxAGhIQAz6hl/g7AEN/cSl7peDlcIXvfSt5RYTAqwGvB8paKTwljLDQXEpjKYgCiAeNfOcQQDiH0e0vKdf4ho2nQ6C/O5zXEE0uk5JbCsbRJr5xMca6UhgX90O8IGxOESmPSyGJBQXvDYy9U3ztJsurzm27zBvhJFaEC4sX71sYe8k4BKrWrF13357du3Zs3bIp44zq35HUrNuA77xn2aL5iIRnHXhXcGLxgvQRLDIiqwfbt22tUAgH1aBpi1a9Xn2+c1Jr2adnj+caN2915S13dPzf130/eGfr5o0Ir3YYASNgBIyAEcjWBEywyNbLb5M3AkbACBgBI2AEjIARyA4EfN4UCAqEesKzAVGgrJSaUo5JweCINwMGfoQKhAeEjeNSCLeEeMBnvDBoy3GtFI1Zj+ChMdi5rmIF9SIlz4U3vpSktfAGbpI8GJ54eY2PT4g8k0E77HQbqsgRI1WK+q5dIp9r+e7LPVv67oXwgJcFY8TDgjBTzKO8FMZTTwrhdch/gcixgbrCAk8Pb24M87rwsrYjAxCoWiO6bkYNBwWeGrXrNdi9c/s2ihtXdL1GTQiBtHzxQjyjQn5kdFbNW1/TJiIyMvKvSRPGJgWDhNt9e73xUp+BI35uc+sd93z+4duvJdXGrhsBI2AEjIARyOoETLDI6its8zMCRsAIGAEjYASMgBHItgR83hQIDnhG4FGRX0olKRjsMfgTN7+0FLwbEBww/iNWePNRSCGcEmGhykghdNQRKbulIA7kkoLAoQd9n3NIAm5P3qgIT6S8xolKgVgRLu9jYuM9kojbw3UKhyTsJsG3p0CuyIuof/BErOd4TBw6B/fi4N4qtjA2xBbECkQW5oSXBZ4geG6Q84Jxb5ayUkoVKcxpta/OQeGD4BFjXhf+Vs7OpReBYiVLXUJOg2WL5p3jvZBeY0jsPjlyREVVrFq91rTJEwnbdsbiZnMAACAASURBVM6B98Wq5UsXnTxxnN+PkB4ZnRWTv6z1tTesW71i2bYtmzYkB8b0Kb//evDA/n3NWra+xgSL5BCzOkbACBgBI5DVCZhgkdVX2OZnBIyAETACRsAIGAEjkG0I+AQK5ktuCjwLCKFE/omqvs84LXAOwyJCBGFedklBsMCDYpUUwirhOVFZCiIFIWrwyuBvB4z9nAuXjhBCED0OityAwMH9zjoQJ5AiYuPiPVEREZ6wiDBPDikRciG3eF3EiICBRwVCBQM7EZPgySPiRr6cEVGIGuHhnpMJRxPCj8fEI0KQTBvxAaEC0QVRgrEhViCcMHZybDCOUlIQNhAxmCNzRdjg3FYpDAuxY4WUOcKNc3wmwbjHBAzXQtrHkBKoXqsuIdj8hlsK6Y2T2XnFqtVqIlr48wCJisqZs2rN6Lo/DR/8VTK7S1W1jM4Kz4pmra68ZvR33wxM7kRjY2Ni5s38+69LL7/qunA58LpIblurZwSMgBEwAkYgKxIwwSIrrqrNyQgYASNgBIyAETACRiDLEBBjur+5YHA/7ZZw+hVDvJ7DG4EQShWkkDybUE8Y9xEVMIRhmCcUFMZ8jPiIG/mk0I5E2zMoIiAURIiQV2Kqz5X39cPCwvaJ1nAyMixsQ7wn4WIxq52Qz8ekzkl5j1BQVqQHnCOOSN160iZHpAgUuUWEEGcKz6nY+HknRHYQ0aIe50+KlwWV8+SIiJfPe3OEh1EtzudxcSpXZHhCvlyRB4/HnMJzggIMxonIQvgZvEFIVozAwriZN/kvmNMJKYwJMYYwUnhXIEwg2CDO0IYQUniZkKybPB2LaSfM0U8oCDsatUrPyal/DxE3zvpsH4xAsASqRdfxChZLFsybHWzb9KhfpUZtcsh4/CXVrlqrdj3EjMXplHA7o7OqXb9xs3z5C1ww46/fJwazNmvFReXya264uUixEiV3bNuCMGuHETACRsAIGIFsS8AEi2y79DZxI2AEjIARMAJGwAgYgUxIAEM7ng0IFORpwIiO9wECRFkpiBDUuVmKN22EFMIiIVTQhvpLfa/U5zz18FDAsH+UFBPi+ECeh1/lQiGpMCVWIjflj4qIzJcr4kIRGOblzRFeSepUwstCdIdK4gExVUSGmFw5wnOLKHFEruURr4mNEgLqcFREeN7cOcLzHDkZty82Ivwfie8Udzw2/kBYbFjMKfG8kA4SwsPCSkQlhG+Tdvtj4+OjTsSGHZS2xyQ8VMkjJ2NnMke51zLf/PAYySWf/5+964CTmvq6yZSdme2VXhZQeq+KooAiKIqIAiKIiooK2AALoCAqCoqISBcpIoKAWBABFRFRqvTe+7ILLNt3p+c7Z9jHF8LMNhYU/8mPx8wm77283LxkknvuPedwLmJDKiqCGafxN8EH0kb5joX1UPjOw2Ml9z6zNJh9IQTCaSvWp04GbfNdrk0IbhxFofYF+xc2IoDBPvQIaBhBX4rHArXqNWqSdPrUyeSzSbzuCrU0uunW23Oys7L8iWEXqqM8KjODQsGya9vllFV1Gzahvg3AjE3Ui/G7xFe5sVr5+Mo3rF6xfMmVjulKbHWl+y5Ie9I6OZ0Ox6Z1f64qSH1R5/TJE8f4PTo2rqQ/wOJanOfCjFevq1tAt4BuAd0CugWupgV0wOJqWlfvW7eAbgHdAroFdAvoFtAtoFtAt0A+FgiQQSFaiawJ0jDx2Z2OdAIP/KSTvQwKAQtmU9yDQgc9swsIUpzMrUehbNahY57ZFbVy+6DzPRWcTBS+pjZFuleSCQykAKA4hR2zfUqWRzqd7ZW8IRYp1WQ0NAdwUcNokELhv/RAbsKKem6LyRAB4CEEgAXkJwxhTo+SZTZIFnwmYVsJgBwWW5AhxuFWbkSbs2CDOqV4lXS722sAG5QXdRKRYZEIiqjdR867jyWnuBLDjFIjE8AQQAWnAWScwZiosWEEQEI9ilT8fZ7Hiv2nAXWIogwGSkruuMP5J+ujsB01PKi7wUwSZlkw84J/E4xgFgqBHgIZ1PMgLRSzM8jXz+0sBDsI/tD2tBvrM2vFw2wMXbwblrjKS2yJUqW9Xo/n/LmzzK75Ty0169Rv9HchHdw0QMeHez457MPx01LPJ59rVa8S5/NVWZg1cOzwwf1ZmRmXpXtRv4Lrjx7aT3q1y5bKN1avOXfZ6s2kjnrojma1mUlwJYMsqq2uZJ+FaUs6qK0b1/0FOQ/eawu8ZGVm8h4tWW3Bl1HrFed5vrFG7boH9uzcXuCB6RV1C+gW0C2gW0C3wD9gAR2w+AeMru9St4BuAd0CugX+OxYA5YlMoUxk/0eGgAMgOCQ0lPzFWMzkIc7GC+i+3du3ihfR/86RX70jiYiMik6H+iSjOa/eXvSedQtcFxags52ZAgQhGNHPjArqNdCxTkHpEiikcKITkc/1LVF8Ti8spHriQsAD7E0KnbykhKKjHdeWAg0KeR8us52oEUTwwONx/a3IhlKo6zzhkDYb3A7gF3KayxzmCjZKQccyPRk7s6RTZUOUMmVthjKlbIZybkUBRiGXUwxSRg7YnbxuZT3+ZlaGFxoUqCaXQvYEVvE4ZGsQEAizIkUBdCAtkxtUUXZkYmBMcjbqlOa2ctHWkL8PZ58sYVYOYL/HAExkZXt8GRSklZKxn2QAGGZkatgdiuQINshJIZC9CDVKhiizVAIoBfd3GvtogrtIJCmsYARSRbHwvkK7ksdJaHfQjlxPYIdgDxeCFLQl6aVYl7RYrM8sDwI5HA+zUgiKkEIqC6AFAQ19uQoW4G/t9G+W/bHs+wVzJ44eMfQq7OIf67Js+YqVIqKiY5C9UGg6KETjc+5KRwKABcVxUMEhIaFV4eRe9sM38/z1V7t+46a7tm7aGOg3OywiIpKUUcA00s6dSTx9JWO6EltdyX4L2pbnsXrteg3Hf/D2kIK2EfWEYDnnurZtcZ3n9p269nj74ymzmlWJs1I3o7Bj1OvrFtAtoFtAt4BugWtlAR2wuFaW1vejW0C3gG4B3QLXvQWq1qxTb+KXi5b99O38ORUq3VC1StXqNUuULlOOUYN5Hdzc6ZPHfTDs1RevewNcgwMAzmP+cc2Ow9/Nmz39o7cH9b8Gu9R3oVvg32YBOqvoUGeULR3odJaT2ogOdeotPI1SGoUi2Iz2Z1QzMyeYJcBnewIVjOyl89wA8IFZCKkyEAl0IeNvMjItlb2eMtB13eH0eteZPO5oryvbkX1q9zagB7udQWHS6pMpOSav021xZub8HNLQfS6mpguZFh6P4nWFm1znoGGx/a7S5qwWMQZLqkuKDIaKdpRJqlTaItlIDRVqNkRGBUlVbUb5BshQxFmNchMeAwCHBHj4IwBoODEiJwaFXUqHKbltkmQeqxxkkEPDQoMcA3bk7I82S940tyQfs0uuG4MlQ5hRNhzJwRHARkitcJ1zSa5yFsUIwMIdCoTiibLSz3FmUFMZJE+4ydd/KLpORl1mXqQByGB2BTU9LgA5FzInaFtqYdBmvJ+LCOfm+E5tC0au34nCzApS9tDp+hkKKXDYD0GldIAWzOTw2V7PuIAVinGpA9ohUgrt27VjazF2+6/oqlb9Rrw2pKIAFjMmjBm56ueffjh+5NCBq3UwdRs2vdlgNBr37ty2RbsPOugJIiz/fqFfMIP1t/29fk2HFvVvTEs5nwzMIvVKxnkltrqS/Ra0bZPmt7Ui4PD32tW/F7SNqGe12Xz3HafDzuyuS5biOs/tH+z2KDNcdLCisGdHr69bQLeAbgHdAtfaAjpgca0tru9Pt4BuAd0CugWuSwswg2LoB59+FhNXslS3Xs++cGDPru3bNm1Ye/rU8WOkp2DkILMpyFvscbvdHvBW8EAZcbhn+5ZN1+VB/wODJs81xSpdsOM/sHt9l7oF/ikL0OnNSH1mUrCQlkhoUpD+iA51AhXMkGiWO0gKRJMOihkX/BQZFaQpYmbAedyAcB15d8uKEq143RUNruwzktezFQDBFsmeflRxuzO854+fNDhSEm1eZ1a2U0nedyohAtkMcpqlolIx57hS2p5gtYc1d2XlZFmyjCG+rCe7kxoaijTzqNM486hvX7zfsWQFGSSj0ys5Q02yt1GUcd1jFc3lWsSaWtmM0okwk1zjUKbnB+RtZOGALZFmOZ7i3HaPdP68S7HGBMnhSMDI+TvFc2DsQafzpEOyoBBUIEVT0IFs3365H46D7zE+cAd1+B32UzznjkqJpSySfFOEZK4VIm8DiGJmByWDpJKofA5IUDr2yf6a4W8CEeSNJ6hD4W7ed6gPwiwL9ikyLlifhYDEDbmFdXqgELjgOKqhHEWh5sUJgBd0OrJ4dfACVrjC5aYWrduwi80b1qy+wq7+dc1r1WuITCBF2e1HHyK/wbLdlVIs5bePBk1vvpV19u/ZuU1bl2Pnup1bA+tXcPvJY0d4v7ri5UpsdcU7L0AHzW65/Y6c7Oys3du2/F2A6pdUYYYuV0COhPR8lyzFcZ4ZENLopltu/27eF58Xdmx6fd0CugV0C+gW0C1wrS2gAxbX2uL6/nQL6BbQLaBb4Lq0QJnyFeOrVK1Ri6KInds0q6NTPF2d03hjjVoUzM3X+XF19q73qlvg6lggD40KAVQIbQrSPFFfgpRDBCd6oRxGoaOQWRZ0hgvAgvRQzLCg45xZAHS009FF+idmU5yWPa5EgyNjhdfjskkma2nT8XU7pbMHMnPK33LadnR1qCX7bFbcwRVZ6ZIlWJGVbCmohCPEXMoWJJu9h6Jbu61ee1iYO8N4x7kV5+aU605ARRSOl3QiBA+4X2YlMCvEALCCn7ZMt+JZddbt7BUf5AZ4UYli2kjtOPHxAefOL487OU72tQkZGEAfFBNAC0OISc4GYuE5bfdakSHBfoR+BzEHsZ9cSquL2zkWbvNpSiATQzlmV0wHs6Wc0hYlu4oNuSQQDO8QJ/8eY5aCLQYpCKDKdmRc/AyNjVuwA2p1EIzg/gj8sJD6ieMTehfMXuF22lwsf+EL6bhIGUWwozLKRygEORqhkKffJxKO808Qicfgl+YOgIaqW/2rPwvcUK1G7YSTx4+mJJ9jNlGBFka6MzOAQQT+GlygbzSbBRVPfp1aEAIPOYY6dEgXBiRgFqbL5XQGokyiBsSxQwf2MfAhvzGot5NmqXqdeg13bN64Lr92PFbIf+ASLDzVYv0mFwCLg3t38/5zyVKrbsPGXLFjy9/rA42B2TF7tm/dVJCo/qtlK+3YrsQeedm6MTIstm1av6Ygx6rtJzrmAr2XljYrv/NM+tEq1WrWNqMiztEOBs74G2OFSlVupH3zA5fym0v/5u1X67z+m49ZH5tuAd0CugX+qxbgg7i+6BbQLaBbQLeAbgHdAvlYYP/uHdv4Arpx7R8rdbDi6k0X0m6x99079KyUq2dlved/gQUEUEGwgVH+BOroFGdWRVcUghIU1KaOArMtWqMwkpnUQ2IhldFpgBM7UDIkxYuiHEfZI3ldK2RX9u+GzKTl5kMrNwTv+GaXZfvCZdZtCzYFb557Jmxx/5TgTbO8ht1LS7jtWVWMzozSkjOnRpWU7TcDoDDbjbYIu9Eadspa1mYBaHFD1iFbSUeSF9tsIe4s0pYIMWsBIohsB64X332USxWCDTcAsLgj3CzfDy0KyykIUGCh859trTkeJRhgBf/2ZrkVI8AKrjfZvT5AhCCNELoW/ar794EkuQbheman8NOY7JKsOzMl4/dnFeOGdEV5/aA36ZUD3qPvHlH2LT6r7EG2xlrsdw6AlFVAEX5Dmx9QVqD8ikIA6DgKs0dYdvhsfYE+Siw8FzwnPDc8RzxXPGc8dzyHPJc8pzy3PMc81xzrZfz0qj7/1V8JALwD/vva9RuRmizggkBx2uKShcDBa++M/vS2O9vdq95wx90dOo2e+uU3zFxUr+e+Xnlr1NgJsxct/fjzud81veX21laoEY+eMnshy8iJM+Y90efl1/wNgjpIzIj8c09C+pp9pzOfev4Vv3oCb44aN/Wz+UtWij4YlPDBpFnzv17+11YKWVOXSmy7+bbWdy3fuPfk7MUr1y9csX7n/F/WbqcDOC873Nm+40Osu/7QWfuvmw8m1mvcjBRjl9mlRu36DdUOfzqou/R8us/bYybPfPjx3v38aRqwE2774vsVa6vVqkuKM7/LDXBkT5zz3fL1B87krNx+9ByPI1BdgjedHnn8adZf8Ou6HSPGTfuS2gl1GjRpRlHv5LNJpEO7ZKlVv2GTpNOnTgbSpqgBQIVj7PLYU33+SVuJfRfGHoW9GJmByyzRotBBcV+cTwTPIOHFjK+LS17nuVTZchU4F+f/vGbbnCWrNnKOtrijbXvRuA7AsPFffPPTJzPmL+Z85/oOnbs/zmvow8lfLBg+ZtIMzvv8jpXXLfv4dNbCJTdWr0UtIL9LydJly/Eeob42CCLwWuW1BUHydtqGPCefL1y6avqi5asnf/X9LxO+/HYZxzxu5oIfx07/+ocx0776lvcIzkfa2N+OC3JeizK2/Oyib9ctoFtAt4BugatnAT3D4urZVu9Zt4BuAd0CugX+QxaohPBOUhVt2bD2z//QYf3rDgVilQ1IsZV46iSdhfqiW+C/ZgGRMUDHOh3YFJ6mc7cqCh3bdIDfhuKjv8ldSPkkljsu6GVLiBhXgqBLcRAi2TsBVpSUvO4E2eveCsqndEPO+ROG9MQcJfVkomXb18nGzDOpwY50o10xWNIVk2L1ptbPMtjkbHNweZdsTo1ypZyClrXdYbBUrJGxt4LNk+O84+yKzChXqqG0PTHqWHAFl0c2psQ4kyWnIciEIrkMyE+4cAy+jIrcT46Tf/soopDNYIkwSfGoyGM0pbuUowezvIx2JyjBesw44N+kTuJ3ZmoQ0WB72orvKgIgUTv6BU2UEND2gRS57XzgR25bfneccV7Q8zjvkkyHcxTvujTJWTdUya4aLB+oh5FVsslyRav0G+ioqAdCJzWzJZjh0oDtUJhxQacesy84Xu4P58Infs4illdV33ksFFHenjs2ZmdQP4PZHOJ4/WZcqPr4V30lUHHvQ916fj1r6oRAA3v3k89mQ+Kpevf2t/uogsRCxykdr6XKlC3/x6/LfuR6OuUHjfjI1xeBi3Nnkk7/8uO3C/g3+fxr1K3fiFSLdNhTKwEJFodLl6tQkZHkzBQ4l5R0mYBzCexg2oKffo8tUar04oVzZhEMeG7gkLeXfDvvS2ZIqsdUs26DxvAPU3NEur3NPR0+mDxrvgJhF/4E3d/10V6Lvpr5GYEEjuWdsVNmMVNjysfvDyew3qrtvR1ff/ej8X26d2zrzxbP9h/01jMvDxrG9rM/Gz/mgYd7Pjngzfc+6nn/HczIubhUQcqGLTg4RAAWdMiO/2LhT/wt5DHe1/mRx8Ijo6Onjh35tnY/Z5ISfQBauQrxlfft2n6Ztkfjm1u0pIOZWSlfTZ/0yV33deo6+P2xk+67pW4VbV8xsSVKEhiiTf5c+ctSamK0u/+hbtVq1anP8W3Z6P/ZhxRNpMcMNB/OJF4YY/mKlS/bp2hzLWzFfRXGHkW58EC3xHu3tGndn6uK0r5i5RuqHj6wj1lZlyx5nefX3/loPNvNmzHlU86XLj2f6jNywsx5LetUjGFWD8EsAm/JuLhwiksx8IaZQuUqVqpCEDEH9FPAqXg/9rsQxBry/seTOmL+igo54Kx69bnHuvhrwPsDy95d27bMmTZxLK/d98ZNm4O556vfqt29He+5qXb82aTTF8FfXHJejj0Mz9hMveN8ZTYQKbJCw8MjwMgaRVCFx+Avc6Wg57UoYyvKedTb6BbQLaBbQLdA8VhAByyKx456L7oFdAvoFtAt8B+3QN1GTX1OBopH/scP9R89vOq16jb4L9IVqFg46HSlk/KSKGu8019Xjst/dJJcvzvnOSdQQYc4neEUeeZnCsqjKBR1VlPX/I1sCT6rh2C23IjvnDpbJK8XWRUelyQDf/A4QaRkdMO3s9OUcvSIJXHHTnvFW5ravQZ3TvLpw2Fb5nq85w/GZBltBpOHGhfe2llBIbLbY0zONoXscckmAA5yiVRz5EkCF0FeR4lwd3psnPOcqVnKhlLp5nDbSVtZ+bw52lU567DHrLgMiZZSMrQsnNlSsAmgBQELghUiY0TMawIG7jiLwXAkW9lWKUQ65laUlK2png0pToVtuF1kRvDTd3AodPLTBsyuoG1ERgKd/OybwIOgohL2FKAJ23Mb11Mcm3+LTBABfghQQ9meKbm3ZyrSn6mSbDYoyoMl5KR7YuTsUJNUB5Vz0HgZPqkfQqCCYAOjnpltcRSF+2S0OfUsuFDwmNkgHLuPIgcLo+npwGTGBiP8CWwQuGE/pP5JRxHARW6Tf/dH01tb3kHh5N3b/fPzt7n3gc7tO3Xt8e3cWdO0R0LAgus2r7+gQUFH96vDR32ycvmP3xGkYPR0y7va3y8AC9Iu9erUtgXrNgAlEQGFD4e9+qIAO/xZis7Vjz6bsygantleD7ZtQZFoRoMzAp3AhRqwIABCJ+jMiR+PImXR6KmzFx7Ys3vHwN7dHyT1VFRMbJygn2p++51tCSQMfv7J7ku/W/AV990HIIjL5eZ8u2whyECwYsHsaZPeHzKgL52x2ZkZGVxH56o6Al88W+zcunE9M1Mmz/3+l7iSpcu88Hjnezev/+uPb37buLvrY0/39QdYuOGQ5s4PHdh7mZO7DFAM2uLE0UMHn+7SvhWj9nFcx157+8NxdABD+5r3Hd9ChzZBHh4zARVxfnv1GzDo+deGvcc6OzZvuIx2iuAQgaFdeehX5DVG9nutbFUYexT1KqQ+BOmYiqJfQRCBAN2SRV9/qd1/IBsyk+j2NnffR2Bt1NBXfBlKBEvufqBLd4IV/Hvhl9OnsPD7lLk//ErR854dWt9UkGPk9cTMBu5jw5+/rxj99uD+zMBpC+Cr76tvvjvhg3fe0Pajvc67P9XnJYIVBPqCLFYrMy1ubX3XPep7xGHM36c639My0JiGvPfxpPjKN1br/9QjD/D+o65XmPNalLEVxE56Hd0CugV0C+gWuDoW0AGLq2NXvVfdAroFdAvoFviPWaAuHBp8wT96aD8jcPXlKliA1AaR0TGxu7dvLrRY5VUYztXqUoAVwlkrHLVXa396v/+wBaBfoNapIGBBKiEKZJNWoyLK7Sg+jngsqSh0YlsAUMAproBqSD4Cf+ffkseZrnjcO2W33WTwuDPclrDMoJQjJqPbfsZuCDrtyTxnysxMVcwn/t6ZcnT7WdOpzdHW7JOVnLKxYo4c5EIwrREAQ3C2MZiOdYvFY7caDSbJLSNc3eu8E9kWRxOsZfbZjZZDJR1nYpBFEZNhDHXkGG3OU7ZynsrZh0uYvW65hONMlkc2GU/YynnRnwAexDEKnQbObw/+MEWZ5arQjKhikuTMMjZDZWQxUNvB50zDwncRthGF7QhaEBAQgIOPQwqLAC+EODm3C7CCQAbr0YHM9szKIHjAwm1C50KMl+eBdpYTL4xEmZOoKKtSlPQ3Kxk2QqA7AY0cGCu37sbBkYaEfQuAhqATMycIOkXmjo16FidQqLFADnnug9kxBKL4nVHXjPBnO46LffuAHcyR60LfotFNt95OQJkR0T6rqRZGa/cZ+MY7XEUHqnZ7dQAGXEeAgnVJT7N/z67trz33eFc6V/u9NmwEMAFmsFy20JHLlQjazvO3oeezLwxkFgijvwlWsA2zI/jpQXqEuuMm0Bog9z8zB0ZOmDF3/+6d23p3bd9aUD6qtTLKlq/IcyupM/8mjh4x1N9Y+Ts26N0xE7ZuXPfXyDdfeV5oRiz44vNJpHoS4xJtCZaQBoi2IJVOuQqVKgNsuW3Pjq2bWOcA1tPBS2ev02HnnL241KhTv1EWhC+of6Edyxujxk2hw/nlJ7t1FBRDMIVfWwwaMWZCPLJi+vZ4oJ0ajPp+3uzpArDg8Wj3wWyMC+dlMzOJ/C4co6/O1k2X1bmWtiqMPQIdS37rGzRt3mLvjm2bA2lI5NWedGGcH/7opAKd5zLlK8Rr5+WKpT8sYvG3r+p16jf8efGi+fkdh9j++rujxxOsIODx/pD+fXjdZ2akpRHYIoDoD7BAZlDDxISTJzh/eX77DHzznXkzp46fPOb9t0qXK1+RgAUBuYKOgVkRDz365LPjRr41aLufTJ7CnNfiHltBj0Gvp1tAt4BuAd0CRbOADlgUzW56K90CugV0C+gW+B+zAEUx6agpimDl/5ipiny4Nes08Dk2AkXvFrnjf2dDQQ1EZ6qeXfHvPEdXNKpcoILnmVH9jKync5uFUfeMHCeXPB3Z6gUObh/lE3SilRyIZp8ExdNer9edJOWkuUEBVcmYkyKbnOnJSlB4TvDJ9SHBSbsSzpRpkuPJSVccRzdFmVMPx8W43RDvVuzJ5ig6xQ1u2WgAyHDqmK1CaqQrLRaZFRWjXSkVrR6H0yu7ykP22mZQvFIJZ1II5CTOhXqy4kAL5QZVVPb+0BsTStoTjeXtJ4NBC+VZH9UMoIqiINtCMXtdBC24DzryxZwWYtmmKiGGsOphhvtlWbJipSnVpaRAx0LMeSHYTQBCABjsh/Qk6mwKOsd9jlYsdDrzehGi3wIYEFoWQidCUEQJjQ22FdkZrMvCRVx7jrOgjUIx9Nvndb5QXj5aIki2giYqEWCLBYM5YsB/+MfzRUCEFF50utGJy3Wlc8dE8ILnWPQvzi0BKRY6nH9GYZbBHyjMthCZG8Iul9wPKNj+bxDlpnOfwP3cGZM/FQel/rwb9EHk76fek78sueq16zY4dvjg/pPHjhx6qEevZ8g53+3uFg1FJDjVr/31y3W16zduyuwIfxoKog2jzXv1HTDoL9AZiSwNbqsGaiV+wvFPHZKLC8EX0kExeyIEKQbM5gikTyUc/nTA+ki+8lheHvLuh8AWbIh4f560NqIq6Ww+HTV8sLYpo753w7nbonXbfbWJaAAAIABJREFU9nd37PzIsP7PPSHACtYl/RVtpAUruI1gx84tf1/2XHJTi1ZtqFXxyXtDXzt14tgRsc9qOAfMHlEfJ+3ArJhVv/z0w5pVK5arx5eRKwJOKqztmy+nfaJ+BZ+J8JvtA1f8LXUaNvUBMgRetNuvla0KY4+8z27grWAziuScnj3104+K0gcpxmjLDX+uoo7OJUug85yWckHrwjcv81moKcHMmoIItLMr0rU92P2J3ku+mTf7vcEvP8exUYvi7o5dHuH2Nb//uky7SwIZ1In4Zs4Mn1bGS4PfHnU++eyZsSPe9FHlEUDLb5zq7cyOGvLe2EnrVq/8hZlQ2raFOa/FPbbCHIdeV7eAbgHdAroFimYBHbAomt30VroFdAvoFtAt8D9kAdI0kDrid0SG/g8d9jU/VBFFu3Nr4GjNaz6oq7NDOiSFI0sHK66Ojf8NvdJpTWc2BZnprOa5DkWh05KO9nMopAmiXovP4YQKTvx3CtkU6xW3I0t2ZFX0uOzJkis7Pfj8AdljCrHaUg6lhh1ddTAt6sYU26lNJtmeYo849JcN+hTRBtlY1S0ZLQASrFmmkGMAIZyp5ohkZEaYoE8Ri8yJKqHuzLLImnCD1slkk3LcFq8jEtkUdkWWY+wGqwSdingMJcgtm7Z4ZYOnUvbRZqXsSccgvu1ABoZi9dgdRsWTjL5dVq/dBcCCx0LQQeuMMraMM8WaDFIIHP1GIDDZa5M9R5xQucYiMh5EhoUQ6+bf6uwjoUXBddwPrxuCGwQwCByIdxmRkcEsCO7AJ+idW19kMQnKKPYpQBFB6UNaK98pSHBIQa8fVFyRJsV1c4S8pz0gpHibbIEex9lgIzJjFMkL8ILC0SVRqEnBjBn2SdooUgYSnCIdFPVJOC4u4hzznFOwmoAVwRdSthOcoTYSszMIaFySCZDb/h//qAytBVIH+XM805HZ+6XXfRkHgjJJPWBmB1SqUrX6IlBFBQVZLE8+P3AIo64P7L0AIjCyHK7OUv4iqLm9YbPmt0E/ykclFWh5ECAIf6snjn73YuYDaXZ69n5+AKmV6KhXtyVQwGhxcv6/89oLvSkcHajvDX+tWkGHbYs72rX3d3yiHZ8TSIu1eOFXs7SZFP76pi4W9bG+hi1eGT5q7Kpfli7+YcGcmeq6ZStWqkw9CW17ZqkQyJkzbfzH2m09n31xIEWy50LXQGxjBsWdd9//4OfjR/sonsTS+6XXhjJy/pP3hr2u7QdsT5zDEgEVyBZwrl6y1KzbsDHHhiQPUpz5XeqBTnMXKMS02gPX0laFsUdecyyvbaT2ol5DUWhDOf8J+HGeqrUduL+8zjPnNAHAW1q1uZv7ziugpmGzC/oa2zblT2vKYyFdG3VV3hrY90nRLwE1kW1EiiitPajtwnUb16xeSfCmzb2dugx4unsnAlZcX7psed/vnJbWyZ9deS1/CGFwXqNDXniqh79jK8x5Lc6xFXWO6O10C+gW0C2gW6BwFhAvBIVrpdfWLaBbQLeAbgHdAv9DFuBLOaNL/4vaCv+m01irXqMmdBrlFUVbHONlRKmgsiiO/grSB3wJkqbAPyyz+Nbry3/LArnZFXRkC3oiCmrToU2HDumg6DynA5aCv3T2IfGAHEreaQAqfpbsGdsMmWfOSGknU13ZqTusSTsdhqzzMU6nPcOYtMeQk5kSfTg14/wep8V7yBNqBhFUebtkLJtjsJ4C5VMyAIh4ryTfbDdYqsEfHguAIgbAxA3ImGiKbIrwTFPo2SRLyYQzlhIZADYIargAaKAEuexGayZACHtyUHQ6hLhLgi6qrEHyxiRYyzqSg2KyQzyZYejLGuc4Gwq9izBsJwjD41SDbz6tlvhgQzholXxZJHaPcmhpouus0+sDHARVk3DO01Yi08In2I3CPkTGBLsgyEBggXVFNoegjxJ/81P0LWim1LRrBJHYD4ugkyLowX7YN79zvSXVLclLkxVvv32Kc8QRJWtGgnIeGRgnXYpkB+aShDqkfmIbfidVEcELgg78vhRF0CJxPDzHPNc85xwP5wDnAucE54YAYMSx8Xj/VYu4Z2ozFTjI+7v0eIIR3Py+esXyJdqBwydfm45XRul36NL9cQAfYWpNBiEAfOLo4YPatuSoZ9Q2AAuCOgGXDp27P87ocZGhRyqo0XB4Unti5BsD+6kb8vecY6L+wuGD+/ZoQQLtTkhxwyjv1u3ufYCR2oEGQVFxOo4hgDy+ICevVv1GTVifmQ/RMXElRr454JJxBiP1gw5i0lVdbtOatbl9q0ZXi7oSzW5teSc1AoSjmH1MmL1o6bEjB/fPnDT2A9EXI9ib3nJ7awIyR2AH7T4o/M11gUSkITnVOK+MSB4bswP8OfGvla0KY4+CnLNAdeo3uekWbisKYHHXfQ90oabK9/O/nFHQ8yzqfTvvi895fbS4o237vMbfEHRV56EmzyynvOoRfHxj5CdT7HZ7zuB+vR4RQBOv394vvvYm2xI8ECLx6r6q1axTn39v37x+7VMvDByyZcOa1b//vOR7UacidCj4nboq+dl66Afjp2HaVnm9b69uHLe2fmHPa3GOLb+x69t1C+gW0C2gW6B4LKADFsVjR70X3QK6BXQLXJcWYMQdox2vx8HT0RAdG1fiWoyddFDcjw5YBLY23l8Z3ccC+VrFlPsp1hXoNOFdt9HVtnHHh3s+SXFROm8KNKhCVKKDTDjtCtFMr/ofsQBBChQDygWhbEmi86YjCh3SpDvridIm93BJIURdhBPwXhOs+NLj9XwLQGKL3ZHzd7rDpWSnnU3NOndyX1JyUnL2ueMhmSd3Ss79K09kndpx2pF6OiY2YWMlqyOtssHrikXWQxQyIxqVtJ9pFObOaIbMiDhQNoUDjEjG95AQT1ZlZENEeGSDE2BEDsS1Q8yK04YsCmYtZFq9Di/WmcyK223yuiLRX4WSjqRbAUxUwXZjsCe7NECLoDRTRAqyN6Qy9gQr9mPAehOyLejg5zELGiYfPVOIUZZLWgF4GORSOD673Ssl53gu0jkJCie+iwhhbKHvQrBCZFwIAELQQBFoUGdhEJQQ+hnsk2MhQCL0LlhfUFQJKig1dZUawOB3AbpcQjG1Nk1RvkpUnAMPeDOWnFNOnHNJPyFjZDkqUzuA4tmHUehQZyYFsyTWoqxH+QaFIroELQhm8Jzz3HPhXOCc4NzgHOFc4Zzh3BHH+K9BM6tUq1GL1ETHj14a7U+al6eef4Wi4hIFfSmgm3t8Fz+q1arrc2Tu2b51U/en+r5Mp7la9Jl9czvBA21b4Qim81O7TfxNbvyKlW+oKgSL6YT/evmarU2at2g14OlHOolMDlG/fHzlG5h9wb+nj//o/YJQPXLMbPPIk8+96G8cjJJv17FzN9I5qSmdAo2Z6+vUv/BsUa9h05s5DrVGBtffAECBTn/SbGn7YRQ8x63NSmnWouWdBGRoCzqfSevz9c9rtrJ9n+4PtKWYueirVbv7HuD3H7+ZO9vfOCl2zvX+AAsCSXSy56U5VREUYaQh0jrxr6WtCmOPvM5VftvqNWrWHAkPh0n9lV9d9XZeP8/2H/zWmcSEU0u/vSDorl4CnWdRZ+HszydTx+SJPv0vy5BR98PriHot+Y2t2xPPPE8giwL3PB5R/8FHnujN64Y0aqQZ47Wu7YvXudB+ufOejg9Rd0Jdp0q16gGvc3W9hzEGCnVP/GjE0EBgWWHPa3GNLT/76dt1C+gW0C2gW6D4LKBTQhWfLfWedAvoFtAtcF1ZAO+alRf8snZ73x6d2iG67rfrafB8gZ/+zbI/ln2/YG4g4cviPB5SR5A/21+UV3Hu53rsC/4SDls4BIVTUTj7LkY6o55PVDZQNgEjQOn8yEu8szjsI0CuI1dBPP21tz8cVwFOsycfbOejXtCX/x0L5GZU0FFODQNGzdPpTId0DxTSYVT3Y41GuGB+ULzeFIeibLE73QaX0+5IOX8myQox7aDE7bIxPdFrDC1ZMjUr6XjMma1nLV6XS/E4bNCyqBrpSglDBkQYsh4SoC0Rh8yJaJTGyHjIAd3ToVBPZkzlrCMt3AaTAl0KQ47RmuEwWnNA5WSCjkVZABpYZ0slABHhSfOeDYq1BXnTalu8Thu2ZQHocJ+2lCEVjTvSlVpiXVSzY9vC66U0S9kQd2PWQWRclDkV5Uo1pZojcwCCQCcDuRQXqJF8AVEuRfFEmuVoo+yziYRPG6iUBLDBVQJU4He2JbjAdbyPqGmRCEKoRblZl/0InQvRl8ikUIMUoj8BjIh9qYEA0ZfQx2Ad9iWyO0SAl+dgtuT68Jji/eGscv7hUvL51lGyARoXjLjn+aYzkHOAQDqdeRRq/jb3mAhqUNuiAzvPXUi346PcwcKMCzrQCW4Q8KBTOTm3HzvmlwBzxNhU3UjXROOCFD4njx45RD0D9c6ZMREdG1vi3JnE08Aqdvhz/letUbsuo/2ZSUGtiXkaHQzSTbFPf5kE1EAg5dDBfbt3XnLQqj8E3U0OeIs+x7MBo8kP7Nm5vXv7lk0OQc1a2450NVxH5/IvS75bEKhf9XpS4JCyp+tjvfvOmDBmpJYiqcktt7UmxVNhRI1FMMSZpNMJX/jRPqDdLtjFD2DRoMlNPDYtHRNtweOiZsgnM+cv5m8rNT3eff3FZ9QgEfttfvsdbXk+Vy5bzHl62XLTba3akC7KX9YAhKB9Iup7IDIdyH51MUZu09IQXUtbFcYeBZkH/uoQIGKG6B+/Ll1c2D669Xr2BV4XpCXT0maxL9rQ33kW++E5nTNtwlhSshFg8gdK8NmKYMOCL6ZNymt8zEZ6tv+Q4Tyn6qwjzuvnBgwezmuKIJg/ijL2e2ONWnX3gT+s2xPPPs+MJC2YxuucQIcWmFOPqVa9hk36vzliNLVoCOLldc0XdJ4X19gKe271+roFdAvoFtAtcGUW0DMsrsx+emvdAroFdAtctxa4q8ODXY1488DLxWWRe//2gyLFAF++9u3a4YsavNoLAYsdWzYyWlZfci1AoIIZFfhTRC2ro6TpXOR6UsWwCAdiwOcOUmOw66sNWNDR9NAdzWo/0/W+O4rzZDJTidzl+6/RnCzOset9XZkFmFWBHuhsphDzPSh0SpP64mGUiigEK8iPT0ogH5c3F3ig58MXuAs0UMlwVJV0Z6eGhCcfqFg6YV2E9fTWEFvWmbKhBq9DTj582nn+pNHiSK9WNuv4rTZ3djnQN6WctpY+l2kK2Q+QAjiAUpKAgcNo8QKEkEHtZAY1VDY+nQAzjEbJA2e5HB3izopHtkUcwIhgbLMgBSo+wxRaDqUkuclAFZV03Fb+j/2hVdfuDq255VBI5ZNob3AZTHKL5NUN+x2ZcFv99K01IMgdWSn7SHSF7OPMxrAS9FAt/MODzAqvxXhRj0Jye6VU6FcIZzfvEfzOuqSIYlaFCKQSwIG4t/BTZG9wN+JeIwAPNeWT2Cb65ycX9s9sEu6L69Ri9yJDg5+CYkrsT2hziMwOX2f7siXP8MOK5/ZNvgMnFRTPL8fJ9oLPH+oXvnET0KA4LjMPFuaOhx8EJjgfElE4RzhXuqNQ34KZF91QGOHO7AQ69KmFQgcw75Xsk/0TDCqHORiHYkMJzs3yYbaPJIpqn0X+Sse3NruCkfLMrlj45YwpdIru2Lxhnb8dVK1Zu97hA/t2kwZo9mfjx2id/ZC38GVvHDlweYYFhb7p+MwrC6J+4wt0PMPHTJpBqhgKVz8MQW9/YAXrMXOBnz8hC0ELwORloM8/Hf0exZXv7/poL2090DD5flPW/7ny14Iamc8WrDtp9Iihgr5J3ZZ249/Aai57TqvXuFnzrRvXUfT9koW2iIktUfLdTz6bTYrFpzrf0/LV5x7rogUrhB327Ny22Z8+BZ3LLMyY8R9NX6c+z0leWh0cIxJy9lFPQz3Ia2mrwtijoOdNW68KADDSc4HyzO/8D9Qvo/77vTZ0BGm1vgO1k796gc6zuu5Xn0/6hJkzPXr36++vD15DXL/178vni7r+Y8++MJDaEZ+8P/Q19fX23IAhw0mFNumj94bF42L1d53yXlAJWdvQ1DjMTNYpY0e+fZmdAHr6A99EPWbjfDD5i/nQ6U4a8uLTj+Z3zRd0nhfH2Io6N/R2ugV0C+gW0C1QdAvoGRZFt53eUreAbgHdAte1BW5q0aoNOYsLIn73bzvQm1q09tGqbM6DIqK4xlyqTLnypJ8i93Zx9Xm995ObVcHD8PHUowinoHD80cknHJOCE571L/Fqqu3AqDq+nO7etpn871dt4T4CObGuZKeMlKUg7bWYk1cyTr1t8VpAlVlBZzKdznQwM5qetD+kUxILxbW5nnzejL7PkhTvMa/Xk2O2p0qO7ExPVnKiLTplZ4TD5Ym3O7Kzw88fCokF+YZJtsUCfCiZZo4wmhR3OLIfeG2lADGs7DIERRoUTwRACnOWMTjdqHgdoGoKxfdgZF6cwXczrlAX6J+CQekUi4wMGfoWuHCJOEpuWfbiQjWm2Q02l8nrjgySHWboYKS5ZHNOefvJ0lWzDsSCFiocbbJIC6VIBhfAjbRDwZVPp5ij7ABJXMjoMIIWSsLYvPhbUDQp4WbZXNpq8EVh4ybhOZbtXZ9kV8Q9gPX4ndoN4j7C+4YAO+n85yJATi01kvhbgA/qe4/6niTuTUL8WoAb3DcBDDUwIQAQkRlGQIHABusK8OSiYHfDMFmKMkvyT+cUpW6Y7I41S6lWgxSOuqR9orgsM22YKcHsCfYTgULAhL8lzL5gNgYFullfLPH48hSKEA7nXGGhw5e876xLsW86qgmSZKBwbvE4NqBURmFWDNvQJgRTjJinHBePi+Ph8VwEdBqUD1drj6iGcunXOAAB6/78/RJn/IM9nniGQMXq35Yv6f5Un5e2Q0PCXwcECOg8r1G3QaMBvbt30tYhJdShfXt2EbRQb6NYN532eUVasz45/OkUZxbByuU/fsesgIAHgg3Val3g2l/+wzdf51VPu23NqhXL6cDvCMBi7vTJ49Tb+RvGbIe9O7dvKUifpLFixh9Fk39cNM8vJdONSJNg5opW1ykyOiaW9INTPxn1jnZftAWB/5FvDOiXF8Ui69E5HYgmiFRS7DuQRkXVmnXrkxqIdESBjpd0Rv6c5NfSVgW1R0HOWcDjzAUEdkKkuqD9xJUsXYYaKx63xz34+Se7+5uzeZ1n9X6QZHF+8cI5szo98vjTBBYELZOowyAfXlt5BfkQcHmwe69nCA6uX/3/oBszVEjRxMyh80ASmE3C8649TlLMkt6KIuugRNtMPRl1HR4L5/tP386f489GzJx+++Mps0riobvXQ+1uy+/dpDDn9UrHVtBzqtfTLaBbQLeAboHitYAOWBSvPfXedAvoFtAtcNUtwBcCf2njYseMgoyOK1HyGKLa/EXUiXqkRKCTIb8BM/2b+/QX/Zdf2/zGml/7QNsplpkAcl3tS1lR+8urHSL/m3K7AwKEpMRwOh0Or8fjEZFffMmS8QIHE5lzsrIy6ZTJqz9bcHAI+8rPoVKcx5LfeaCjPS+ng3osfFmF+GodTIqgnIy0HQcPHqBTz6sCMUR14VCko9A8ffr04MqVKwd0bNDhzzmrpbcorB18pwMB5f6iZhllV71OvYbaF+nC7sNffUExsnPr33Qa/meWgt5P/jMHXPgDocOd0e81UOgIxrxXSDcDOp/L5AfIbc577hEwpDX2uF2H0zPTXIbUEzFJqakZzpRTwfbEv61pTi9uJimxJTIOAigw3XgmuKLJ5s2OthusXopeI5vB45XlCGAPBoPXG44siRwAEKkeg9mbagrbBGCicognuzKonapQHwOj8DJLAiLcbo/BeALbLRaPg07qRAARgBssFoANRqvbHo424ZHuVIvsSsV1rWQaJMXokk1OUEylMqsj3J0WR9ACVFChjVI3lzkfFJUJsOQUtrmTDCVdRELQL4unUrAh0mzwOeSlLLey5c9k9+Zs3Dkv2MiXdSXABn4XAKcADdR0T+KsiL61AKnI0CCoIDIp2J5ZL4ISStBV+ajpcosQ2xaUdkLoWy3WLVUNlqxhJjmkrEWyRZgkZ7xViom3yfFlLFK5UKMUhY7DkOIixNUJVLBQi4EZE8yAIFDBLAruJwWF4AHtwv35W0gdJfQ0+CmExglEUAeD/bEPzrtDKMzcYSQ+98X5SKCEwC+/MxOD9iVNFQvnIHU3SGHFsRwDmMH6tA9BEfZ1GcUUtRvo3E4+k8Tj8C383aAI71fTJ35SqnRZAnYQ071cNJsZD4ycZiHwkJWZSZDl4sLfJ+pP/Lhw7hfq9fwOjd4a3L4b2hfabeq/wTIVQ779FUt/WJRXPbGteq16DfhbXZSMPo7zhUHDR9Jhqv69J4Bw+uTxYwXRw+A46jRo4suuWPTVzM/4TOFv3KDYqbN5/eXaHSJifpsmw4KZfnzG2Ljmj5X56UHRgcx9njr2/zoFYgw8V4yS59+BIuIhYlxv765tAcEZ0ggxQ2POZxM+1h7btbJVYexRkHkTqA6fX/hcXtCsX1IvTZ23eEWpsuUqDOz96EOBhLADnWd/4+C87NLz6T6k+RJaLqIeqcUICPL5NdAxtL67QyeCFgvnTJ8i6jCb6O2PJ89MSjh1gmBgW2Rmc1vCiWNHtf3gVPuylm7Evvp079hWu53Pz1y3d+dWvxRijz374iu3t7n7vo/ffeMVNZUUnznv6dS1x8plP34nnlMLe16vdGxXMjf0troFdAvoFtAtUHQL6IBF0W2nt9QtoFtAt8AVWeCeB7p0fxg8r3yhS0d01Cpw3/618uelf/7280/ajumA5cM8xfD4orPql59+eO25x7uqoxHpjH1/wvS5d+Clg+25bdq40SOm5qZl8+V08IgxE214I+GLFaOwGOXGCC++YLvQgBFUv/+8hBHAF5c3R42byjH27NDal1LOl45nXn59GB0MjLwbPXxQf62zuzWEHJ8F3y2F+xiN2PfRTnerOWt9kVRjJs/8etbUCXm9VNNBQucG6w8cNvLjeAg48oWLPL14v/dw7BwTAtTc+xDVOGPix6Ou6KT4aVw7F7AY8v7Yyfn1zWO8+6aadFIFXOb/sm47+aTHvT/MJ5DY8q7293d9vHdf8nr/tnTxt9M+/XBEfvspyPaCzBn2c+9D3XoO/eDTz1rVrRTH88hxUAASAo23glb75CfvDX2NmTisy5fr8V9885N48WRE69D+zz6+esXyJX60KXxRu3jB7fD0i6++1fCuzjWpAdL45lsf3Lhm9V+ofzGql2OtUbt+w1+XfHeRLoXz+YFujz1F+1PU8+tZn03IyxHEcb84+O1RbTs89LDJbDJ/NvaDd7S2JB1J/6HvffRwu1sb7Nu1/RI6MY7hlbdGjV276tflf/y67EdhY15Pd+NapfCjNqKWUbZtIAyJS83J64HjG/Dmex+xLQEpRiPyPPuj2yjIORR1mjS/rRUEKLuOGPTSs4Ha0dFASgitjci3zm3qa4MOhV59+78OmvPEiaPfeVMtwir6z+9+Upjx/xfr5tJAMUKe1E/I+PIio0IG37xC/ZLT0JhYr8gXfO8y/PLIbEjAH8sALqTKHnuW156+1pB5Livk3Emz89wRJfLUTlup5J1mh2KMt5gj7GaPMzTEnVkuXPJUyzKGHkcGQyUIwER7JAOcz7IdyvZBgBrOAbxIRwaEA7oUJ6ElUTXUk3UbtCqcuLrMwA5CiJ5gv+mEJZwGsyPTFLEXFE5lcfndAJCiLMALB8S4czAuAwS509EPsyVYYl1yEEYuZ6CO1ai45XRT7GlQQYWjfnhZ+6l4gBRp+J4I+iiCIAQuhYC1j3rp4fLmUlaD7HOK0hue4fLRQQnAQK1zo86S8IEduU1YX03FJLI3aFgPshnMMWbJAsVyJcl5Sb90xmspn3yXZW4RtFFq4EQKM0lGqHCYSgdJwcieMMchEaW8VYotHSRXtxqluDCjVNWCAwU4UQ+C2xloDKIsKZ5jzRXfJhhAOifOi9MoBBZ8gA0WZt/QUb8RZS8K6YNYj+AEAQ6fAHTukolPAg2k02MbAgxnUM7mftJJTIqpG3L7Yj32w+Phfo+iMMOCNmZGBgEdZlawL/ZDyiqOqwwK7UTAQmS+UDT8soX3EK7Mzs7k2HxL75dee9MLAZaZE8d+wO9cx98MbeMbch2ZfO6YO2PKp9rtdF4TlPCnUQHAwqdt4U/IW91POO7/BRU7pjOe2Q3fzp01zd+x5rdO0DDxuNSABZ+pqOGRX3uxXTxbMCPEXxuKWhMUom6AdjsFnnm8alFk1qEd+OnKwzEt+sIp9c3Nc2f/H4QS2/q++ua74pzv3rblsqxHbuPzwJJF86i54nch3RWdzVs3rV+jrXCtbFUYexT0vPmrx3N5YM/uHXkBAqIdxa8/mDRrfnRMXInX+/Xqxuf5QPsOdJ791Sf4xud+QXemrsNn+B35ZH+0aN22PZ9bVv18YTx8Jho1adbXBCOZ8UBaMF6r3AZ9cAKnlyxiv7yO1/7x28/a7eK5EY+Tl2nR8Jm+36tDR/DZa7ZGy4Vg0DvIvPii+rjRBDMKO89Z/0rGdiXzQm+rW0C3gG4B3QJXZgEdsLgy++mtdQvoFtAtUGgL8CWAD98ELAhOfDryrUFVqlWvRWcqUxm0gAVf5EdPnb3wtjvvvo+ObioHtL3vwa53dejUdck3/08jwPZ0rv4G8cSDe3fteKjHk89SJG/d6t98wncU2S5VtnyF83jJ5YsSB84o9DLl4yvRwet2uV0hYWGM2rxkQTR9Y2hl+qIub29zT4cPJs+aDx+FF77nRPI4MzpQ/SL0+HMvvUrHMfc5D86JTt0f7/3My4OGDR/Y1xetx4Uvd3SUE7AIZEDyL5MPt3v725sguDO4Rt36jeAr8YEXpKDgi3rpchUqIrEhiE7ac0lJdNQU+8KxUoBw3PtDX4cPHQuikfnFEmShU5ffuFNms2zGCNO5AAAgAElEQVRa99eqvAZApzrPg6jzwutvvf8EHMd05PPF/vE+L706c9LYD/LKoCnIARZ0zrCvWnUbNqaWCahpPNQFmfr1j78xcpQRf7fd2e7erRvX/ikAi9ff+Wg8HfM8r7R5l55P9Rk5Yea8lnUqxmipPNj3s/0HvcVzz/nx1ecTP+nQpcfjL74+fDQ23Zyrf0HafKUKXqYZFSrmEUG58V8s/Kl67XoNuJ/7Oj/yWHhkdLQA37Q2YATvtAU//U7qLtIiEPx4buCQt5d8O+9LiqWL+vDP02ks8RxoAQs6V3gNoavyArBgtOKgER/55iivLVw6p3kNiv5Id8FrNjszI4P0DgQeeY1xTjLrJhiIW0HOV351eE3lBdbQTjz+Qf16PULwSPTHefDSkHd880kAFpzPU+b9uEI4oziP3x8yoK92DPndT/Ib8391ey5QQSc6HfF09MKBQ5BCbisrbrsM/y8yEIJkxVOBUIUCn7GsuFKMSvZIRTYnmJxnzpucZxXTyS1phvMpYYbdvyjpdrfVopirBrky3UhHsmQZbCZkPrhO2sqlQ2+C9+o4ggMALNwAHsqFuDNAMSRLELoOARCi2I3WIFA4xSLrwgAgI8LqdZjcshH1DW4AEEEmxWWBJxuDszqQpeEEUGECrZTZi3GiPcGFVPyNep4YQCsuuPVToHFBXQxoUzhNRqwAXVQp9Os4ZS17BNkanlPWMsczTOFp6Dso3RTuAZBhwFilVINPX5vvF1boV4S6vAoc3PKJZKeyA1kKstN7UUOC902hD0FgQuh7MCNLAAmCIkpMJ1/KCkACA7IbZIh4+7ImQoEIZXgkb7bH53RXa10QROF+xPuOD1BBe1/2BsSyXeUsUlCjcDm6ArImAH5EhhjlEFA7VcT3ZkB8YlGH1E0SAIrjACWcaEsnPzMXTgH92I9P0j2xw1rYTmomAgAEB5hNxuADOvZoFI6N9fk3syIYGEAwgZkJ/N0dJvrCJ8EGgh1cWOcBFDoAf0ch2MHMCGZDMJtLAA2/4btI6eEnCymkaE+ReSL0OQjckCqKdqeGBvdHWwfMgLOAmomDYXYgP3nP6f5kn5cYdU2gm5lYpKXxl4kpss8YIU16o9zjuvhBOij+cXj/Xmp8XLKUKVcxnivUlEjc97HDB/argdZsDMKKBwVte39/UzeA65mFkF99/t6TkkodWMF7O9vh8ekyikM+q2j7ZLAIufa1VITM3mSQAzUe/I2DwDLX+wNySPGjFTRm3eysDF/2CjNi8js2B04m62jHzN9CPj/yuY/bDucGLKj7K4FnBP597MhBzmm/C8XS+VzEzEl/Fa6FrQpjj/zsFWg7n10qI+33u69nT8+rD2acMFCg5zMvDCTY1Lvrva3zo5AMdJ65Hz5/cF6K7BwDXi4uzEvXZfOSAJ06GIlAWNkK8ZXU2TM16zVsTDFtnjM+Zw96Z/T4m29rfdcHw159Ucw1PBv6Mqn8ZcKK63zBF5/7Ffbmew4BEUwZ3sMuLrw2Rk2a+TWBMwbAaJ91eIykoCKNrWhU2PNa1LEVdU7o7XQL6BbQLaBboHgsoAMWxWNHvRfdAroFdAsU2AIDh74/5u6OnR+hk3D+F59NZMPGN7do2fnRp55jFLe2IzocCRS8/erzTzMikC8SN93a6k46mtWABZ26dDIP7N3jQT7wL/1+4VxGjJ9LuuAg4EO/yJJ4+oVX3+CLUK8H292WFxUQgQFGRc1E5gLrEzhhFNnA3t0fJCWTliuX2QIEK5iaPmzAc0/w5SQO4Vm1AHqoj6spxCnJTxuIG5nixe2RAi4iIOmY6NWpLSNXJUZi0R4f4iVKHQlf4BNQiIoEEWrUadBo3ozJn65bvfKXQjT1W5VcwNyw8a9Vvz36dL/+BCt4DkcMfuk5B7wHSCgJv1Kwgv0XdM6wbsNmzW8j7zIdM1PmLv6VTp9nu3W4cwPGyPNPJzzrEWxhuj4BqlFDX3mB6zhfmX3gD6zgfCRYsWD2tEmc65yTdCo9hbnX/LbWLdf88Rs52H086nzxvjBHN65nVs3kud//QgDghcc737t5/V9/fPPbxt1dH3u6rz/Agk75jz6bsygaL729HmzbggKgzOyZ/8va7QQu1ICFO5cf/RDCYLUnSIifCvoNZh+9OnzUJ4x+JUgxYty0Lzm/1YAFr0n2Q9q0NXsTMhZ9NWPqmHeGDLzSeaJuz+Nr0LR5i09HvTXYX7+co6BsmIXMqdADe3ZdEomLCODadAr98esqX8YInRQfIivpDKhQxr735quDkHHFY/IHWOR3PynOY7zO+qLjlvoUpH3Cp9IKpQUyKiSDkm01eHMkRTbiMytBkYMaemXb7iB3wuYg1yEpLGPlgZDUdalO6F8bDx2OsCd7TGcdIaGphuhYxSuXPW+OygjzZNqiXClVAApYIIp9HmDEyWhncjWPbEqFwHYqMipsoHuKg35EVpYpBPoRDitAiRjqUkA/IhGZEZkWt6MMwAYXwIlDGFUM9C8yAEBkI1vCU9qRUMficZYD2AFuJvl8uCedIIgJ2RWRXskYgn7S0TYMbVxYZwToYQWAchRjO30iuMK+xSXv3XvGUiKnjD3B0+bsL5XRh+mGrIPhoIUyYox2tHOQZgq2MUw57Nx/X2lzaohBql/WZuhQO8Io9A8E3RGd6kJvgo5+kaEhHO7sRwAYPiopAAzmaiFyECoYQccUlOKWXCfsCsEKZhGI7AxB8eTL4iDAgcwIuVSQZClnlS032KQoZE7EVLbJVaFBUTnKJLUC+EHwSQHwsRadx6I+BdQvLthewe6VtqEvjidLlqVQpFVYMj3SB9j3eZtROgxQw2AzSHbUOYn1CaCPIhBAUEAABvxOZzcLKMN8AAaBCcwhiVoKFI4mrQoBDV8kMxYfUICF2ijsj052/qYzSpmfPs2HPHQo1JoQF7Mjcvss8EcO0sREZf4WjJo48+v9UGv+fv6XM7ie1DG8r/jrUAASgTIaKLjNdsAyCKJcsvDeyhW24NBQZqrxueCdsVO/4G+DOriDzz63tr7rHv6OiSh33hv5rNUYGWrqgAnQLPmAAPDs50kzxTrU6OBzlPhNZP90OvOZBL+bl9D/nTx65FA16DqIzFC2J4g+/ZtlfzDAQk2T43u2wO/Tb3lQWFUF5RL7oMaF2igMlCCdlD/9CtqIoJA2yp5j6oJsOwabMCiC/dFmfN64HcEw4lmSzuP3J8yYy9990nsRNPGnJcBnFfaRFy1nw6Y3t+Bzpz+w/VrZqjD2KPDFoKnI88hApEDPswyQuPuBrt27P/nci2G4eJZCw2H024P6a4XItfvP6zzzvMz67tc1fCaiEDbb8nmSbZDBegkQx7lmAMrGZwTW43PAZ/OX/Mbn8x73tvRRnnLB414sniF28B3jjZGfTKEexsLZn09WZ5Zi+vsCdARgoB4zr3MClj99+7VfjQq+S3BeOXOBMrbl0N4b//lXDFJ5ukv7Vv7mGgEZBoWIwKkL+y/4PGf9ooytqPNBb6dbQLeAbgHdAsVnAR2wKD5b6j3pFtAtoFsgXws0veX21hSv+3z86PcEWMFGjBziQ7k2u6Je42bNH8FLDuuKl32+/NEJSRok9Q6ZKbEL/Pni5fAoopj69nignb9BMVuBL6v56RaQioYvFBRlHImX2P27d27r3bV9a8FBrX5ZpcOC9FGMXKcjV2g0YKjBbgxWPY5GN916uy8yzI8wJl/8+gx8wyckSee4dvwcO9eBOvmqijNzHxXBR5GXKGW+J1xToVmLlnfyZQ2JIukEdvgyOGLwy8+JanlpjhR0X4WZMwSc+OI75eORw/mCCp9Q2JMAsUQkqPrlsUz5CvEcg5rai3zh/jjDSRUx6N0xE0idMfLNV54Xc3LejKnjTfBAhQVbSJshnJISwTC+6O6Hw53ZR+UqVKoM8OE24VCiI97njEKUr/pll+Pp+ewLA5k18Opzj3UhWMF1InLTo7lGatSp34hz3l/EZ3U4HdiWAAXnIOcyxyOo1/q9NmwE3qkZXX3Zwhdxju1qzMma9Ro09mWfBBCzbXf/Q90I0Py18peliQknL6FpQCTyxWPioHkMuE4jnu58T0s60MhZfW+nhx+lg0LrVCrM/aSgc/N6rpcrrs3nZtINMesBDjtlDLIqbDJ80vBVSwawIpndpwFYmEJM7rMpADA+B3DhQgLAusjzC7aHZq5xyfZsj+GISVE8cpzBYjW4PZHOTDn0bGR26tlzQTF2i93pjHCnSaB5ys40hoYACECEvxwFGqeKADEAUgQfxzaPQfJEAYzYD9qmIIAOGJOcDnDjFISxa2Kb0w5NibNBcXuQeeHMNIVmV8w5VjfCncFsAROuPDNAhf0Qz04Jc5sq2Dz2KGRdKAA+cgB6gOoIghaKR8k0Rp+0eXNC8d2VEhR1+ExQ3Jn2SUviIlxpIRVyTpRDVkZEsjnmzNro5seQcWHHek8wjoHgCa/vWuHGIGRV0DlsAJLgPZzlZYaTcKALeihWFvRNvCcIwWuCD3Ts+347AATIraPl0MbhUtl0t5Th8EreLI/kWZOmpJ1xXszI8LUFYKCgGCNNkq15pBxd0SqVqBMq14IGxa3YURY6NQNMaM3+c7zSbuyUGTO+MYP2qbmYp9jHIQAiqwBEZKM/83G7siXWLEfg++6jdiVrW4Z0dHmykoGBhiIbIy0U+hapLkk555IYue7L/rB3iuRxuDB/RLc8ViHkzXUELpg9QTCCDn/SsXCOabOzGLnfBeU+lGdQOAfZKaOpedwFEs4WgyjsJ3+bmEHBrDpGiBNQ7v/UIw9c1HLCcwJ/1/z1WwnR54zcDgT6qykGte2ZScF1A4e9PwYMe0mkxeRzEu936rrLvl8wl/dC0hvSYVoR9JGdkSVQCRoY2sh3AgH8bQukG6Dul/sizR8BGmZkMAqd2SQfvvXaS9rnpx8WfjWLWZNjPvvq26+mT/okAqkVzw0YMhyYRdn3Br/cR91vPFAa3tf3BODzZ13Bu6+l7CtboWIl/sbxmeurn1ZvmjxmxDB18AaDVZj9Qgc2n8caNL351ocgpkwqrOGv9KOgu29hlDzpfxggMjgleSIj33s83e9lUlG989oLvZnVazAajP5+HzAVOG8lCnNzbtzUonWbLj2ffO7VZx/rIrIGCJjj8DYS7CeIIuh82O5a2Yr7Kqg9CnNNkNIUPvOMlchovhmaEWxLAILZO8ykYLYq9NIb1EWWCZ87CKL9vnzJ95998sE7/jJm/O07r/PMZzQCSk/2Gzi4CvTokPhQgdnQzLDe8OfvK9T98TkbCQqHWrW7tyOeEY63ad+xc+Wq1Ws+0/U+0tJdXM4mnk5g4MYPq7ceKFexUhU+C73/5sB+6jrb8RzCIAdm1g54unsnAQ5yPmIMFb9HlkkgHTJe51qQhpmwfC/iPkjxSiqp1SuWLaEWCJ/fmLH6ALRU+JzKTA/1WAp6Xos6tsLMB72ubgHdAroFdAtcHQvogMXVsaveq24B3QK6BS6zAF9Oh42e8DlfVqZ+POptdYXmLdu0Q7DiZu2D/kuD3/mAoAB1BET9eNAkMd1fy2ss6GgKYno6eNf9kX/GAIEFRjU1v/3OtuQ7ZpaDVjBT7I8aG9GxcSVe6tW1g4i4Z3QkeZ7VjgoCIBQSnIusBX9jvRtOB2pVMFXdn75F7fqNmzJqXk0RUZBjLkqdWvUbNqFDZtvfl3MwF6U/2nMr+np1+AefkP5o5NBXni9KP3m1KcycYcYHnREImrPe2b7jQ/16PniPlrZC7Cst5UKmBcGI/Mb88pB3P4T/3oZMjOfVYqKkQfgEFGgw6UVhXXw3Llq5sdluRLuSQ5kRscP6P/eEOvqVFEucU1qwgpG+vfoOGETnlTrzoRooQzhGRguqx0pghFGx/iI+6VygA4vRrA/16PUMKQS63d2ioZjLpH4KdNyCi3zH5g3r8rNNYbeTw5o2JHiibUtg5WmI3nL9N3NmTNVu5zFxHe1DDms6G98f0r+P4D1n9gY5ufyNqTD3k8Ie03Vanw7keBRGwYOmR4F2heIDKwzeTMkrh0oeQ4hkUbKTIWCSafSm/YySEJM6wxbkOh5udIKhCVRMSMQwGjPcYV6DId5qc5aICzmXlWKMOgIAA3oU7tAck80DkOBgmDtDMRo8QQAQSiRaSu2McSbfBEAhDGLZ5Uk0ZfJ6JFAwWQAOJEW6UqlXkY6Milg7BLTR5hQyMcLDXWmhLkPQkRhXcpUSjjPVUNecYQqjzkIUMiMiQem0D3ROScjYiAAgEgsgJBzghBk0TzYAGCloVwYMhEY3ZDPis49VqJu+4yarJ8cKcCYV4MgZaGYkoo5U2p6QfSQ4Pqe0O9FMcAP9+7Qn7illwlh92QWS3aMcSUKKAhb+x/cPFtIL8W/W4d8iQ4KfXOcDNeJtkqmEWTY1CpdKh5ukkO2Z0gm3V3L8naHYAVb4MhYAaBhCwF31QAk5pkaIVDPUKJdGRkUdUDvRmWjALAfOIFkAQhzGME54AUKA8yoUK6OAHqSjE0aMk1pqfaJDWnEoRzm8PFk6kOBQMkqC4A3bsg5kQ4DE7dPhENkcPB4CLhcoWC6MRWRT+A7WuijVA9DiEhFrFXgh7EFNiT9RKEZLCigCoww2YPYFs3nUC6l+7kEhzQ4j8JmpdhTlEiFrTZsr/pP3TAYQPNHn5df4nMIsS/VvBdhcEtpCZ4cOWy3dHm5TRmaeBaK1YxbCWYhf+NOg+HXJ9wsffnx9P4IRbP/z4m++fgv0ktq+6LCnFkD7Bx9+lIUHTE7/gc88+tCKn77/Rm0AAry/Yl1eNHuiPp3Cb73S98nBIz6eSMc+n7teebZnZ7Xekqg7d/qkcbe2anM3M0hZuP4MyP5feKLLfVqwhnSX3E4QJtDJ4bMSnc3aQAZqD9FRzHOxZtWK5Vs2rOXcubgwI7YVnMoET7iSvx9/rFj2I6PxSW+prjsOv8fMcGSGL9cTHBnz9uABPNd0vDOrko5oZtSq2/F38ocFc2Z26Nz9cTqwuY2O8gOgIxX1gJ8fY3v+rjKgQN3+WtmK+yyMPQp6oRBo6v5U35dInSjajJ765SXzjDRGu7Zu2jj/i2mTOF8COfID7TOv88xzSpsSHCNdJYMVmGkRSAPt01HDB7/36bQ51IkgePTyk906MhBJvW/WoVYbMzBIITnxw3ff1IrB87w1xnNs01tuax0aHh5BOlP2EQI+Weq5AJB519/xMPODeiJqbQu+E/Xq0/91ZtEu/HL6lLDwyEiCKgS4OPdFP6Supa4FqUiLMs+LMraCzgO9nm4B3QK6BXQLXF0L6IDF1bWv3rtuAd0CugUuWoDp1Yxc63n/HTerKXSYgk/H4pxpE8eqzcWXSIrzMSpNLdpLOidG9jFaS11//Z8rf+2ISCSK4jGaMZDpGTnF6MhtfoQQtW0YbZWZkZZGRycj7tQCk+q6BFC6PPZ0H/Lnq/Us+DJLfQFSRIn6dJxeEJK83AFLgKP3S68PZd2l3y34yt8xkMIIL+irr8XUqlWvUROKfRb2RdPf2KgZwAgzOgEgIVKyS5ub6/JFrDiPo7BzhueXL6TUE+E50katqsdGhwWdFLfAIeMv4lLU5THSsbMY0aYi48HPMfroXVC8XR/uFvv6h1NqfD1z6vhXho8au+qXpYvpCFG3KVuxUmV/c/pBAAvMgJk4+l3fnOHCudiz9/MD+BKsdrLQuU+wa8608R9rx8PsiEqIeF0EyjVSfjz5/MAh8zAe4Xzhy3Ys0iv8cYazLwI/dAJonTrFcW7r4T5Ah48WrGHfpEchuMf5qdauEPslPQn50ekMfOWtkWMZtajOWiL4RGDCn+OuoPeT4jjGf1MfGmcyh8Z5KrQW6IQmfc1j8K1DWNsjyV6HZPKcl5CSsMvkTk4MzV6dY3adTMG6CIOSs9XqPGBHlkU7SE20Rk8pslXKluMg2JysWJChkBUSlhNVIeuE6YStfFqp1MS6Jpcr3G607c8xWCsDhCiNOsEAD9zUrwBgYQ13pwdDS8KdZQxJhYh2IqioMgASBIHyCToVSngQKaO82UZQPoHVSImH9kQ1ZGmEgV7KhmwM0EIZeAzp0JwIAtARdDQ4fn+EO/3GUE9mONYFu2STC1oWLohsnwhxZzXFPgwOxZKNzI3K2E8ZZHnA52/IQb0EbDsT6zx7yz1JS+vvDqv1N4AOA/ZrRT8O7NNrMcg2h1c5iM+qEMZOOI2shFx7iuufzn4BVBAQFBkWtLsbB+BuFyOH3BIp1TztkDIAMmQhq+L84RwlNcEh5ZDTqrRFCn6whFy+WrAUCwDCWT1YfjLYKN2F/Z0GGKF19kvoszJ0KcpCpPtLbA8DeJF5yq7sQ38nzrqknB2ZUjJAirQM3Jmpi4FxOJFZwfPPrAmOm2PmWH10dihCIFyALlxP2hSCGj7QQruAvkm7SsG8I3jDfbAd++LzQBUUOrYrovhojHIXZk61R5mFwt9CM9qzjRA0L8g+/Q0tz3Xj4dBc/sM38/A7cFibXcBsQTogBQWluiPqUOXV8UtPPnx/IP0JUhY9/kCbWxgMwSy8QAETvIe91Ovh+xnNjkeqUrzvEWzwt9850yaM1Waz5jU+/jYu//6becxA9EdZI9oyuIO0NgxMKAktpDP4RSDFoD+axzWrfl1Oik6CKoH2zUzViaNHDCXooa7D+32Pe1s1Jb2Tv2h9OpE7tWpSk9mWBPv3IRpAOJa1++Lv6v23NahKqk2On795FFdmPWb10q6Myvc3RgYWzJgwZiQ1Ok4dP3aEvzPqeozAZ6YBdbC02bTXylYcT2HsUdCLgjRJLATbxs2cv5jPdaOHv/5yZnp6WgYMSHo0ZiQVtD9/9fI7z3y+at+8diVq0uUnOE/QrgWez5mVkwKUzF92M7MzWPIaM89b30c73c1ndfXzK/d/d7OaAYNZ+M7DsVKHTvRPcOyem2vHq98rmE3OdyIGl4RFRETyeuM7hT/qsYKe16KM7UrOm95Wt4BuAd0CugWKzwI6YFF8ttR70i2gW0C3QEAL0MHbFfzBTJXXUrs0b3VnO27nS526Azr76aRU8z5TE4Bi3W8N6NNLvFSKNt/O++JzAhaMDs+LR78h+PDZRhuVpx08I5zA5FDbl82Bl1itE1ldv1Xb9h35IkStB7G+ecs7273+7ujxixd8NUstbsm0ddbRRr9z3f1dejxBwIXf/TlgCfhQEDq/sRfXVKSOQSAndWH3QU5pnudSZcqVp9h4IKHNwvZ7JXOG1Bh05DNTYfwHbw/Jb9+cY8+/Nuy9Fne0bR9IP4QRhzxORMOND9RfLgORz5l3NjWjIetXA2jHF++Rbw64hIKAQA8pOJaB5kLbH68RXk+CO5qp/x9Onr2AfMh0lqjrM2OCfTHDRdsP5zntsH3zhrUdunR/HIBamFovgyAftwdygPGaulpzsia0anZs2bheO2ZmRzzbf/BbXL/uj99+0TrFaFOe319/+m4hs7KYQUORT7WjIh6UZ4GOqaD3k/zmzPWy3Q9QIYZO5zSzKyiy/QR81n1B8QQOLZcFzEnwsF9g41FkSy0Ibu+Cz93kNFc4ZXPsOGBz7PSinhUu7QxUqa3YJa+Sg8YmKVKOkCK9SZILgIPB5sopFes5Gy4bvcEWpyMMgIUxIyjcJnu9pahJkUvXxCh8DzQlACi4SQ8UjCyLsgApDGctcZnIqggHaOFBfTtACi+AjiPImJDwtyndEJZq8HjjghSn67wxai9AjRLIkEjKMVrPcvDHbeX3IsMiHABFHDIRsnF04UhYcIe4wTKl2EKCPTnhAEvMDqPFCqAkxSh53GXtCdVACxUBMfAoaDmUq52+c3O4O81zOLiyBGFuQxzgkxrhhupmg1waXv5MoBwHd6V7GI2rBi14HIIOiqCA0LOQ6oVJlg6xcuVosxRc3ipXhSh2OrQqtq9KkRJQ0fRiebl+lWC5otUgxSOLojM0JiIBZvxBsIInDh1dFJ7FvnfjZqOcdUqr0Mfe827p7I9nlT0AK1zQmjCmuHCwiuRwUSH9AmhCIXJqR/jonGhrFGY2UBicJ5zbuYjsEAG2kBKJbVgETZPQ6cjvUhDt6NAjtRsBCoIXPEekgVIv8fiDwEnf3LGI7CpqVKg1K/LbZ6G2896hzZ4QHTBaWxuxXdDO6ZTk5M5rCeRw17YpiC7FT9AQKOjYRD06XPMCK0Q92qggYt501qqDO/yNh5kVgWgitRm22vYc799rV/9ekOPkWJipoa3LZ0xGtufVh+85JoCoNgEMLYih7uta2Yr7LIw9CmIzUYeBCmtXrfiZ0QpXQ1Mtv/NMQCk/sEKMle8TyWftiYU5vkB1ixJso6YTFf36C4Li8agFwvMab3GdV39jKw476X3oFtAtoFtAt8CVWUAHLK7Mfnpr3QK6BXQLFMgC5N9npJma2kk0ZMQ6v2sdqeDFvYsvQHxpZNvX3xn9KUEApmkLoUv1zulYJyDS6ZEnek8b9+GIQC+6zNrgi/eRg/v25DV47pNgBetMH//R+3nRJ3CsfMlY9+fvvxK4ePql194khzJe5JYLYWKxL4rf8SXjON501funA/ap51/xOc15zMxs0I6PY+e6LTjOAhn+Cioxqr5arTr1F/mh2ilKt6ShYDu+6M2cOHZUUfrIr01h54zgyF6MCNJA2TPqfTKKloKjTyCN39/LOW3WrmPnbnQa5ec4ygUt5Buq1fIBWPWg0Dl5zPtvaV8cBdBDijD1WEqXK1+xYuUbqo584wLHMnmQSWeA5KFyjLRVU1NwO7NPOIf9AVCkMWGdPdu3bqIoNUVJ1dePEI097OeaYQYRx/LF1HF5OnbyO3f+thNgYRYEwQPt9vu79niCAB7X+8uWIsjC9rvAIU6Bd1KSqB1YFFRn1PLq35Yv8bfvgt5PinJc11EbRsrHcfqgdEPp4fNFI7MCC6LhDUGgeULyhPO02XVqPTIpNgTnbIiAjkWGxXUUosyumqheF1vMnPgAACAASURBVC5wUvuUwWcpuOeXwhUeC3d2HSgVQPxCCTM7XO5IQ1rQeWsUJbAdVq8dfnjvObdkCjIAnABY4MLfwQA3FGhSwEtOhiPFbPHaK8O/ngOqpwQAFmbWAS1UumKQg0EXFYsMCge0LCygcDqH+mmh7ozgcl53dYAVWCc5S9ldIdHOlCAIZR9CsoIX+hheMlZh/+WxD1IoQSvDGwNQAoLahlNGjAPZE7QHx2NOM0ccwNiOAUAxdUz8rsK5oNjjp6zlFNT3Vi0d7wo2yjgOn+OfnErHs9y+DAI694WOgxCkpuNfFEO3UnKpVlFyfadXgXaEnImMCFeKQzo467RyCtxX5p6l5UY1Q+RuoIciNdLFBZRQLcUfyMZISXRK3yOTYufmDGUfwAn59xTlPEALD3Qr6NTnueU+CT5wTAJkEILgIltBAAkEHoT2BMEVtuc6ZkbwOHhsBDf4mymyLvgpsjDUQ83rO/dH4IFUT4dRmGHBfTHQQEQwc19CjHwAvpdEIaBL2jgCHAJQKeg+9Xq6BXQLFNECpFIqYlO9mW4B3QK6BXQL6BbQLZCHBXTAQp8eugV0C+gWuAYWaHd/524Um1v586U0TnTS33zbHXeR61atycAofDojl347/yuKEDOrgg5UilxSCC/QkCeDw3bq1z/+xmyOz8b555JlqjXBkfz4mxmRzv0QiPhlyXcL8jITKXF2btm0gXRVj/bu15/6BRRyJp+ulgOXlEEnjx45pI3QYmR7dGxsCUasAavY4W98dSBgyDT5gooWXsmprVqzdj3SA20DEHQl/Yi2wp6MHNOKIxdH/4WdM8yqIJ0B9006poKMgXOQdBqk7SKFhDaitgl5jYFY/bx40fyC9EfQYuz0r5uy7hlEY37hJ5qzKsQWuV0LWHDOcX0O+NI+/2bZH8xyYDRi9/Ytm/jT4ajboMlNXO+P3ov7IN0Infy0izpTiPsgjdmFMey8BDThOl5P/Nz29zo6GIt14X6ZKQHhWfLVX1x43+jVb8AgUnRxzBTC1O5Y2I1A1IChIz56CkLb6jpC6FZrV3WdgtxPivWA/12dMaqeItUUYe6OcnuurrEDVFAWWbFnBblPrjR6UksDoNgf5DqaYHPssQbbt5YxelNzAGSEwAXOPsqjJIJU6oxswf8uqYIXfxmClTQ5RooyWz0pymlXssHhLWM0hUc4rUEWr1sp5fBYSAGVBeDADBomo1MGkKHYswEmRABwMAOYyEH2hAXAhAM0UVugTdEG47OCLsoMwCAEYIUbGRcysjVSAUgkumWjLcjrjEZ9EzIvZGwLBtBhM7rdEaCAcqBNttnrDAWNFPz5Bjrto1ASAFBkQJE9CJRUZuhi+JAa0D0dwb7D0eYMNDBOlLEn1CnpSIqNdp5PORJcKftgSBX5RHYFGfRLZYGshMOrrwB0qBofYgjame4RVEnsi453LnT8y6HQoGgRJVs6l5BvRcaEEVoVm6FDYQHQ4VyarGxzeiVLz7Jytco2uRnQFNrWt8DDn4ZMie+gZ7ELgIbpvEva90eqcmxtmpKeDVonrCcIIN55CCpw30JHh45/fldnevBvNYgitrEu1wvdFwFiCNqwMNUUFn1Sx0KijkUhFo6RNEDcr9DyoCA3wV1GSLdEIa8UgQmCGQDSfPOMmQPMIDuCwmwQfdEtoFtAt4BuAd0CugV0C+gW0C1wXVpAByyuy9OmD1q3gG6B68kCdDjegsyIVb8uXax13t8COigkJERp+ZTrNb6QSQAu/cF0sH4+fvR7syaPG63ljdbagVQEpMjp+kTvfhTN09LEkO+fTtCfFn39ZX42ZGQ767BuXunfpN8BtlKZhYKTy8BxPfmjEcOEsK92P6T3OXbk4H71ekbmM7ti4ZczpnR57Kk+gcSLKdbNyO/8wJb8jq0g2+mIpoP+6KH9ewtSP786FB9nnbyotfLrI6/thZ0z4vwyE0KbjZDXfr76fNInj/Z+YUAPAFNawKJZrtAo9Q8KeizU0WDdKWPeH0bQQNuOwBHXQav+ErCgfu41MnzMpBmca+TT/nHRvNnaa0z0Rz7vDX+t+s3fuLgPYAK7SWc1+7PxY9SaMawPeQtfVtCRA5dnJXFOklJDO76CHn9e9cqWj6fDXNLqd3R8+NFekVExsYsXzplFbZy9GiFVthF2Y1YSsJRVWvqR/wcsLgdhxJjyu58UxzH+S/ugk5gOcTrUGbEODQH6vOGpBkhg8EkxSKU9oFqC/PVyi+uQHJU+P8LozThh9KYAhnOXQPUQ1KEzGXxRgClc0ndKulRTccHp7JTWQ3x7LXIPWpjD3JW8doPTkRbkMMV4jaYUt006L5VyK6bTNjn7qEGSYyG96zK53TYAExTDPpZhDINDW7EBRLBDS8KE7IgbARiYQNfkBqDhDjI407EuAdkb2aCvCgFIYQXYkIWsiBMAGsqCLioEdeMAYJyIcqWkAhiJwd/J0Kkg3VQQgIgsABoRKPsh8n0W7Usgs8OAv6GVYcySvIYzyO6oVM5xuk2OK2Ub1rudUlACPnOQieHBOL1m+3mTRwnNgCefzvwgq1GOAIBByiShU0Fnu9CwIAjgahYhy73LyjHhRmmfR5H+j73zAIyjutbwna3q1XLvvXebajCEToAAoYeEFmoSSgghhDxICClACoHQQ6+mN9PBmGKDce9d7rZkSVbXtpl3vvWOWcuSLduSsfG5753s7sydW/65Mxbnv+f80emVZp2ogPu/rnAWz6s2Hkn9ZETLYmPfNFMpehWVEjXxtkRShIoi5oXn1ztTvpJZC7nhSGqnkJwjasLVdYAAcHUnkgkHjm++R5ujI5J1INyIC95J/PeSq0fB8RIxIke4x5S4yHiiDt+pD2HQqKZE4rrGPugDfCAtysTQECAfPlGHEGgdEhcydregc8FaZc2ydrk+TjBpUQQUAUVAEVAEFAFFQBFQBPY1BJSw2NfumI5XEVAE9jkE0GQg/crUSZ9/Wn/wx5x0+lk43+s76ElrQ120KF5+5tEH6ztQtwcCDtc77n9iHDoD9aMxBojoMNoUc2ZM/XpHQJIOiToisvnC9uq6Y3375eefuvfOP928o1ywBZJCh9RRyW2e/pMLLwMj0tOcd8mV1zS0YxxhZJywpKfa0dib4zyOXsif5iJH0BMg1dWXE7bNFd0c493ZNdPU+1t/bAhJuo5y8ZkXJIshovkBwbZgzqzpTZkTqZRIS0SkQHnR6qcE67ied/K1vUSRnqib5AgkzqNlQtTSn2+8+jLWeUMikm47iILyHD50999va2hckDdEIvQbPGzEry/dWvuC+qSEWrpw/lxIi/rXQ2zNnz19amNESVNwaKyOBMDEHZPr1qzaInrKc/Dzq2/4A1EgjAsh7XA4tE0KGOYEPj88/ezzf3vFBWfV76NHn74DWNvbEUaPX7K998nuzG0vvhYnMHoV6FYQgUQqqISDWGgA8U1LdIXx2tU438uivjaLcipfr0oJL/mp+L3zxXAYs50e4VqeA97lHYSg6Cru+S4SZZEj1s+pNKOdGqefuKMzfaFIpmgvZHgqS50qb3qtzxuJbAzk11T5sqpTIrXVQSvkF1HsWrQrhEzIkaekWnQl0oUgIPoilhmt6kMkhKSF8kn0Q6ocW1fqz5uWGa1sL/WyJZWTR0beVnQqWsvnRvlcKZ/dpJ5H2qwTd31r+ST1UEzaqJX2U4XEyLKDGZnGn+PzRGpTUnLbtrItv08IC39qfqcjrJpNOU51qS+zw6B2tSl55Rmb1ub5YuFuF3XO2dQtxTv7Fccun1Acve/Ytj5R/7aGVESc+zumeVJPbue3llXbdek+E8sPWIHSsGOJ9kRQ0j8FhmQ4fomsGCJi16EpFc6ibyqc6Mq6OJEACRAsEVHsSeVmTdRxHhdNC3tjxFQ+t96JSZonr4SFuFEPbmSDSyJwvZv6iWUHKYHxLLs6F1zLfYOEcEkL6tIGBmlBGxABEBPJqtn8txTt1E8d5b4r3HHRXqMFIe4GdFToG00LGDLWG6R3bzFIDCJgkgtrlLXKumNMrOONYpoearvI60lFQBFQBBQBRUARUAQUgb0RASUs9sa7omNSBBSB7xUC7k72xeLFTZ4YKXz6DRwSFxyu76CXrDTi+DJm3JOP3NfQrvPtATThvbdfx2l82FHH/bA+YSHZmOLpdWRX/bQdgdx3wJBhOHHnzpw2ZXt13bG+8/qLz+2IrEATgyiPkqINW4T/ROA469Krf/uHZx+9727xz5LWwjQkBCz6wP1IhTNPdAZ2NPbmOE+KoReeePi/zdEW6b2IpEHss37US3O0Txs7u2a4v1z38btvvrqzY3hLNC/O/OnPrzz48B8c+3ZStA6kwLrVK1c0leQZNGxUPLrilWcff/jjjz+O1ScrONer34BB077aVrOE+RJZ8dE7b7yyo/ETBUGdmVO2TduEBgX3BoMMq66qwkG4pbDm0Mpgzg31gzbJa88/9eiOxrAr5/MKWrchuilZ7PUnP7/qWkTBSZ/1/DufT2tM6JZxQdS4WhT1+yfCYo3g11CKrOS623uf7Mqc9uJrcCzjjEajAcIBXYAfick7yfFLZIXxODXGG6swvtiGl7Ir3yhKr5saDkRW5vujq+RZsvOkLjvaNzu2LTNNXNgd5bOPJBxqY6WIA9lvikTyYrJQGn2ccJwEWS/u8BJPimP50mPpwfJQhRW1lwVNqK23KtazyNs66pfYBStgqoRZCNWZFFsIhRSJkmglUQ9RIS9YqyLEbWXI9zKJnCi1Yk62RF0UZVvl7TOiVZLuKVrn+HB2i6S35amcnj3syQ51ayLdapafL4RFK0n/VCpjtDlX7UtfLFEXEkYRPgqR7dTMnDa+7gcE7cIpfvnMMf4UoRXSsnydhqU7oUrHLlkZ8g867qwsrz9aN+vdL4O9Du7gaT+g0zm+1M+OiXpeFrTClVEzw/Y6ZWk+c8bNfYPBDSHn0+KQsywvYKWLMPcRAct0lYiIslU19ie1EXt9VWVdK9GmaHNYjtW2TcB8mu+3MiRaIjRug1Myq8oJTS53YpPL4w58N+LBjZ6AbICsgCjA+I7D3yUMXAKDqA6ucbUr3CUJ4QAx4Ypk8xvyAk0KV2ib9cFvN4LB1ZIg0sK99y7JQbtxEqOp6aAgLRootBETMgNdaqLMaH+FGO+0i5LqMzb+/TxdjLSRGxJzQejcJVQaal+PKQKKgCKgCCgCioAioAgoAnsdAkpY7HW3RAekCCgC3zcE2ksOJOYkKfrJQb2l/PLGW/+6VjyuHTp36VY/N36WeGOpGGlg5/SO8GEX+LyZ075xiZLk+qSDKlq/ds2OnJQ4b9n9/upzTzyyo/6+HWt4hzs5EQGmvZqaKkRF4+VSEei2HdsWIeo7+N4QVhwTwiKuI9CQGPeOxriz57v26NWnQEIWpjfgKN/Ztqjfd+BmcuCLT95/Z1eub8o1O7tmJHBhGMRQQ+TQjvqDxGKd1V9jRFygP7Kj693zA4eOiOtXQKxZ1r+2iqzgOEQPhBbaFPXbZL7oqzSlryEjDjiYug2lKXNTdUEkPffYg/fUbw8SBtKiId0UyA40O1pqTfK8SLapLc8KmiMXXfXr3z0i+jThUF0dgtwb3liz1XuF8QsvmNZBUrTxnQiJhjCCsGhIrLt+3e29T5qC/T5UJ66jIObqKvxQvscF3cXnLO82Gydxii+6brFoV8zKqJ1UJmRFT1+spJ9oPBTKuY/EEEXGod028dlFXNaSpEg0BSSkQUiKNU6RWWhlmEOs1tKXT6zGLJXIC4/HcoLecCwckIiBcMwvpES0g6RWCkVjXidQF0kTtsTntWLyf14R0k4JSwqnmUJUlATsEJESGUJkLJY+Q0JkDJXIilZZ0cqoHK8R+iEq34uk+/WiXeHpVb2oMidSnimkx5diw+T4yoAjPUYieVK/QEiPjkJWxJ30Tm3ZSm8s3NWT36XOm1ngtTLy04woYHja9CwTmYtO1uATC0xNWZkQGVn+/keu9uS0D3hSMw8OGOuwAp+pczweI0rg7Pp3BFiiViKpXqtbtzTTQ9iGVcIotBaNC/59DGRleU+sjXke+KbOOycWi7UTzYthnVOsKiEvhNcwh93Y1Vou+aamL69zZj6+1myQCAyc8K52BO8Ol6Tg/rnkhKtd4YpfQ3IQeZCcHorr3GsgM1zdCG489TlHeic3uoI2Oc51EEau+Db/TcV4XCIlmfigrd0ttAuhwvMOCcFv/k4gEpJ/e7uKHZQw5v+/xNjddb3N+3V3B6TXKwKKgCKgCCgCioAioAgoAi2FALuPtCgCioAioAi0IAJpshua5sUf6qafMINHjD6I9EYIBhMx4O6693i97Og04qOM7/JGvHpHQ8PxiFBwcj1L0j4l9+eewwFcUly0JbqB6A5SH9Xvo8+AwfF0UOSw31H/OzPWoEyI9sTXGtcqwJF/3sVXXnPv3/54E/oc6FuQcqihqJL2Hbt05Zrk1EBcn5qW5uYR39FQm3z+wMOOPIYx1M/73+QG6lV00y9N+fKzHeK5q33szH1AM6SbRKw05f4yHtaruzb57ZEf8TUti6z+eHGW1z/GTn9XMyH53AAhLIjKKVy6tai0W6dXQnC7IbKA+crjscPng7ZI20SkQUPYumLon7z71muknqpfh7RLHFu2aAH547cq7Tt13mZN8oyRrmpX72PydaR/Sn4WbvzzXfeWCvHyzCP3/dvVtyAKqn5fEJOkfmM+9aOsqAuxhDU0p515nzTHHPeGNmT3Ok5d3iNEPYwVw/F72uaxwTTYIrId6WHZdd+khBd+kVX9geOPrK7wxkrXCgshTm4brRHewby3+duaZ6CnuK9JKdVRmoiJBSyfpIPKllRTKSbVEte/RE4UCGnR3ZRLBEe5XeqtjbX2ptsdJUqiNmBHwllOhS/NqdmUYVdm5UY3FaRZNZJdyd4kpIKdate2zw2XZknKpyWiT7FByI3eIrQ9QCIqHBlxpohsiwyE/BMSq8tJj1b3Fn2KGvkuhMWSsQXh4h9J9MVQBLvleBvRqeghpEU7ITTShayQrExOWKzEE6mLWcWLHV96jmWVr6u1qktDEgsRdRZPLHaWfjnb1G5aJMRFwIRrgt6ashEmFm7nRMM1xpaoDjs2X8JS2guwvPNx+oNNrWhP9BHrLCDlClnRSc6nivnlWCfRuTivU26K/WW581TENl+me+NRLsVSr0AiMY7J9plf9Uu3jrupm9XjlcGe3D/3sNKEyEi7pIPlkgcQC3x3IyJw5LspobiZOPmJznBJCrc+9VwBbTcFE5+c535CSmBcD4Hoau1AUjA3frt9uaRFcxMELinDv99oVUCgvSU2Ob7WNo/PLaxd1vBYMdZ0emKNJ1XRr4qAIqAIKAKKgCKgCCgCisDei4ASFnvvvdGRKQKKwPcEgfJNpYhlmvadNjvc2bn/t3sfe+5ff775NziC2eWMfsMjL46fgPYEdVYs2yxKXX8H+7BRBx16278efIKd1S48/3v53Yn/ePiZVyAfODbq4MOOGHHAIYdNmbQt2eD1+XypaZujHCg3/+3uBx8ZN34Cu9iT4ZY0PG7qqB2mX3IFgeuPFfLhhj/ecfchIsTttg1B436HZPn7fY+/sGj+nJmvj3v6MY7LZvWcogYcsJxj7HympmXEx3/iaWf95NnxE6eOOPDQwzcfT0vv2rM3edh3u4w9+oSTp0+Z/HlDmgW70jiOd4iWYgmz2ZXrm3LNzqwZyAqiBhDc3lHbjP2J1z788rJrfvt/bt0Lr7ruRkiP+gTM6sLlS/v0HzyUtF9uXaICnnz9o0m/vuWvW+30x6Heb+DQ4VMnb6vt4l6L7gff0bioP07mS/RDIBDc4qijTdbFLXf9l93F8cI4ST3VGPnkEhKNRRMhuE074vtHAHer4pVFmbwmScP03LufTzvnost/tSNcm3K+TsIr3HoIgv/g+JNP+8efbvo165JnJT6uepFbHHPn9Ma4Zx4npVT9vlzyqKE57cz7pClz2EfqsIYgmVhvOHt/K+a+Y9eJbsXHgciKX2fWTPyXL1Y6LbVuxlJ/bEOxx6kTx7eTLXWJqMBpjFOZ++Lu4EdPAHWFFDG/kBPthag4XI44ErMRkixTRF+Uye+w/GrnSbNT/bnRgmB2eIVEU3yRmlFblpktETY+q8zxWOuCGeE1WWmVS7OtitWtohvr8mJlOdnRco+QFUZIi1QhMqJeO8Y7ZrHPic1NsUMlQkSI8LWzQVI+fSNWLNEgPJtzxKYIORGVKItcOR+S4+XyfZ7Yajm+QWydJ1ITtcI1Zc76hZXO/A+L7QUf15l18x1n2it59hePhuw5737mLP58nj3/4w3Oks+z5HuVs37BK7G189/0lq1aK4FzX4go9guSIu5NUR7/WsCZZ+zIEsexZxonukS+T3ec6HzHDn3jOLFZxg7Pq446y/6w1Fk1rsh5uSpmPog6ZpEwL+/LeGfIv3AlPst4WgfMVW2C5rdjc62LTmxlXXFhe+tXX4zyHPfOME+723vG/x2Mp1GKY/+tVoUbZeFGTLjaGHxyzhWp5jvPHfVcQtYV0YascMkRzkHGQJrGCdxEO25KKvq2m5oOKnH9jj5cMW70LIhkQyPlz2KXiaEL5RKurF3WMGuZNc3aTiY0dtSPnlcEFAFFQBFQBBQBRUARUAS+UwQ0JdR3Cr92rggoAvsDAiK2PYGc/r/549/v/mj86y+f//NfXseuZ9ndPJeUMggx49DF2XrnrTdeAyYfSr3f3nbnPTfedtc9D/zzL7eS/uaHp59z/oFjjjh60bzZMyslDMHF7tMPxr9x8hnnXfDg829+JL7JyAGHHP4DUk09/dC2qWBw8uLgv+qGP/yZXdhHHnfSqf++/Q83EN2QfC9wFJM333WCb+8+sTt+/uyZ03522a+uXy/iwBKYUHP4MSecfMKpZ56HWPhrL3yb31+mWkYExZk/veTKn0p9yJvrLjn3VFfzgMgQkRDYaixu3yuWLY6TONeL41uiRDacc+Flv/z84/fHf/HJB+9Afjwn+fxJY/XCEw/99283X59I5bLzK6xbzz79Rh869gfTv/7ys4t/ef1N4hsOE0kQ5f8IW5EDfID1t+c2/8Y5TCQC5NG0r76Y6ApBg+eMb776cudH0/QrdmbNEN1DyzObMKali+bPJW3Uxb+4/qYeffoPFJmRzv0HDxuJ9sXXn08gDc6W8sZLzz7xK0l19s+Hn3312UfvvztbQiuu+PXv/4h49F9uuvbK5LpdhQmAZJo/p3E9FVmiiMya2iTHvdvGu6KZctwpPz7n/+645+Hxr77wTBdJ43XGTy6+HDImec2Rco2oDxz8z47/bOoD/7z9lokfvsvO5HjhfkO6Tf7skw8aQtt17iNgXf8817F2EYpH5wJSobqysuKJB+6+s+l3rvGaEnqyBMLnroeefpln9c0Xn32C550reFb4bOh5YU6IgL/8zGMP7eycduZ90hxz/K7bkJ3n/C2MbkU/MXQB4imMxCTFktNL5B1mOMb7su3JqIn42uQHI0sLvXZ5tURcoDMEIYHjGAc3O9pxVhPxwjusUIzET5DBraTFGiItpOFNQlzMEhd5uURcjHHSTZp42CvlSu4n4uoZ/txYvkRdlIi7vMbrjaYKsbEs5vVE/UEnP9XUFYer/SuD3pBcEOvuse18aXe1x9hLhXRY6zeRfsSECPEAcYHmwVghJKpEl6JGSAhSHrWSeu6cs+Ucjvdl8tlVPom2WyzXfyK/DzShqgJn1Qyv8QYqjKiGm4r1EcefErWy2i6RyIp59jt/q3NC1TlWalbYpGZXOmm5U6whJ31qr1tQ6x14bMikpC9wMtu87zgRy1s1PcupnOV1yidVmUA7n127IuypWylppvr47ZqVNdFgh0hNSt/KzMIHhCiYEXlkjWOJLfxRgeU5Nt9aNDAjHpVxht+K48x7YYlgS5rAHmJEt4g8uJkg2hfXfzbSskXIe5VEZFQdNMWGgHBLcgopCAUwd8klNxUUGHHcTf3kkhYQGBATySmlIDlcsW3uPW1CEMbTQjUzWZE0jXj7bIRgPIhw8/05MfQriOohPRgEGtiwHpl3laz1daKTsQ2BmdywflcEFAFFQBFQBBQBRUARUAT2BgSUsNgb7oKOQRFQBL7XCCxeMHf2/Xfd/n9XXP/7PyHkjEjxXX/63XWH/eA4cqSbK3/9+z99MP61l2674VeXusQBZME9kibpuj/cftd/Hn8x7lxdv3b1KsiF5x594D/hJG2Lu2698VrJQtOdyAq0KRB2vuuPN14LOVAf2Mfv+9ffxx574imX/PI3vyfVzL13/On3DTlX2SmOA7yp4sn0d++TL4//yz3/e4Y+ES5++ZnHH3rkP3fenpzCifYQWL7wymt/y1ivv/S803GIu+OUIIS1x5502lmkpFo4d9aM5PF/+PbrL519wVe/wElNO++/+fILt15/1cV8J7ICsoL6Iw8aM3Z3FtTAYSNGQzj0Hzx8ZF+JAAhKHis3uqOp7aIvcMJBg7oxd6INSBN079//+PumXr8r9XZmzXB/IZoaSrVUv28c3zdc8bMzISHY4c86vP8ff7nlkXvuvL1+3ecevf8/h0pEDYQPxnk0U3514Zkn1ScEuiWiYSCfGpsvJB6kT0NrGdIB5/qJp599PkYbaGtcf9n5P4YYdNuUDErreV5Yc19++tF707+e9Hlyf8Ivef952++vb2ytQxgQGdOQXgbHnxaNiPMv/eWvBw0beQDE3Q1X/PTMspKNpGzZ7cKav+za390C7hBEt9907RXfPiubo3XOPP/iK+oTR6ReQ5Qb4rKhQbRq0wanpmmILNqZ98luT/A7bCCRIgfndK4YTnCICtLnUHDw9sIXLc77EaJXPT7mzY5lln9S2mrTI+ne2CYICTAcKIYjm533tDVSrCRxfWv5xJmMAHdQrEjczBNk//8GcTN7xU0+UtziAdIiOWmmu+WXI3RHpTP2nAAAIABJREFU3IXf5Ppa2yvsKusdK8Xu6jMiZJEtPvR0M9sbiq7xVMe6WXVOrrSX6vXE6iS1lEQumJkStdGTNoRsIAqNvklVFY8oEJKiq3y6kSBoIECysE4ZL+PH6Q9x006uny+fRBT1EGbMsnLa892RVE8+k54XtPK7pEt0RYqJhiF5Wjs1ZaQnwmnuOIs+xYm+Pjb5kToRGjei1RHzjY5HImQ5jgdyRvQ6SDvl8TiOZZvKL+ssx3KENbByjBNLkQnH+9ps1mvFji0WmTTKQ0o2ogkYJ8545ogGDvPi3zrw9ksEBuf6ClkB6fCqXMdcS8VR76S8Ar+0JfLCJSTcvlyNCEgI/vsISx4L80q+Jpmc2Op4CxIVjN8tECncPwgxIiiI9GD9UWTtbiljE7+Zz0RZ92AVBo/kxvS7IqAIKAKKgCKgCCgCioAisDchEE8fokURUAQUAUWg5REgmoBc/ggII2p95wNPvjhSSIa//v66K196+tEHGxpBxy7deojYdD9St0jqpFk4jxsbKTnpcew2lAIm+RoiAPLyC1pXSKRDMvGRXIfoCKIXGnIUN9Y/aa0GDBk+ijQ2OEIb2hXPtTihSTMkaX6W1Y/sIOXV+Zf98te333jN5Y0JKue1KmgN2QIp4o4FguGoE3/0405du/f8TBzZkES7c0fRDoB0cNuAsBC9hDT5/7QUhBNEDRl9EX5DaEjWoQAployMo04mvkAc1+74OX7ymeddQMqhphJAuzP2pqwZSB0iBppCWCRjzLrZkdA195conjaiNk+6omkiXN6Q1gXRFehHQDK4kSj1581zAmGwPVHrfoOGjmjVuk1bCJjGBMRZb5Kext6Z+bpjYV1zyxvSinDrILwtt9nfUBTG7txLruWdkS8TTCb23DaJLpk3a/o3jb0/Guub9d1eCL7GtEO4rqnvk92d33dxfYKswIlO6hwiJUiTdIMYO/Zx6ktBSFt0HJzQXEkB9VRB2UOrsqrG9/U4tVxHtBcO8ovEcGTj9EcDAyfwO2K8p4eJdRVDz0I4APNPcX+3kjN1QkmsEZLhTPnNDvhWIsa9OWVURCIzIiSMMuvl99NOuVlpZZqD7Ih1iNT3iVh3hcRdLI6tNAdbIcd2aqS2I475oPnIqRLndVTIl1h8XDiyh4vhzIaMICpgiRiaDJAzpA4ihRCRVpAuru4MUQIQiMsT44eQSLNyOxR6Rp4Vttr27WnSJBVZbXmVs2ZOaezje6dK5AXEQbnYV2I4zekLcmGupL+q8w41EU/nODakyuIc2BDVgAMdUsFN3YQDnv6JZKqzjopjuaXIPUv+yXf+G4b+SF+IoPfRYpCkpLviHkG6LBTDQc/nInHSu4LY8baEwHD/O8hNI+UKVCdHYriEBveZsbp1aCKZ0OD3ljG3BGnRAAb0CY7gy70iNRTRJ6zprvFJCnkkxv24Q4x/M1mrRPLUKWmRQEg/FAFFQBFQBBQBRUARUAT2OgSUsNjrbokOSBFQBL7vCAwUoeG/3//EC+y6Xy7ZlE47chROMi2KgCKgCCgCewCBBGGBU5foCpz1PxW7Tox0OYnoY+dDj117l8euCrQtvbMir/wZS77jaMfBj2OaqIKTxdqLuZEKs+R7oRh/Xx8jBvmBxgUaLI/LVWPifUqkhbjqj5ff/cQq4kSDFa8Xc6ISiRESIeWAON5jptYKmlFyLF/iIWJCqwRF3vk9e6U5V9ooEKJjkpAa+fLdL2dxQq9z6qS9mEQfOOZI+U3UBymBcOhDVqwSi6dZk0KEDjvzOQeRQGQB88cp7wpXE3HSXdI/WZ6DfhbwDD81VUiLNFNZXCuERUnso7tfdtbOxQHOjn6Ep2EViLRYIfOZKQRLkXegCXu6xIkFnOoY2OD8B8tkrQn6ZYybhKzYot2SGGv8oxGHPacgPiApIInimjPxMRizQIx5YeX1CYvkthPRFw39d1E80iNR1/3uEhwcjpMULUFQJI9vB/NnzXKvIC3AEfLtqMT17ppGQ+hJMTCGxClRwqI+wvpbEVAEFAFFQBFQBBQBRWBvQUBTQu0td0LHoQgoAvsFAojxXnvzn+98/81Xx6F/MK8Josf7BTA6SUVAEVAE9hwCOJyJROgjhlPfJY23/F0s2hVrciuen+yPru+SWf1JF8upJRUR1+Dgh+wgOgJHPw56HONEJnAMooDiOuhxIBPpcKa4vbk2U9zr6XH9hc0kRa78xoEM2dFKUkNtkBFVyrE0cT1L5iQz1PKaFaI0sVpohJ7i+u8jrv4F4oLPtrKE3IhIyiefEBS1pkzIir5CBayT63BK48CnfcgH5gVpQD/x9ExiEDU48iEc2ojheId0wPnPvCA3KHLOiTmrZ9pOx8HdPP2OCprWPVNNRr7PU77uB7G3/zzJxCKdEnXBgqgDyJBMGVu5zMDVdqAKznOXrAAXjP7c9Epx8WtHYj+EtNimiIN924Obj9hCZjDnL8TQCmK+ECK0x31gDNtNgZQgHBqr46aToi+3zh5PqeTOvwHiBvyIckGzhLxX5yYB5a5p1njfBBZEnMRTeDUGqB5XBBQBRUARUAQUAUVAEVAEvksElLD4LtHXvhUBRWC/QQAdg1vvuu9RhHP/dfvNvxn3xCP3fbFwbeW4Jx++b78BQSeqCCgCisB3jEBSOig0b4aKkfotLm7wbZE8S3bVa6JXEfDFSjwisp1iOTaRFBASOIdx9rsC26Sfw+l+ghgedQznOQ5zUk1BEEAIEAEBCYCeBdoStEGdgPxmDOyQJ41Rrrj0IT3Widt9nbiUU6T1Lla6kAkSVSHHOwlRsUnSQeWLRsQYZ5NcH4kfZw5B0cRoL4IQnwg1UCH1IVbog7FS0LUoFCP9kktKEImAWDNjJRqD1E0QHZArnSS6IuzpfbjjOfKXOaa6NOxUbIhaKZkeSROVarXqlmF1GJTqrJyGoxxiAFJkc9SE/K/odEeld/AiYiLNti1vJOoVKC27to5hWSbgj0ZSU8OOKFqAAQRKo2kPE3No8COJzKB/5ueKZdPmbpd6ERR7m6Of8YAx6w68XxG7oN6kWR/dxViPYF0oz0KtRlns9tLQBhQBRUARUAQUAUVAEVAEWgABJSxaAFRtUhFQBBSBZAQ6d+vR6+5HX3iDXPSXn3vK0VO+nPgJeffRNiD/vKKlCCgCioAisMcQILoCsgAHO15zhMyJkNhSLCd8tS+6scyx/Gm+WLFPPOxyzkF4GmIAZz6pj4hGcKMXcPZzHMNxTLuQGHxnJzt9oh9AFIWrvcD1kAI4+SEWMJzKlVsiMSARLDNFjrWRFjeKK5oUUo6njcl1aiV9VLmpEqVq0ZQQ57xlVgl50Ufc/QWWR/r1mHdEhPtHUt/tl7EcIAYxMkOMSUFQ0Ce78xERRw+CSBEc2mhJ1AjrMMgRuQwru22ByW5jnOVfVTgZraqszIJaq++ROV6vf2Ps5RvecUpXQdi41y2T8RRa2VxvnA8mDPAVbczMtG3PgPTUUFE05m0VCvl+7vfHgl6vva51q4r7e/XYUJWaEqnOzane28gAmdbeVRqINHGEfCB6hULEECnKfil2T9LIue9ofDwixtrnGeB+Kd571+3V0SgCioAioAgoAoqAIqAICAJKWOgyUAQUAUWgBRHo1rNPv4fHvfVxbW1tzfknH3mgCE2Ty9wMGXnAwQhoL5gzc3oLdq9NNyMCIpgdz2Muutr7rYNHMIhD0JCTS3BpRrS1KUWg+RFIRFe4KYmIcvi5GKQBRIRbSCu0WMS16yQtVMhyoghUI1xMRAJi1ERQ4ORHL4Hvo8UgKojYgMAgxRK7+nEQQ0ogeIwTGT0LCAOOUSA9IAcgEuifCA4ErNHV4O9zHjaEsUnjRMTFQHnyGHuRnM2TFkPyuchqZUY7G43jVJtUSSeV5niFyAjJWSfeHmLeafKddEATxCaKnSE2UgwiAwwKxRgz0R/MAfIFhzdpniAy0q3cjtkmmJFmgukBs2FJheX1G4msQC/BWAOPPdVZPjkW++ietkJu0BZzJbrBlh6CM6Z39qyvyu4v0RWnOMY6paIyNSoTi+toxGw4HQF1RcGhy1YUvOL3xe79yZmTGMd++46NA7JrxcUMIoo1hsg6a/mQRHPop1BY8whwc84rz4SjURa7BrhepQgoAoqAIqAIKAKKgCLQcghs/i8FLYqAIqAIKALNjkBqWlr63Y+98AYe7svPPukol6ygo+GjDx6zaP6cWXVCZDR7x9pgSyGAR95KOO1bqo+9ul0lJfbq26OD2zECrrYBjvkLxSAr6hV7npAUda02PbwuJTQP3QoEpTsnDA0LHPoniR0mhsAzxIRLVuBsR7/hZbH3Et/RDYCsoC9XKwMigIJzGWIBJz8EBoQEf5u7QskQC/SzWWPCMnPF0IUIWQFTZqXJTvmYEAoB4xdx7nSJaKgUC3nammoRvK6WeiXS2myxpfKduW8mPDb3Rx/0SdtEV8wVI4oEIoMxQMbkCRXitee864l9+O8iSQklVERtjbNh0dfynRRXsk8/t6/nqGsvsXocJMLhHtJJkdJJyAvTPRLyppdXp2ZEY54rJUbjLOE7+yXICua9pcgxSbVl/UbSRd0x7rVR4Ktl1xHgvi4Tc8my+i2xDln7rFkigXTz2q5jrVcqAoqAIqAIKAKKgCKgCLQQAvpHagsBq80qAoqAIvCzy6/+Taeu3Xtec9HZp6xZtYKdufHi8Xq9B4w54qh3Xhv3rKK0zyHAv5uuWOw+N/jdHfD+TNbsLnZ6/XeLgOwkxwmPMxyC4RSxnvVGRJok0aqIfZVZM7Ewp/K1oOVEIBogDXjm2cFOJASOYJz5vNN5H+D8hwSA0MQZjMP4QDGc/+hDQAgQjcDxOWLsfIewYMc7RAgkAroCEAWk6HG1LSA+iNRYLAaxwFjoBZIkXSiFkOhaWPJ/k+RXLytmKpxKGYs/Hu0xSPQtlsXKJeLDkv490kdMPp34nElBxTjph/F1FCOaAmwwIjogaogW+UqsytSU9Talq/zGF/BZA4/rIN9jTtHSTVa3PMZvrPwubX0XPDoq9vzVq4XcIIWV3zaW/bXdM6PQLrhTxnBqfOybg7PA72kJyJrrsZx0ITIgS86U45BBVk1tcLh8TthcX8suIMA6ZSMEwtqTxVhnrCv0WtzCOuAZILpnjTwbmyTKYisSaRf61UsUAUVAEVAEFAFFQBFQBBSBZkNACYtmg1IbUgQUAUVgawROPP2c8wuXLFrw6Qfj30g+M/LAQw/Pys7JnfTpR+zA1bLvIIDDkx2plF0Sht13prrDkTaYFmqHV30PKiRSg7nz35K6RqNP9o6bK87XhgbC/SKlE05/Ujgdk/Qsu/XRl/jca2+an1X1tu2xK3Da90lcB5ngRj2Q7ohIAt4F08TQAyCNU1xYWoyd66RaIt0TxASOeAgOUkshqo1WBVETrB2IA/QzID0gLiATqsQgQHA6k3YKoWT+Xof4IHUTc4nJ/46XKyokkmKYjCxNJKs7QGIg1C0pogJOiels+URkWyIrnFh8vLRPfxAS6FPQDoSDq2EB0cGYXA0LrtlM6tixRSY102PqKrsZXzDorF9YZc97f533jLvyJV0UBJCx2vRu7z3vv6c4/zx6qlO8rDZk/Hkr7fwfS1jIqbQqBMUHlnEWi4L5FJ/X/jolJVI69tAFJRuKss30WZ3vDEd8l0q9mGTe6/voM2M+N+YzV5MhPgQtO4WAK3QOQfZPsUPFkgkL1i7PAOTZJLFaeW4a1LNoQC9jpwailRUBRUARUAQUAUVAEVAEFIFdQUAJi11BTa9RBBQBRWAHCCCo3aFTl24fvv3aS/WrnnrOzy6prampnvzZBPKTa9kHEBAnNWRFPCWUmF9+R/ZHLQuc8jJ3nJr7s2AFc3dTaoLF/k5e7QNPcHy9EsWAc32IGLv465eJolsxKxBZU5pR85nUt3D6oikByYFjn98QExAIkBScIwKCv6WJEoBM4DgEBOtC0hzF18ZUMYgP+qc+kQs4iSEnjhaDGIEEIXoD8oCd8URkEPXAcYgGnPdcC5FBhAJjypVVSNREutT42koVwiQoOhaVJt2uNn0lbmGjXSbkR1jq1cXXK2PBKc31r4uRqqq32Ddi74qdnDiGM5s6RF4wRoiWmfb8j3sYy7vOBFLTrLQ8j2fMJR1cskLOx4vVqntHz0E/HR1767aJpbEMT9R4f+iek7fGXK/XeSjgj5WGwr7B4Upf5y+/6jkhK7MuJmRFV9JFSQsL5ZP+2/3vwjHgDWmz6eLHPlNNCxfIRj4hFuqRddxr7h33HSx/Wu9SngGeBVJ7UY/1pTjvAGc9rQgoAoqAIqAIKAKKgCKwZxBQwmLP4Ky9KAKKwH6GQCwWjYZDdXVEUiRPvd+gIcOP+eGpZ77y3BOPhETAYj+DZV+eLo4czI2wwLmjO4D35Tu662N3CRt2xeMIxqmqpMWu47knrsTpD6mA6PX5DXUoZMVcX3RDUV75E+FgZDnRDERFcH8hIUiVxLPPvXcjEiAaSBdFXd4FnOe9wHEiKSAccBq/InawGCQE/x4QuUDEhghCxCMr+FsckWvO0QbkCMdZV0RDEDJCm9TjWr4zJqIl5gsV014IiwPE1gnLssnBNR0zQScqhIktehq2yRQxbsuxzBQZZSf53U5mARkBHvRJyiCEmYkMYS70CV6Mj8K/Uz0kLVSxidYt9Bx60VhPl5FdTUY+BIz0FQkZr5/oFYkxKS3yDD6xlf3NuA2RNcWwRKEkD/h8Sf9UWxfydxdSIlciKQYXbczqI4aGx9lizPsjsf+IcYw2SVnF/PX5StyMJn4AO2QX95AVMbuR63gWIMFIX0Zkj6aFaiLAWk0RUAQUAUVAEVAEFAFFoGURUMKiZfHV1hUBRWA/RYBd6J9//P74w44+/qThBxxy2LxZ075BaPvWf9z3aCQSDj/xwN137qfQ7KvTdiMKcCRS3B32++p8dNy7hwDOVNL/UHAM4ujT3cm7h+luX91IOihXuwIHP+mgcPrXL9Msu9ZJDc21sqrfd8kAHPI4cTEc+ERUcK8hG4iGYA1ASvBOILqClErsVsfxDvHAcVIqXZG4Bqc7kRb0T6oo2uG9QhQD17g6GbRLeip2vRMFAYngtodjGVKESBEIBzQmhI6QOnbcotJKraxMn8RbBOR/WxPPYRWI07/S9HIqZNzU29wn/UOskLKK3+vFIAfoHyIDsmCJCGlnm5TMkNV5WJrniF/kePofTb/fFggLO+aYaDjsrJ07yeo6aqj3zH8dFL3n59844XjbbnnQti30OLgfRJ/UL6TUghxxU24xV46pE70BsJp4iGgeyDQwJH1Z/cgi1iLPxMTE/YeM2wpvnilNC9VEtLWaIqAIKAKKgCKgCCgCikCzIaCERbNBqQ0pAoqAIrA1AnfeeuM1fQcNHf6/l9751D1jS/nj9VddvHrF8qWK1z6FAM5oNzULA99vUyIltBr2Z+c8c9+8j33zLncKmgD7MyZ788OMgxzj+T08MVAiGiAdKDjIP/I44Uhq3YwKX7QYogIHPpEGRFZwHiICRz8kFe1AIGCQGZAVfCe1Ejva0a+AyOA4zn/qrBbjb26IAEgL6rOzHQc+RAfRHFxLRAbjYgyka+IaxoIjH6KiqxhkB+OhDfr6Ot6+FderaCdi28bTydSIjsVGJ00iGYqMI8fynRqTZgVMrUQ3rJSV65PVShtfiF0txjxxbkNSQLTg5PYaf+p6q+vIoGfkGcO8h112iohub46kSCrOqplvGn8w3WS27mt1HCIC355UT+8xF7U66LSJ1qdT58lD0T+peq/61yd+4ygfL/asGLoKYFcuqaA0sqIRwJp4mPsICcW9JXplUGLdcLn7DPBM/EvMfU6UIGoiuFpNEVAEFAFFQBFQBBQBRaDlEFDCouWw1ZYVAUVgP0dgw7o1q88+9pBhaFb0E+KivKy05I0Xn358/uyZ7HTUsg8hgF6FFJxnpGnh306clvttSQhPM//9TnQ6oePBWnB1TTQ12N77JLgRDDjNzxODGKC4ZAXfZ1hO+CshKza2LrvX43HqIA0goiAW5onhwMdcDQsiLQrFXI0AIjKIJIC0Ygc7KZt4P0wRI0pirRiOfvomqoF3CA5kiBDOcxwHPdEEkBMQEawpHMoQCVxDtAFzILqBY6vE+HeEVFNoaoSFrKgRKxGrkJHOk9W5Sd5UY5yIsZ11QobEJCWVpIeS44vkO+ODfHFTXzEn5si6XiFRFUVWRqsMz6gzTxBNCp9ETZwpx7cpTtHiz40d/dTUhR170cSp3sOvuMrEomVCdHQqOOOWE7xfnv63aCTyD7kwGW/mjbn/DQKhIyLb5r/MSUgKcNXSPAjwfgZPomcmi80QG5Vo2r0nrD+ejSfFpotxP5R8bR78tRVFQBFQBBQBRUARUAQUgV1EQAmLXQROL1MEFAFFoCkIVFVWlD/10D04bLTs+wgkO6lttKcT0Qb7/sx2cgb7o+B4PYhcEeQNchwHtDr4dnIN7aHq/J2LQx/y4cBEn0QrQAy45RuvXbk8t/LlkMeuhnzAgQvpQDQA5AC/SZ1DlATEAtEPECG8D4aKQVxBSHQVwzkMmQD5QFtcBxlAfY69KMaYaBPCARKEdFDUoTA2+qBN6rE7nkiID8SOTPRHW/kJK5TPw8RYj6vlqo2yEh2hA+Y4IfleJ0RBnbQdMLaIcluSEsqWkTBWtw2uJXLDTcO0yXh8IavT4M6eXmM6eE+/Y6hEVWxLzoaqC52Ny6aZaGSdvWpm1Jn99mIhNoTrKZ9mpea0FhJjquULVnTs1uvdwkXzwP8kMdJjQYqAA22Shgjn+Eyx98TmKlmRWAW7+OGmbqqXGo13E6QXUZ1EAbmEBb24zwLPBunFiN6BpGM9bCmaFmoXb4hepggoAoqAIqAIKAKKgCKwywgoYbHL0OmFioAioAgoAvshAm4+cHVQ74c3P2nK3H+ICooryL5/I7J3zh4HOWmY2MF/W2KIyWTFh5YTe0OiK1ZnVpMxJx7dAMngalW4zzuOXJy7RDjQJg7/tmIQDcuSrkHcGAFr2nAjsnDK8xuSAdFvN1UU6ZcgI4aIIcjNOiK9E+QKpAL98Em0x7BE3xAYRHMwp+PE6A9ihHEzliohLeYKpVItva8TWmCKxFFke9pKuijbxJxak2LZprXjkXRXdnw+ZdIrBAJ2mPF40z2Dju/kPf7G0VaPg5lf/eKYmk3/jX3x2CPG6+vm6fuD7t4Dz/uRM/y0r01d5XTLG3hfUkLliZ7F105dxVc/+N2DG/934ZjbpZFnxCCAfiE2Qgxcl4vdIxYXfBayQlMRNQB4Mx2ClGK9vZ64D0cl2nWfBdYYzwgRN6y7rQiLZhqDNqMIKAKKgCKgCCgCioAioAg0GQElLJoMlVZUBBQBRUAR2J8RSKSFcrUsXNFtzbG+ny0KImukuDoWSlbsJfe/AcFtSAV28hPNgJMfZ2xymSo/PrRMuCS99qsKSQtF5AR6EjjqcdqyG520TKR0QiQaRuNsMYiBCWLsSucaHL0QCKSDWiA2VgySAu0iIjBI+4RWBWmVuIb0PB3FLhB7TAwnMg5iN7UYTmTW1SIxtDAYD6QI0R6MBd0KiBNIBqIzuJb3EQQa5EVQtCpiQht0Et0Kn6eDaW/5zSC7KE58eBxbIje8Zp0c+1yS3K2TXr0SVXGolZYXtAYeN8R3zn+6mtTsraMqHDvilKy8O7z4ixXFE57+IrhsYnUgp83UzNHndrJSsoJi6U4sMif61KUf+i4bFzMBn/EE0+PvRiEimNcSIS4gZxAL75KYHym0ljcUVSF1wZ/7BpGhKaIAcicKkRYNRFmwJsH8QzHWK8SRW3g20LcAa+49z46S8juBuVZVBBQBRUARUAQUAUVAEWheBJSwaF48tTVFQBFQBBSB7zcCOHJcDYsouhb7a1qo7/dt3u7skp156tTbexcCTnwc+KR3uquBYb4i0RUzjGOz+9x47QpXowJioL2YqztBrn/SGuHMRRyaT5zpOH2py3lICKIw+I0OAMcgF3DQk46nUAwRb6Ir0LaAGIF0gAjhGMa1XcWIomBMr4mRSulQsZGJfjlOaioEuSEoIF3QtiBaYq7YgeJqtsTlPMTKkRiLLBOzwjK1tSJk7UgaLEuOOKbK09q851RK7EWtjCMYWOXpNqaL99S/dLe6jWbeW5dwTa2zZs7tlQu+fGbD+HtbF9eYwbWmc6yqNCUcuPsmZ8RZvwym57XuHQ1bXafZ/dYcaVmNkbg8KxBAjBvsSJ2Flke8CEnBcwXmzI05ce+K5Pj7QlrE75F8d1NlEVHiam5A3MSkzjZD358PuOmhEhg4CQIDHFmfkBLJhAXV7hO7PoF7HNP9GT+duyKgCCgCioAioAgoAorAd4uAEhbfLf7auyKgCCgCisA+hEAiyoIdzTjXKDjQNJXJPnQPd3eoSfodSlbsLpgtez1/45KKiZRLCEzXL7mWU1OYVjejJLfiBZzfREtAROAMhzzgN0QFTnYc+RyDLKDdgWKQDrR/vBgaE0RRcM18MZzy7FrnPUEdyidiXRNtstud86PFICggNYi6WChGZAXncNqj+8DYIUomJNqFmLhKjEgPyBg+WYtELvA9S3rtJbOYLemf5ssbqsAKin5FwITlM1Pc/Gustt6gE/Z2t7J79xO9ism+M+85y6TnQSJsKc7yrzY4xctWO8u/ftWe/uo7KSUrIvkmxS4zbdeWm+x0j3HWbli+6IjZ7zyb3bbP0B7rFsy4a/3CGS8JqYC4MwQKJA4kjavxwjxIC8U7E9IHgif+Hk1EVDBX0mmBCY51rgODCjmPzgXv2WRCBUKDe0Ndda4n37yGv4MfJBF4Hd1AFe4PzwpaFqWK6Y4B1RqKgCKgCCgCioAioAgoAi2HgBIWLYettqwIKAKKgCLw/USAFCc4CHG8KWHx/bzHOqt9GwEc4UQwnCZ2shhpliAaISMoUy0Tmxy8MoLYAAAgAElEQVSIrC5uX3yzFYwsJyICZzgRDzzT1IeggEhwneE40DEcvkQCsAvd/U09HML8JmqA9EcQFehR0OfhYrPESOHk6ltwDWmaXOcwYyD1E2PAac97hr/TcexDYNAfBR0MSA4c9hAZ1GO+kCUQLyH5FZA3VIVTbubI7+6SGioqIwsbjxWRZFGpTnjIMd6jzhtg9RzbyaTnX5BMVjilK8vsD/75nrNqpmOvnrnM1FbMNXYMTAIZpi5/qKdwYcCJVhQ5WYEyO1a5cuaXlZvWrWxjeTx9HDt2g9SDdGFuOMchGiBqwJN5kxILxzj6FYw7XcgISKGDxdzoCogg7hX4U/ccMbBlrqQtggwhtVH8fqS172n3vfxuj3ksS4ljAaSxIhEXtkRZsIaKxCaJEZ3jRlmAN/eIZwVs0RxB80JJ2e1gqqcUAUVAEVAEFAFFQBFQBFoOASUsWg5bbVkRUAQUAUXge4gAKaAkFZTrHFMn2ffwHuuU9mkEcN7jfEXrgUgIHOIUl6wgJdPj8hCXCFHhCURWupEYRCvgaMdJDknBJ8QD1+GwJwKCujPEcJq/JUa6JoiGUWI4g9GjgEjgeogICuNwxbNdLQqcwuhdEBWBY5jrcQ5DOLjC30RhIKoNATBGjEgOhLtx9JNuirGhj3GYGOQMbS8RI1LCI6TFJhltUFz9jpVu2js1wjd4uno8HQ4Z4Dnk8tZW11Gi6+EGiknnK6eX27PHlzqFU5ZKdEWtU1FEuiwiTnBqQzYw3jiJ0t9aHepvmeqXYgfeFbL9J1ZtXHdQZusOY3zB1NxouK5c3o8bpN4RYoiFnyvGfHGKQ8aAK8QN0RN8DhbjPQrRAyHBJ/MgOoOIEe4lmDIvMKJt5loqaaCk7mdm+uV3e8UZ3yh5XC89kly63xZwBkNSkD2awJ215z4bPCs8M6xZiA3WuZIW++1y0YkrAoqAIqAIKAKKgCLw3SGghMV3h732rAgoAorAXoVAxy7deqxesXzpnhhUWnp6RiQs/xcJb8lhvif6bcY+kkWX4822bd+xU0lx0YZ9eE7NCI82pQh8Zwi4YtsQAezKp+As529ezsWJCY9Tsyqz5pNKX6wEkoC6OGhxzOP8d9MPkZ4JUoH3FM77rmKQD0QNzBODsEBzgX4gLAaIfSmGo56+aJP+0AwgIgAHPGMhtRSf9IfTnuM46Z8SQ/eC45AR74oRYQB5wVhIqcS7B6c/Y+onhjOf7zj0idjgOgiTblam6eaEPBGTk+31dBibb/W/ro1JaZ1ute6NCPm3JRqKxD57eI4z802JylgvJEeUaBMIERzbOLHBBKKAdFREmDB258feycVPx8Y8FYtGvoiFQ8W2HSWCgugPxgGRwydjARcwIgoEAgIHOQQMZAxOceYDgQG2RGYgZM494BjEBfcHDEgBxVzjRLFEZyDqbYSQiAlhAd4qFg0wjZSkKAvuLeuOtUlhTUFGcV+4T+Ct4tvbwVJPKQKKgCKgCCgCioAioAi0LAJKWLQsvtq6IqAIKAL7BAKDho084Mk3Pp581rGHDF00bzZpPFq0/P2+J15o1bpNu3OOHzO8RTtqocYTQttbdp76fH7/Sx99Pfe+u277w7P/u//uhrq95ve33TFo+KgDLz79OHZEa1EEFIGWQQACAkf+QWKXJ7pwd5DzMyzpoGzLCW9oVfYgju9kJzfOWhz/OGtxtOOcx5GL4WjHaY+zvqsYEQSdaE+MyAxSN/Eb4gLiF9KC63G4MyYiAHDOQ1aQ4mlNok3Ocz3joJ9vxHAo47wnqoMd7/SBcR1RCNSlL7QgXMIC0oNxM775xvK0N/6CNqbtaROtsqJqkzmom9VmQIEJ5pJyaUuRyIrlsY/+86kz7/1CZ9NaCAHOtxXjvxEgNhgT8yCyBNKAedA/+Dg/8X7G+UVPbxzzf8H0rHSJruA69Ch+KwbJw1zQpgA/frtY8J25gRfznyAG2cE8EYYmQgViiGPVQkxsN5pNnPEaCSBA7agkyB2INO6fu2GA++k+IzwzRNOQNoo0ZqwxLYqAIqAIKAKKgCKgCCgCisAeRUAJiz0Kt3amCCgCisDeicCIAw8lx7qpqijH6dbiBYJk5fKliNTus0Ucc1vyqch8hqVnZGRWVVQ0it/Bh//g2OqqKhxzWhQBRaBlEOCZxNGPBsR5jXTxmnGi67KrxifvyGenOZESOOsRHib1EkQCTvPjxCAK+JsZ5zyOXhzyXF+YqMN1XEPfOOdxyrvkBSQHznQc8x+KQQIQtYFGA1EI9DEtcT3tXpioT5/0BUngRmFARiRHR9AuRAB1JO2SxzH+vIWm4EfVpnZJlWl77ggr/8SbjBNzjG23TyYrnPXzN9hz33/X/uS+RU5JocfEopApjIc5MmbaxaGNw5pP5ug6uSEP6hMIsVB1BeQChbRbpIJirIwdBzlprWgDwoNxgzntEbUxQex5MVeTIyIEhRIQCTBb4APcicR5TQxyr37h2aEOETCQVXovWuAmaJOKgCKgCCgCioAioAgoAo0joISFrg5FQBFQBBQBM1AIhNKNxUVrV68sbGk4Ctq0a5+dm5c/59VxCHvus0WiLISzcOLON/BjIrOnf/NVQxPy+wOBbr369Hv9hacf22cnrANXBPZ+BHge2bkPmcDu/fplvkRXLPJHNyxPr/mcaAR3Vzl/DyOQTeoj0jHhWHc1KPiEaMQZ7zrcEY1GR4LjpGmCXCCVEc590iDh4CUFFE5hnPekdSJyA1IEc9NEERXhRngw7lMS10J8oPdA324qJeqx8x0SgPPzN9exWhlPSqpJ6UgaJ9ukDzrLZA7xmYKTl5nMEQeaYHuiJWREkYikeooaj8/nLP98bmz8Lc+bklVfO6XLq000SrQI86BdMFwvRrQF44OsIP0VpAgGobFNtAOpmZIK88fRDSarJHUTWhzgDXlB+xiEDQQv7YEVkSIlm3UptLQwAtw/UpBxP1hH9UkLnh3WG2uSe+4Kz7fwsLR5RUARUAQUAUVAEVAEFAFFYDMCSljoSlAEFAFFQBEwA4eOGN2Ys7254endfyA7mM282dOnNnfbe7o9IS1sIi0GDh05uqqyorxw6SIcituUHn36DSBt1NJF89lNrEURUARaBgEICJzsOFiJEKhfFjvGyvE4df6U8CKctmgn4JglOgKHOlEVkAw474mCIH0bTnfqor+AYx1SEicvpa8YaZsgLogioA3aJCUU1+CEh8zgE20KxoejnnqchxyBaEDjgQgH0icxhpGJdiAQ3JRP9A1JgpM531j+dcaXmWcCbdJNev+ASeuXYwIFIZPaPcVkDm1jgh3Hbh5iolh+vyn5/Et70YSFzqo5a0zdos+ckvW2kBWu4DfjJh0g/20AfoyR9FWFYpAXjIN57pTzWsgK7gN9gCUYEn3C3BHifiPRJ0QPOFVIfUgLSAwtLYcA99AVmyfSsT5hwT2jDs8Sa3an7nnLDVtbVgQUAUVAEVAEFAFFQBHYXxBQwmJ/udM6T0VAEVAEGkGgVeu27dq069DxpacefWBPgNR34BByu5u5M6ax83ifL0RavPbptNFzZ0ydQshFQxPq03/QUI4vWTCPncZaFAFFoPkRgHjAIU60EynuSJ+UrF1Bj5967NqP/dG15b5YMbv8cZLjnMUZj+OWyAcIAaIYOA6BgGN9mRhEg9veCfIdJz6OdpzrkBUQG6SBoi13LJAZEB8u2UH0BcQDkRNEaTBO2qQdRLUR7OZdAWlB++743FRyHYzlSzW+7HRJ/XSocZxakzEkajIGBuRYlsk9KsWk96WPbcv6Z94whXe/ZQrXLbJnl8SMU7tCaIOgjPQ9iQdhJz3kiauzQb8IL5OqiqgSHNdgAaZuhMUO0wQlyAoiS04VY1wQFa4mxrPy/WExSBGIGdqrE7JCneMN3sBmPQjWRO58JAYxdXK91rnPrE03SkjTQjUr/NqYIqAIKAKKgCKgCCgCisCOEFDCYkcI6XlFQBFQBL7nCAwWIWimOHtGw+mMmnv6/QYOGY6Ww4pli8mPvc+X7JzcvM7devT64O1XX2xsMv0GDx3BucUL5iphsc/fcZ3AXooAznYIByK42MVPNBMREJAFbgk5lq8ms+qDqkBkFXVw1uK8hTQYLIajHqc6DlpSQOFs7y5WIkYEApEXkBL8/QzhCvEA2UAfXcXQgOB3t8R3HPH8diOrjk60Qx+IglMfogCyhPFQv78YRAeaF9QjAmOtsbyLTVrfTcYT7GZyj3SMNy3FhDdUCWGRb1K6EFWRI+mf6hM0QqPcc6ep+GqFKf3ANpHS+Z6c6Eanvam215hqJyJ0hcRYJMboRncgBg5B4qbEgrBh/pAoOLIZ03bJCiEqIGwgfIaLudEV7thwlKORQTTaqkQ0Be1q2UMIiPC2PX1VBameiOphrScX1iv3hvXIszQxsR6USNpD90e7UQQUAUVAEVAEFAFFQBHQlFC6BhQBRUAR2O8RQH+ByAAiBPYEGH0HDR2+cO7M6baUPdFfS/cxQNJpSZSFNacR/Qr67z9o2IjiDevWbiotwfmnRRFQBJofAZzkOGBJm/QjMZz+7sYcnPHviQU8Tqikddk9OGl5/+CcJSLCFcEmqgBHO0QG5xDB5pllJ/qgRJtEWuDMx4FL1ABt0ZcbbcFnoRiEByQHbRycGAvX4uyHqHDT7hCdAeEByUH/aDgQ4cH4cPL7RKPCMtkHRUybM/ubSEnIeNPDJlKWYlI6p5h2P2sn5MXWG5Ds2mpTPf9hs+jqL031PKEkKkpEaBwyBEqk1tNBCIuVMu5YfJ44piF7ZiXmxPggWCBMmANzdZ3aTXVa0yaEzPFipLviOvQqSJXFJ3P/sRjO8ML4uLTsUQSEtIgIaQERxb0i0uVYMaKLWItoWECkEfHDM8WzpUURUAQUAUVAEVAEFAFFQBHYYwhohMUeg1o7UgQUAUVg70RgyIjRBxUuWbQADYaWHiHRCB06den28btvvtrSfe2p9sGPvhrTAPH6fD50O77+YuLHe2pM2o8i8H1GQByt9aeHwx1yAKFqBKS71qsAKQFpMdsfWYsjHgcs9Ul3hIMepyyOeZz2ONiJqqBARBBRQeQFO9Jx5CPOTV3aIPqB1E2QCwyK6ARIABzyvE+pS1ukXCJqgbRPOO8hIuif8xAVaGjgzGcs7G4nsgNSY6NoURSZ/GPaC1ExxMTqMo0VqBEx7c7Gk+oxvqzO25AVS29aaErem2XqCguFqOguRAXjoG8iJLAiK1vGG4iPw9WqoF+XSMCBDekCccJx6rgRFU1JAwUpc5bYWDEwwfFNFAeE0WNiR4mdL+aJOdYJV5zywye/LsmhPwr3kUI/mBvN4Uz9/OnEKf1oRgR4Foj64/nA3MJ/H3YV41maJFadiMjYapOBkB7NOBRtShFQBBQBRUARUAQUAUVAEdj6D1LFQxFQBBQBRWA/RcDj9Xr7Dx4+8v23Xhm3JyAguoJ+vi/6Fcxl0PDRB65dvbKwdGMxO6W3KT169xsQTElNXTBnBvngtSgCisBuINAAWUFrOFghK9gZzq7++oWd/J+LTcupfBXnuW+13cEWAe4NQSssghDV1SlWne01sVLbeBZ6jN1V6mA430kzBaGAc5dIC0gMjGMQAZAP6DAQbeGmn8Lp/6kYehroABA5ATmCAx8vLyRG28QxyBIMnQgcxBuM5ZkkxMR5QjYEJIrCY1J7DRdh7QyT3i9iMgZ1kNRPm/uJlkukRXGtCYsmRc38sNnwQrGQFXVyXMbmkIbO1dYoTPThRkjY/iNNLPx8nBBILi5xkExMUCcWfKRezQZ+Sioo5nCJGKQEpE2lNDRNiIk1RXXB5yZvzFk/Mr/81bYpoYECfnefx7m4U1pd6vQy572IbbHbn8gS8CJFFHiROgqMwyMO/Qn3rVHCRAmNHd+fBmqA6desJDH+bUZrJLnwLCGMztqHrIPE2lJ4FpW02CXc9SJFQBFQBBQBRUARUAQUgR0goBEWukQUAUVAEdiPEejdb+Bg8aWnzZk+FadFgyU7Ny9/5IGHHj5p4kfv11RXs8t4l8uAIcPJZ27mztwz6ad2eaBNvJBUUAMlJdSkTz96v7FLRG87rl8hWbC+aWKzWk0RUAR2DgGiGnCWE8FQv+D0/oVYXJOh2/LfOsf6hlsF1kb/aO8U7yG+SfmWZafEHO/qOhPMTjO1OelW9UZrs2+cNEq9xWifHehEPkA8jhSDfCBdFI51oiyI4CASw019xHj4O5t3JsQBhApRFW7UAudog6gHCAiIkcFCVsiv7nNMzqH5ojmRYfKO6GHyj883aX24dutSPafOLLt1kaR/qjSxyhQTq/YaJwYpAcmAk3me2BIxnP5upIQbWWGEhNhCWISgGTY7rt2yFZkhhAHEDGYLOeASG/G6t519tK8gGMpxjPMrCTs5RSYIWVFrO1abhRXpD8wtzywpCfsz5XfwnbUFdo+MmvcPyN90nd8TS80JRI4bnlu+9KuSHDAkGgNsSb+F/siHYhBNOMpJ9UVqKr7Tf3x8MhZHxka0yw6jP5Lmpl8FASEbHCEdwHOyGM8OqctYw8mF46xlngEtioAioAgoAoqAIqAIKAKKwB5BQAmLPQKzdqIIKAKKwO4h8OOfXHTZz6645oa//O6aKyZN/HiLc9wj5dJrfvt/RElcf+lPTg+HQ1sENHsJGbF4/hxSnDRa0K/g5JwZU75qqBLpjJ55+9MppHH6283X/+KFJx767+7MBOd9eVlpyeoVy0l/ss+XLj169cnMys7Znn6FK7g9d+a0PaIRss+DqhNQBHYeAZypCAQPbeDSZXIsozxqrEfWOJW5fuNdGuvuLbHyCsqd7NSo8dUd53t/6VKnTXGGVdkx1dRV5JnSL3KtTfyNTCQFURaQEuz+5/fdYjjkOySO8y57QgwH+gVipJA6VIxIARzpEAeQEbTH57rEuXbyibOYsZcJUREwnvRck9Jxo+l4ZaYQFEER2pbeh+UbX+7WZIUTsc2KOzdJNMVq0aj43EQ3hSUag4gN0kgRnQBpQnoqIj9Is8RYXN2OOHFhHbW1gz8RQbGNrlCCDICoYZyct+UYDmyIlnj92lhxfsTxXO8zsbMcx9hhxxOuiXorllelLZ1Smj1aIiyYJ2Lbjnxfsrgy3WmdElraNb22e03M2yXDHxue6Y9tqIx4SY+VLJJOxMkrYoidPyVGuizaYS7MrVrGwhA88gmJAd5uFMlWBIZGYADT1kXICvDiHhItxD3lWalPWJwrx2aITd+2BT2iCCgCioAioAgoAoqAIqAItAwCSli0DK7aqiKgCCgCzYrAtTfffldaenrGeZdcdU0yYXHaeRdeetm1v7uFzrJEH2Jj0XqcYebE0876yZ/+9eATB/QoSIlGIziwGixEB4RDdXWL5s9tkNjw+fx+8cfnIspduGzxwt2d1IAhI0bNnfX9iTQAPzCZM6PxCJV+A4cOL1q/do17b3YXQ71eEdgbEZBXRLIwr6tFwFDjOgQSjNRSw6YvCIRhYhc10Ik/ZJuRhbXmmy/KnUhZxASjVuuatU674CLTK2+e3dd6NPyz2lSrNvd0/2ttC6xi76HeL9ukWzW5AROmbXdnOVESON4hKig4zUn9RCQAmgxEcLwmdp4Y2hY419m5TlQCJAYEBamgiCKAQOBvcJzzm4SYqDbezAqTOTTH5B7RyuQe5Tep3ToYT3Dz3+k1C2vlvPABVTFT8u5XpujFUlMxVZQo6qRP5zOpARECqYAzHwIF5z3vdEgFoiaYB21tiUyIt9u0ggPb1ZOgDfCgPZzcpLLi93GS4ulUiaBIrYt5itfXBdfPK8+oXV2T2k8uJEqFSBIiKDzGsgaIHTmprNUgY20y7VNqTJbfThucH8qbvFGmZMeXywLHtsEVfM9ODBNtkXfEwJ0+p4otF+PfN1cknfkXihH5wr3ahoBp2pT3j1qJCAtXU4WUUKzV+uViOfCo2AtirFvFdP9YHjpLRUARUAQUAUVAEVAEvlMElLD4TuHXzhUBRUARaBoCNdWVlSkpKakvPvXI/clXSDanuFDmJ++99VqyQ/zE0885f6mwENsjK7iOFE0L5syaHotGk1OBbOkiVFdbe+rhI/oKb+HfsG4NO1p3ueS1KmjdtkPHzm++/OyTu9zIXnYhBAzYzW9En4IIGCJdvpjwwbt72dB1OIpAcyOAExuHJ85jd+e2K5rM+8Xd+d6c/dIPf8tCCCSTJFv6qLPNy5VRs3xJrVO8LhR3gLevdDIr/Cbql1H6U01thwyryqk1qUV1TkpAeJWOZU5uQZZTkSXnK4W0YE44atGegBg4JTFPnPCQFOhmDBbj/UjaNxz0OOchCyAocKhzjHaItuA344AEqDCWP1v0KXJFWDtoWp3cyqT1DJpA265bgRQuqjFF96805V9IRMXCLyX9E3MlxRS74l0Chf4YJ31xnvbpz00RtcWBXz+6Yqu+kn5I1AL3Mll4GwzAmogP0kxlpHjtvI2hwMlBj53lCUai1TFf+ozynI3FtYHeQmF5PR5vTFJFpVrGGmJ5vN1FN0numZwIBMxCCQiptUtNtj9kcnx1pnWabYpq48tH4mCkYzsqZhuJ2mAYkDvJGgsHym+0SVwsXS2RxxPjAw8IjChpoxqb4/5+XEiLmERaQPCQOgwtK1Jy1S+sJ+47kTusX8Vzf184On9FQBFQBBQBRUARUARaGAElLFoYYG1eEVAEFIHmQOCWX195Ua3oR0yfMol83lvK0w/f+8/Z06dMnpekj0BUxIgDDzn8teef/N/2+k5NS0vv3rNPv+cff+je7dUr2VhEDvjdLlv0K7YTjbDbnezhBpgTxJDwOjgKtylduvfqs1kj5JsGU27t4eFqd4pAsyAg0RS0A1mAI9M1HMo4jyEpIChcsiJeV65xCQW7GaMtGAOOavQjCutPTkY5bkG1eaEs6lTftzoeAYLTlbROq+Wcz28iwaAV8rXzrM+sdDLSv4qNShX9iizRssgtclrXZJiq5W2soqCIcRMdATmM0585kiIK8gLHPZENkAJETnQWmySGs5xjpJFCTPoHCUxw9jIOiYqw0ozHn2fSB2WbvCMlXuF4n+hWbKtTUfTKMrPq39NN1ZyoiVVUSFIlIj3Q1eCTaIouYkROMC7ICo5BpqCdgdg3pU5Iil0hjLinzJn5SmCERSTLaElf1U6+TxI2YVSKN9Yu4HFMSTggqaB81ctCeZ9VeHMLhbzo5LM8Q33BlBS50AhxUenx+hiDLxoW5ihdMm2lpEt+rDwBZK1JdTaYVukeU5smUHt9PWKRsIlFQsaOybTDdfI9LNEXcvnmtUfhXiIKTSTLhAQO4H1IYu6Me77YGiFeuAcxJS5c6Lb5JFJmsRg6IRAWZ9arUSi/ecZ41rYrft5oD3pCEVAEFAFFQBFQBBQBRUAR2AkElLDYCbC0qiKgCCgCzYEARIFkYaqV1BdNTq3w5YQPG9yhT6qmGVMmf5E8rs7devQKBILB7aUpon7fAUOGyW5XrxAejTrTuwmhsamsZKP8PzuGt1vQu2A8diwu+rpNGeTqZWxH4HtHfezp84hqg1FDESjMt0//gUPefOm5RiNG+g4cTJoaM1sJiz1967S/FkIgQVa4JIUrRo0T093ZT8+k7UlORcffm1iczOA9IY/WTu/Slp3g9WdFm2hMsNsf4mBLiecwckxlh6DJemq9idTE4ucZL9ZKtCvmiLC2Z4PTpl3YDnjyrZK8LKsy0NZanxIx/iKJwvCWOPmbgp7wNDl3HOMWYwAQFTjywQCSAmcv/UMY9Bf7WmyuGHoMpFM6LHEOokJIBCtg/HmdTcaQmEnrnWXyjk4z6f0Cxpf17XvTrouZjW/ONSXv+03RS2UmWiE72236YuwQLpAURHewK55+KIVi7IBnLJyDrKgVosJ2PjQejO+Jutv9EAc/c4M8gYAJCeHQW7TAfUI6yHfvcV5foLO8GFvZkdCxIV9qatRnTxFVDXtJXU4s5M/3ek3kPG8wrafH57e8Xr9wDNKtZWXKbxmE1wQzBAqPd7PghCfFlEWzTK5VYVKDfhNwRLojkBZPDSX/mMQJi7rKMuF2IiYaqhW+xo264A473AuEoiEkGCtrAbwhKrhf4IF20Htii9G5UNJi21ufJL7N2trmIZNjPDusc/DluYYMiheeSbm+KctK6ygCioAioAgoAoqAIqAIKAJNRkAJiyZDpRUVAUVAEWgeBMZ9MHnWB2+9+uJ//nrLjbQ49pgTTznrgkuvEqmIvI/fefPVR+658/b6PXHuvJ9fde2Bhx5xFDv2P//4/fH3/+Mvt0Qi4bjjADIALQvhCmJoTnDs5DPOu+Dwo44/CedgTU111ZMP/OcuogHctgcMHT6K740RGzjrn3rz48lff/Hpx9ddcm5yKo6thte7/6Ahv/7D7f8YedCYsaSg+tefb/5NQ1EbpE9at3rViuSIjcOOOu6HRxx30qmks2J8lRXlpPBo9hKQXb4/u/zq35xw6pnntW7bvsOalcuXgSFkw/IlC3FubVXA++qb/vT3Y0/+8dk+v8//8L/vuK3+fenVd8Ag2t0eMdR34JBhEFPzZ0+f6vcHAj+9/FfXHzz2qOPWrChcds/f/3hT8YZ17GhtlpLYwb5LjuBmGYA28r1HIImscMkJfM6uoDS770lR5DqKeZZJNYPjG0cnUUikKKIQcbG7uhb0DUmA2DTO6hOTb4DkITKSDiqwLmwGlkedOYlx8Xcv70w0JroJKVESNsGIpIIq9nhsfxureECOVS6RFdXrNzk57bwWQtZOpm08tR5jQ1IQ4YawNYQBnzy/eM6ZKzv+0XXomRgT5AK/IQnov4uxfP1Mavd00+HSQ0RUO9+kDygQrQrm8G0JrQmbBZevMBVfLzGRkvbioed6PMJxwWsxoiu4xhXsdiMpiITDmUwd0lNBMvuEqIhftyOyIkFSQFQwT8iRPhIY0dsXtDbJ5zES2DDK43WyfCTkYvQAACAASURBVKn+TsaWarbTxh9IybA9QbMmag4NRxx/rZXSzopGekskhfAaPuMLBIVoCAgxQRYo+V9hPeJwyfc4iSG5ooT4sKoDbcwqISrSfdUmW87hGY96N8MCacGNZu3xPRIKmVB1WTzqIs75b4644N5DTjBXOikUw/EO/q3EiI5hzYLZrkSaxMfyPS+sV8gvV7Mlebrg+2wCP9abpoX6ni8GnZ4ioAgoAoqAIqAIKALfNQJKWHzXd0D7VwQUgf0KARzhHTt3Ja95vPzqxlv/euFV191YurG4CL2DC6685obH7//3HcnaE6Qd+s/jL76FBsTcmdOmRKOxKNewwx9ygHb6DBg8ND0jMwsyoFXrNm25PijMRscu3XoQIUA6KXQoksGGQCgvKy1ZvWI5KUS2KTgUizesX0cbjd0knO//+t9zr5UWF2945tH77x5zxDEnXH3TbX8f/+q4Z4R7IC3KlsI8vvp8wkccYOx/vOu+R088/ezzE45La8iIAw6+9KwfSm6U5i25+a0KHnzujQ+79uzd980Xn31i4dzZM4447oc/AsOF8+bMrE9YQGg88uL4Ca1at2335kvPPIFo9hXX//5Pb7/6/NMQLu7ompLiqk//QUOXLV4wj2sefOHNj4aNOujQEgF1+OiDx3Tr1aff+ScdcUDzzjburFOHXDODqs1tRoBUTjyv8hWnNiQEqYhwBEMaQFjwyTlIC8hR1iL1MMgKfM84ljnfHKQFY4F8OFkMomBL4UEQse0Zsyqd5aJdgSMbUgPhZq7hdDvHWJkRx1cSsXzR9XabnGyrwhESI1RgbcyQtFBtC0xltuhZrAma0GIR4W4rs2f8z4vh0KdP5uoSMjhyIQ1IH4Wj/GOx58REhNs6TAS0M0ywQ2fT7f8yTNaogEnplG48qd++kyu+qZVoinJT+l6xpH/aaJwoURLgBCkCEURfYEfhHAQQv6cl5uRGV0BUQKAwRjAn4qLBIiSFq4QOO0AfECPgiZZHf7lbJ/oC1qDUbKt9rbRuifxEQRdH9CfsaN0mT1q4VAgEIRGqTabfFn1wn0RTUHyp6fEbDUHh8fCfGoK0RFRQXKJKzsWruAPbZOXIhFLFWy6hGklyJFznT8vkMmEoYgFfME2qSJooIULCtdWSKiruO0fMO9sVu5ADpOBCkBscwI00UQxgpsy5VqIsGtRsagyn/eQ4UVGQ96ynC+vNmWcLQfs3xEgdtVXRKIv9ZIXoNBUBRUARUAQUAUVAEdiDCChhsQfB1q4UAUVAERh+wCGkqzBTJGrh/J//4jqc5m+//PxTt990zRWhUKguQ0iHZLKibfuOnf779KvvcuziHx9/+LSvvkBk1Nz92Lg3Tzv3gp//52+3/o50RS89/eiDGOdwzhOp8NOTj0SUtNGCwx0CZHt1iOBwHe7163Xv1bf/Px565mUIgCvP+9GxVdLpxA/eefPhcW9/cu7FV1z9wD//eqt7TZfuPXtn5+blu1oOt9xx7yPHS7TDv2//ww3PPfbgPX+555FnfnD8yaeRgqqhiIddXTnoefz3qVfeadexc5dLzjhh7KypX5Nf3uS1atX6gEPHHuXi6bZP/X88/MwrecL6XHT6sWMWzJk5nUiKcR9MmgVxUZ+wqJXQlaUJQqKhMSK4PfGjd9/63Z//+V+uB6dJEz9+/54nXnr70COPOWHwiNEHuWPa1TnWvw5/cjNqBDTXsJqtHdkx7pfd4vF0Q/LddXqyg1xLCyIg68oV1HY1HEgfw+51dmXj6MaB7upXQFaSpofoC9Ii4dRnxztOY0gMN5Iqvnl+F4ft3nvWAn1tVcLS6qaoKVghlEpFNC5MTQQEO+wZK/2vE8c4c2kj6aFSYsabUWy3WlNl0ld9FjukdYmTt2aEd5pvWmzomvaedUuP9n10nGheDJH6ESEuSKPHuxMCBJJioVhXMRzhEAWbtS0snwg0+NtK6qc+JqVzhml1QobJPVxEtVtbJloZ2kJYVM8JmXkXbDJ1hZtMrEawc8AJgmWdmKvT4abhKZRjGNErYOpiSWQdBBIGptQnWKHB6IpERAXaFBBOYALhBJHTl7l4/Z6b03Idk9veEb0Jb7Fkg8rzB+3aYIYTDdWkSu4ny2yqCxuPL8V4U9JMMJAq32WJyPuHTyIoHMnJxaeQE+AS/28OiZKolOiLBnMISbSLTLbB5UA0jkeY7ogM0PIEReJb2vUIQRKLyu2PZ4faopFCN0TAQByRMgsjQuAksdfFJsncIZErND0UUG0pPJesl7heSQOFZ8zVYNmd57aR5vWwIqAIKAKKgCKgCCgCioAi8C0CSljoalAEFAFFYA8icMCYsUeFRcCiSrz7pBx66an/PXD7Tdde4Q4hOSqByIjbxZGPHsUlQlYskXAAt943kz6bQDqlDp26dFu5fOlWOx77Dho6/P03Xxm3vWllSt6oTl2793z39RfZAdxgIfUUotxEJdSvwNggGSA0rr34nB9BVlAHAgCi4sO3X3sp+ZpBw0fFyZNZIhAO0XLSGef+jHkzf47PnjZlMoRFu46dujQnYfHzq39zs6RlihMFycTAgWOOPHr+7BlT66dkImXTwKEjRt9wxc/OhKxgbODAZ0yYoeQ59R88bOT8OTOmNabZAUFDVEymgH2kzI20WpAVtDF18uefQli0l3CbZiYsXCfurjqB9+DT0PSuhJhwU/+w03eT/MbJioOV6CB2kFfJsbjQsxIXTcd1J2uCOY5/SAic4ezIJ1oMoWOO8zclRMX6hLkEB85pHKFcQ+QBaxOnOsd2tbhOfAiTn4j9NLkh0kEJSTFDKtUUR0y1+M0hTZaJkRqojxgRH0QpjBZ6LzXkBBcErXBdqZOXfn/40k6SIsq0skrmppq6vE1Otj/Nqg2EHX+VT1JEiUMdogbCgnniGGcdsj6ZF2QF8xasPD1MsN0wkzu2t2l9Rqrx5aabnIOl34T2uD/fb8IbombtwxtN0ctRU7MoZJwIURqQPjiHISLog13v9IHINmN2DTy5Jy5BAXEC0cH1buot6qBhYXguEhEVYMe9guAgEiEkZEBECCnuJzvrj5IsTSarbcC06RkzWW0ijgQ05Ao54E3Prc0I1dSZQGrUeCXlky0cQc0my0TqomI1JiUzJx5JIe9EIRNEo+Lb5EJb/nvD8njYyd9okfvR0DlAY64Cn/AWHr9je8IidZERJ0Sikh4qSYx78/WWaIU4DumzWHPgib4IGwaIfHlUDPICvLVsRoD1y7qBeISMi6eMTCo3yXfWPn9vQKSxtr5X/87oQlAEFAFFQBFQBBQBReD/2TsPALuKev/PObdvr8lukk02jUAoARJ6aKIiRVRERQH1PbA9K4g+u/LsvWAXnwWRZ1f+iqIC0nsgQEgIaZu2yWb77t29/fy/n7s78WbZFCCElJn3xnvvOXOmfGfmZPl+5/f7OQT2HgScYLH3zIXriUPAIXAAIDD/+IWnPvLgfXd/8KovfZNAzF/4xAfevb1hQ+zjOuhzH7niv0rFCsorJEXRzQcupkqfJ+A2MSwQAHYE59x5Ry/g/o4sLOYeftR8XDcpKPfT6nr1G/7jrbih+tInP/heXBzZtojX8IOvf/6qsW0TYwMrEVxfffcXf7wJEcSKFZQlvgOfVvjYHUuB/l36ris/8rvrfvLDe++49R+2TvChP9f+6NtfK20HLP/zne//8F23/uOvxBix9+YoDgXfn1q65DF7DXdbsxRx+5c/+f63ttfXmbJA4d4pLznr5b+59prv/evvf4EgKyYEq909XtUH02dPsO8OCPd4HSJWIZI5GQ2pXDw3rXyEMmQqrskgg3E1BHkLiQkB/agywYW3BoLd4x3fDxscjVfByCzBDRnfqswnpDMCEXufU9eHKEMOQ6ZDLCNiHKa8Rpk1SbwHSE4sEWw8AYjyXQoCTSfGCbjNOwOhhDWzNVGhXEH9XNYVS+/sDfrlEupgXbOuq+gX/YGs50R5lwjyGuUn0ybqDwWJU4YKidkTvI726f5q7kVm+ysnzfJXVoS9fJ/iWCAaI8DgYmjD6FhZl7OVeSdzcn+L3D/NNqHKOQqsHTONr2oyDedMNnkF0i7I7sOPS/PIFczgo/1m1cfXmp7bZSaQhHFHUEH4pV7WN66ZcGtEneDHONkPYMz7g/5bYcISx+wJa+UCJlvxHRUr2D/8mzEiPnneLHkinCSVYb4XFBbISVfxkZqmgmlszSsGBXEjCl44WggX8iFTJqQUWiLZv9kk00NmQrzSM5HooOnrCBRPYsQjE56eRud1VJmhG6MpCB7VCGR1UnLtGX7F0CJaXplVnAyFy0iHZK3hZ+UaKjuM9kD/vWKgbgUIx5ojrHWMqIVoYRPzh8VFUpggIOMiyhHvI+AhIvLvHO9S1vpY11CsQfYcApB73z7DteuKOwQcAg4Bh4BDwCHgEHAI7DoCTrDYdaxcSYeAQ8Ah8JwQKCsvr5h50CGHyutTdX3jhImvfckJR+DOabxKsWAgSPTqp55c+rtf/uSHY8uUlZVD4BrcSJXesy6nFj9039076izWAdxfsvjhB7dXDndFiAxPPPrIQ6VlEBcufff7P7JuzaoVv/75Nd/dFVAOP+rY43Ed9c4PfvwzA/29vV/8xAfeU/rc5GkjcT3GWovsSt3bK/P2Kz78KSxWvvHZkTgfNh138uk6QRwKPXz/PQTQ3ZpeffF/vq1cPrm++5XPfMJeRJh441vf/X4sRzauX7vGXj9o7mHzEHOeWLxou/gRo4LyA319vd/6/Kc+XNoWrr/4re5BPu7OtE9YWEiYgDTldDoWE4gTuL+BoIWYJUGKQ4YzHnzQ88nJX8hmBA1On0Pq8okFzFTV2SfRYqt4tjtBPUDrGo2QXMSc+YKUZy4g/Zk3vvN3JGuZawgWkO73K+Mm6kRlRDqsYIj9AvnOJ9YCRSJ9JO52kSV/pon1AAkNgbqVjMayAldQYvI3y0jALEma8mxQFEgg9m0QcNqiv1wnPoTsAUKNw0GiVoJEfSEIxXtNbfmywsHNG4NJ618W/rtsCIKEYkoPxL0URC0nzxE8EGAQayxTLqEinpZIcYapOGyScsRMuKDWxKYQ10Mrtyxsum7qE5s/bNq++rAZXpmVCyj5TsqDH+6d6COEMesckRR8ESb4BC/Wu7WqGFEW/i1IbIPh2ADbo+6fmCvI+9OUi3GLRP5PUEyIE0KR2BESJnRhsM3389MmH5Y2tVOGTC4dMrFyAViXkhVDOBNJeFm5hBrwvHz/hiWJZFntcEvtlFQ4kghMT3u55lNQyvZCogViyohgEQS3qSH293R9HjHqrm5EWXiWSVYcyVAs9mBgclUKAD7Ti0cTnpcoz2VyRbFia9UKxKH2Wb/4ycvoO/9eHqnMv3/0CTE+I3wKEi12WTx7lt3eFx4DA6ykmJvx3qWle471+mz27r6Ag+ujQ8Ah4BBwCDgEHAIOAYfAC4yAEyxe4AlwzTsEHAIHDgKzFAsBdo64FL/62Q+/s2blU5w2Hje9+OxXvJrg3Fd94F2XjedyqLF5EqccDUGzSyvAIgMrhrZVK5bvCFniV+AOqbNjE6TbuAnBYuljixfhwqq0wIte9vJXTWyePOVrn/7oldsTXErLQ/pLpzkCi5KXnnv+az/w9je+RgYiRQsDmw5SrAf609vdBXG3NZ31yte8Yd6C404s5Av5TllyMN7B/v6+YUURR/iZPHX6jCN1f8nihx747lc+u1VowNXSKS8+6+U/vvrLn03KnKG0TlwxEcH1kQfvvav0+nmvuejNWKY88eiIiIMrqC9//9rf1DdObHr/Wy46v7SsDbhty44HIPE4uP6La77z9bHjramrhzg0G9augeDdXelZE4C7qwNj65GIwDghBiG4sTjhE3EK0YH+WmITUhHyl9+cnLfuhyBoOc1v/evbIMIQ6NQBsYvrLsjcjWoPAhqy/A5lTgjjjx0hY5v19nyNd3+od9SygrmBcGYuEIQg+JlHyEzm6nBlBAnKMUdyOmTWjc4fZZlrPomHwBpnPqiL8ggH1mqjGIvkWSbIU06AF+MCwbQiWGT15amh4IENaRNePRzE5A6KucdKAWGAfrWOfuc3/cCqYc5oPIsB2RRsUeDtqiWFQ+pa/bbH1wYtHalcvHk4FM/NDS3dpMDcixXuGUHNuoHS+BVZOlReZ2oWtpiJF04JymZXeWUHNZlIPWLDSJJ9mVn9qb+YXH+TxIqbTSENs05/qIt+IKCALX+bI1rYGBXgyB4AZ7Cjv0VXT8pbCeNRl0/FpuYv3NoqX5hHBBb2Iu+ks/XP0OOyTDhZn2dHFH8iHEsoeLVcPcVD0xq0e2IVIROK5OT6qZAury14lY25cFDIypohCEsDiCeqcvVltbmBwS0mGY4F4fK6XC4UCVYPdEYnZdORBsXh7pbI0yGRQNYb5m4JBQ36PiIIBEFOGA+rbY2TXBSu2vQbPFu36fnTf1AH41knwbg/FC5Ph2oKvqeO+eGheX2bymK5dMSkB/uxDBE4+j9pKHIbJQOSAvUXLflG0zz16cyioDJCzm/z79xO+rG/3ub9i7DIgQj+PtlGaNdv9hpYfUl57f4KghuXQ8Ah4BBwCDgEHAIOAYfAC4+AEyxe+DlwPXAIOAQOEAQI3sxQIfl/+t1vfHFHwz7n/AsvgWi/8Q+/vm68ctSF+6SOTRtxH7I1HXnM8Sc9/MC2lgPjPY+7px2R7TxzhOJO/PWPv31ajIvzXnvRmzOZdPr//fbpsS3Ga+uQw+cdjTUC9RFs/OYb//S70nJySeLPPOjgQx+8585/lV4nUPfnrv7xuOO35bAAefzhh+6/787bbi599nVvfus7iTnxq59tawGCYHTSaS9+GYJOqdhD7Aza+8LHrnwX9Rx70qkv+ujnv/H9ic2TprzvPy98xVPL/u0OivvgB/5YmWxvHltnzp6Di6wbfn3dT8eWoa2uzo7NiEu7Y/lzUl312BPxe+SkMHEkRJKmRwNfQ/5iHYGwQCDis5URFThdbklvPiFpLREO2Qqhy2+ECIhb+3eJdWtDGa5Z4cKWhTSjDKf6ESWwzoDYJbAumBIzhVPklL9PfYQIXqb+LtJ3f+wJ9N0xB/tZHeBFZj7BlU9Ic9w8QVpiFYN7ITuXzB2kOOuAeYdsxzKLZ7YoQ7IjMHCPWAs8y5w+W8Gi1PpjBHrcEWkXSLTI3dJjtiR8QxTmYS0SiHr6xvv3tNGx0D+smxiX7XOPRIunFIGhXREYpuSDeP3GwqSKP2bPy1SaQe//5c5e/fboNcMnhO7tavY3ZSRa5OQxaqU491iucv5Rfv3L5gXVCyd48SnVXqSmplSsKAw83Jlb9p4/+IOPLQ8Xkowbcpx+8cmeQGhjf7DWb1fmvU68AAQixAvWNGWx5igG0h4Z8b+TrARKf/LdvhMQ/4jhMV+5Ra/Ai/xw1EQS5SOukxS4WlYWEicUOLsibBI1nWZgS30QCieT1U1DffHKfLXnB1F5YtqaCH+dqCpkIzGzUoJFLt7nyfVSPl9e17ulq83vTvaWI74gpmt/e69QT9inIzUgTBSCtESEHgXMhhSXd6fIkAJe4KZpZ6looOGH8oeEY/lGubDaVFFfyHuKVB6vyN5UVh05pWtdrCYUrjepgb5ibAseGHk9Pi1FdPXDKkD8jj8KPxv/YxtcZXmxsz7tT/etWyjECPsOHvvfiiMWKyPzuUf+rdmfAHZjcQg4BBwCDgGHgEPAIeAQ2DUEnGCxazi5Ug4Bh4BD4DkjQMwDKiGWwaaN6zmNPG7C5dLxCs59601//uNY6wYeiMbi8aOPPeFkYmFgKWArIcgzgbR/8/NrvrejzhKrAYL+T7/+xU+2Vw4LBSwLxlohlMus4diFp55x3x3/+udYa4jt1XW4TCCK98QcfeWqD18+thxxN7DCWP7EY4tL7yEqnHrY1DoCe0+RJUWd3GjpKK2flxIxPJRM9nR1bpFesw7RYmydZ5736gvvuPmmv5TG16AMAbgZ152KU1H6jHWlRb0//t3fbsdS5amljz960TmnHbNy+VJiJmyTDpYIQ1DuUvzHlmmdddDBq55a9sTYPlDukMOPnL/8ice3Ge9zXGCWPMLHznOsavzHCdyrxN8NkM6Qz/W6dp4+IashUrkOEd2qjAWQnRdECchYiFaI4+JheGX6THl+U4bvw6LCIiI4+Q7ZTbYn0CkD0QwBixBigzxzip9TwbgHog8Q0dYigACxr1CGFD5S/WUtIlpAECclXOxul1yqdt9MYywrWETMH/OAAAW2WAO8avQauHEN6wvmEVwh/8EZcp3YAIhQiEmc6mcOmX+IeMpAwlP/s3EpQ3u0S33bnIrPaCXJBVRnddgctnxI8aBzxVPguLJivfCMJVpHyfRifBTWFfUUrT8kVrCu1ormbuwPKlsGgooaaR/pJn/TzD/nzupMmVj2pd7Ng43h5IAfaz7Uqzi83m+5fKFXefjJWpLxXG4g7QdejEpkTJDPbfrtY6F1X1+dHlie9wLv0JgXmSrXU40hPFGN4IIFCt8ZD5/0BSshMGKdsj+wEsNSBOzGdSOo66XJihXMH20gMr1eQzxlRKBQDPBoTFYIiks9GirGC8X0iq4xmWSkP5+LdiVqsvGK+iFiVuRUZFjogB0YkoZ9P+hUcO5fKVTErER1IZLoMx1DveGWRHW6Mz0UO1MupBBcGiRMpEaf5/WNkKE4F355PpvZIqVittzzac96OwzEbQemV5uMKQopX/Ye8iQ2HI7mw2XVmbCiVmwur/cflmwSjZX3H9ezMVzb1RYvBuQ2EiuCzLDxIxqrrC5GXEYVU0xrfo5q/LYf1ivH825Un/pdPIvi+rIWboiLRWvOksT6ZK2yFmyQ+DFF3E+HgEPAIeAQcAg4BBwCDgGHwHNDwAkWzw0/97RDwCHgENhlBGYdPLdoYXHDb6776Y4emnPo4UciStx/1+23jFduwQkLT+P+HTf/7c+l97Fg4PdYkWFsHQSj5tqyxx9ZtL1+4IapWNcD27pNOvq4E08OhyOR++64dYS+3oV0mAJcU+wvv/u/a8daKnD9oLmHz+PzyXEIfGJQcK/43Bgrh+01jfUJLqu+8+VPf2xsmbNe9do3cG2xxJ7Se0cuOJ4guuaqr33vJwpVseqTV7zjP/78+/+7djx3XNFoLDZD7p52FHAb0al5csu0sdYktIGoRP9u2IFgtAuwji1izz9DeO72hFWCKsVNCFYUJyjz90OrMoQvbmqOVYb4hRy1AgWn6nnGChd8jhCpliWFAlUc32J9IiN1B6JMrGJRuKAkhGuv7oh9HK1nRI+xlheQ5GuUqQMCHYKNfmGBgSiI2yhOl0OwWTdE7EMI0gc1Lj5XYXlRrPXAThYfiEiEBkhySGccDDGvuPLCkgWXaexL1oKNr4CAAYYIEggV1MGJfuaEOtYr45YJYamUnKbNXRItjmophn0h+DbPUAfi1Wu5RgUSKowEisX6WDeYNw1PDAZdKYW21i2I/hZlLBuw9qBPBMrm04osrA/EAcq2Ul5BD5qVl+EqSs6F+juD+ujd+RPSGwqT1x6UyFRWN81oiZa3TvZrTjnZk3Bh/ARRpwuFfFo+67oGslt+8MTifr+9efBGf27waKi90BIeDMq9Jn8zFhvry7yhWokWNmA448HiApECvPjN/mFdMwYy19jfOzvVDj7sG+pmfrB24t+Gk/2QLzkmbAq5rIj7qESLRNHSIiQyX8JBkMuEvMxwoaKshvgV0Uw+Gxn0TKZfOCRF++POjbbJCck6E6PhAMGyUxYYqZpJydZkX2W2t71qmh8Kiu7wRpKXLuTS/XJBFZFtU0rCAH3K6+eUoknMiADDte3GtSgW84J+P1QwkVjudu3k8nA0V1/f0pMuqxkOJXvKyoIgMl3FHq6bmpo9YVZ6sO3BSHXn2lDVcL8MOvK8cnwJNbGi1QXj35qCoFbBub/uhSJ5CTl/0PUDPZg084GrSIS+e5SnKRO3xSb2HAcPWI/Pjzpe0pj76hBwCDgEHAIOAYeAQ8AhcGAi4ASLA3Pe3agdAg6BFwABiHl5Eeq9+18337Sj5jmZz31O8I9X7lUXvvFSTvbf/Ncbfl96/3AJFlgjENx6R/XPmXt4UbDYUbkj5h93AsT9WOsAG7vhwXvv+NeuQijB4liI/x9+84ufHu+Z2YpvMTLe7Qsou9oW5Yi9wedD99yJb/KtiUDbZ5x1XjEWBbEqSu8hIGAx8pkPvfdtWLbgyml7bc6cc/ChuLh6csmj28V54qTJLbi6ktenp8UIOfmMM4uuTwThLos+Oxr/qDsoiCOdOn5WAYx3CO+oOyUbXBniGvIX4hqhCZIVAQCCGwLLuqqBYK0USzji9icQgR2MxjDwJE6EolkTkpYRqfNMotU3XrkIy5xnBpdIGJHVUBgn+rUFk2rTuHQ9Kyra46R3ZkAH0/uL8olXJHT5hiBhXUZBPPMdSwvuI4BYSw5LuiNqQFyfpQyxu1ljPEOfkHOPMQ4JGAeiP3vIcYQGsLMBtYlbgTUNFjKsZcSp4v5SojyiBuwv2FIWwh1hA5ITQQOXP7iGwnUa82JjlIDv09wajda7Kx+oF8wZ82eZ7nYtlkcUICFTGTJVEjAUR6EonhDLhPXaqsxznPJHSGOtEOsH0YJx88m7txhfRiknsaJI3oqwzw4FZSLvQ7019bUTWuZ+7qBoItoQjlQcH/gVCuAst0RivCHW+7Km56crupfU9Hf3VOY3lHeYqemsP5S4LbewJWuiq08J39kzw1+VCQe5e6NeJibRAix4l2AFgWhyqzJiA3sIAQicsAbaiRj5C8WuuJi1ztwxXixjWOuIsW+SdYOJllWNuoLKY+VQFC/C0XhOQbL1nGQHSQZDvQlf1hFhXemRBUNeIkE0WpbtjJZlmE/mlzllz1sRpUPDps05sbJ0c0V9skVAmWw6LIsGTCK8mIJ61xPhW+8qPRMIUw+TBgQK1g/C/LjuNT5LaQAAIABJREFUoPQEvXokVp6OxcqySdW3OZLILImVZw6VS6jKSDQbCcezTbL2iCSq0muaZvcfppmQ5Uc+GqvwOnP/iM6LJsp9xbYw6eSw3DFmigw7WBStL0aTZKYJBZO9OBIpu+uks97dftdfr35ehN+tDe79X1j37APWH8IgVhasKRJ7jr2HG0Znobb3z6XroUPAIeAQcAg4BBwCDoF9EgEnWOyT0+Y67RBwCOxrCOBiqUq+mIhJMZ4Lo9LxNE5o4lS4GY/srm+YMPG0M895xV1yadS+fl1b6XMErl755NIlxJfYET5WONmRW6p5Iv0Xj7GuoM6p02dx6lLBots4Kb3TVNfQOIGx3/2vf/5tfdtqYgo8Lc0++LAj5IlpcO3qlbjvec6J4ObE/9goxaW0MsQKhAju4aqp9J68ZNUj0IwVgcbrzEEKysH1FcuegNweN6m6IumpGOHbBBHn2ssveMObiF2xM0uYXQGiRKyAYNulk+q7Uu+YMoXRWBU25gCENO7NGCPt8rcELnYggfExM1QUJyQzGD+mbxPiJtYSMrGmhElMD5tycZ2+V2WST+YVqLhgvKgvQUJHpxs8M+lS3+T6dKBdx7+9aGBS6wckbsgdjZ826c0pk3wsaVIKMTAshz/ppMIqF10/dakt1jxudFiXEKqQzxDTXId8o2+QqnyHTIeAg8xlD/EbIvYK5WXKN0vAwCKgU+PeJqj9s8Bun3hE68iKOogVEJPgZAl8SHxcK4EXlivgaONbQPpzDdGRU/WIFhDwENGIFOAKhsxLaSwS5uUZuy+TdQX9hDi/QPkzW8HVytf/N8d886K+jLl9Y9psyAQmIfECawXEKYQA4m4w1zbuBtw1Y7WxVayYAZMNEWstgtjDlRNj3pZ3zKwub0kE8ysq6l+aD+lkvq6LkvdT2Ux7qpBLLevp77lv9Z2LHu4JZlSZGdPm+LlcWzB1cEl+bn/MyyiAxLrI8sIsP2bS1VE/o0WewQoIQYj3Kv0ENyvmgC347YpVhRUrEF4QOxgrghzr/FwsGXB7JHHCROKyqJA7qCJpXyj0S1DQeD0Ex2Ii3kNmKFLWs6FmWi4dXl1eO7RZ46wORXMdoXAxcDW40Df6mpb1Qn8+Gwqlk9H2zFB0kr5nAjm/0r2i+yhZLwyqnYzar1Nb7MPi5dGMoIh1VlF4sgnhpyhWeMGgPtfo55AEk1hNU39vJJFdPtwf92VpEZeAEU4nY7KcyG6QyBLVc5OjidxGvQ86K+qDGdOPydySTuZb1y0um9W/Wb6tcmGTHZYDKUlRip8xammy1UXUqcLk1Xr2xxJ+kgewayjmBlBYm1hWvEzZihV2ir6vL1gw/lYZF3A7s/opnV733SHgEHAIOAQcAg4Bh4BDwCGwUwScYLFTiFwBh4BDwCHw3BFQ7ISjqOWuW/++TeyE8WqWtyeIQkM8hbH3L3vvBz+GS6brrvnON8bemzH74LmPPfzgfTvr7YyDDp67avm2hH3pMwonUSbxY97vr//ZNWPrqq1vaEQQsa6adtbWYUfOh4wyWC1sryxCywq5e9pRPIidtVN6H1dMHe0bIJy3Jlw0ve3yD31y04Z1azeua1sz1oKiSooFQbB3pR3w4/nVK5ZDbo+biMnBjdSYOSQoOmvh2h9e/dXx3E3tSvu2TEn4Ei5B/j4vpJFI+0AEPu59OKmt0+RFEovT1RDSkKMQwA2iIGOirSRSiDasPFROWw4PTMWhMROVu35fxULluq8YyAWdfQ/V5Ez1SSmT7eOYt+wvDk6ZUDxj4tPKJVj0GU/fQ5UiRL1O4xWqTLa7zuT646bh7LAZXpWS5UVE9XSaDd9rMzkVK2Q5Ok0Gd8hXiFFIZ8hfG1vDximABKb/3IeARXiB2Ca+BqIHLk84eb9F416q8T9A/A597pdpVKxAgAALYj1AniMogCFEMoQ511pH8fydPjlhzzoAOwhsGxMCEhvRAnGL9xd/Z/Is1mIISfZU/rPFkv5g4QNhvpVkZ+EPqZedWbP+b13B3YsGgozECvrP3FvRCiKW9co4SdalDdcZIwS7HS9iF+shpAAJwdQyP3bZ9OhJpzeGT6gIe9GysDciKqcL6yJesHZRR993rlmxOehKFybX5MP+UBBv6g6qvWqvzySDMqyDanNBuGaDmRQbKFRGZFWxudlrPzhjhitCXh4ri0nKYEf7rEXeRbinsi6YtuI1TnBt7rEH6TOurhBAECqOVtYcIanIYCmiLVNQV2RZgVihlMxn08t1z9f/y92TRMTRhGiRTYVNb3t1pmNlww+rm/svlBARkfVETu6eshISHpeQ0CPBIDPUl5jWt6myabCzIiehI5rsLkukBuXBTdYVJNVfQfv/rhsLCzOk9xV71QZPB/+theSdSSJEzkgs6ZJ1RRCvTLfX4f6peniB2jtm0/LGLZF4Ll1eN9Qa9vODw4Px+nw+lKht7ivo2WnqX1z6TO2EWfm0BJN1dVNznW0PxY5PJxNmsDtqFBhcYkVxzre2qT7GFMPi0EI6jwtD1uuBbD3AnsYyincmAdNbt07gyBf2HnuQvYh7uF2KQTKmDvfTIeAQcAg4BBwCDgGHgEPAIbBdBJxg4RaHQ8Ah4BDYAwgQl4JmHrj7Dtx97DB1bdlSJM6xTsCFlC08W8T+ay+59B3333XbLffeces/xlZCIG0CetvrBMiePLV1+thg1rgrwkJje52Ye8TRC3B59OhD9+MiZ5vEwVcEE+7nc7mtR1O5dthR848dG/PCChb33n7L0/pLxepiNf2+5/abCdK7W1J5RUXlWCuWi9/6risW3XfX7Wec9YpX//76n/6IhnARZUWDoeTggHSiosiwswR+sk5ZO15AdPvsoCaO71a4sNff9cFPfBa3Xf/3kx98e2ft7Oj+qFhh41Y8l6q2+6xIek7Ss24hnDk9T4bctQQwhC7kqHy/iIj2xTJWHOaZ6ERRhSdFTOV8HWfW8g3kNN6XFUUooec8sZCtZRInJFwMd5twdbuJTw3ps1ZeYlYYP54VmwrJTIIsE/OZH5SFhshbrb7CUNQkplWZwN8kAaTMTH5bh9n4w4hZ98MnzVDHYtGfM9SbySrapD7hpgh3UUl83usTcpIxQa5DDDMuXJ4gYLQqI0AhWFAW8piyC4QDUsWP9dmHpclo3/aLj1ELHbBg7UPkM2bGz7yCEzjwPgID/mZ8dLQsc2NjVUCO85vnOTHPO6u4/pUeUMZ1DNZT3QSEt8G9n6X7MuqHiMfCZ2tiUcqiwrQNB+sHcqZKMSw6CkGRkIZQRQDgORsgnOJWOOEdxpzSd8ZsY3JkffH8TXG/8sT60IKLp0Zb5lb6tbVRrwaXUyL08yGt9N9tyN21Oll45Mb2RPum4Slz5eIpX+MlpkRMtqvO695U4Q3WygXUMokRc36euWhKyJtQPt1vy9R73RUDpjIxEFSm6kx3ssIkH1FMC/qFJQtYWcFnG8up7YgVKAOMj/6/XPvkLMF8gpQCCQtFl0x6aUdlVZGQS6jKonjB+CVabFT8igrdFRYep+kRmmxMjSK2cq80ecMTTXO61tWujiayNZMPbX88Es+uloVDYziSfyhanhluXzbxP2RdMWGot6xSMTBk9SAxIL/90AbqjshwD7IbzK1AhDBjxYOs2ihInAhVNAymJFrU1E3pbdK1Jj1bxxuorqX38NRAbJrcV1XIHVRNaiiGuME67ZDFR0XIz2N5NRySXVc+MLIMCfzKhmy8ZlJ2Zu2wVxkvi5j1j8dChSCk0Bgy8kLAUQTyfC7/Fi1QYnX8RFjfAE6ytDgg3EMRI0YWTHZPMR/MEXOCSzVcQI1N/NvAOwEhcr96L44zVnfJIeAQcAg4BBwCDgGHgENgDyPgBIs9DLhrziHgEDgwEUBsIB7Els3tuCbZYbKxHE59ydnn/fwH3/oKhREfPnf1Ndel0+nUZz/8vrePrYB4CXJD7ifKyosuNyj/o1//5RYsAS4+97SilYNN4vOrero6cT8ybjr62BNPHh4aSq5QFOyxBdatWbXiuJNPf/FRx5yw8MF7RuJYIFZ86fs/+/VJp734ZScc1FRear2A+IHrKdwtjdcY1hVc3567qJ1hNd59xenuxu2VFSQWnHDyaRdf9s7Lr3zrxa9+zSWXvYOA21g5fP3H1//pZ9//5pclHlzdtmrF8oUveunZBNS2LrWA9KxXvuYNC0485fSrrnznpf/Gr2qH+I2OZxWCzqxDRgKtky5+yzsvn3/8wlOv/dG3v1bqroog3MTPKBWndjRuS/iqDKwgJOdut6wQOQ9xSeB1XO9A+kNcsWZwDwSBV160qFCcgGI//EStqT01Zia+TpF8a+TeqVpxKzy5bMqmTfwICQL5tASLLhOuldP86iGJGxDDuNqB6Oa0LkwZAoONiwCRyYlv+boPieAM5HRf9fla3uEKnoWQXGmC2mlmpkKjzPw0QmCf6bxxhVn1qb+YLQ9MNrHQqWJpTza54aQQ2iIxY5N6Sp1YBfAJIQeJDY6MCeKd9jldDNFNO63KCDUQ+rcJF/bvkxIudjvmqveFSIwd4phPyHuEBoQI8IGEJDM/xK+w6w1MsGD6mzJrBHcxYEXCXRPxYXABhasYTmnjfg3hI6y1a+NWPGP3ZaPuoGgHKxCCSBcTFUk8MBHlnpyJtKWCBnn8oR3Gwzrhb10yfbNWFcw3ghvzypgtYS7bAhOEfTN4RHUoc05TZMpZTeGGSQk/npCRAp6VcnkT9OQLS/6xOffo15/KbN6SLpTngtA8Ud/TteZXJU35xpDJtZ0Qum+gP6h6fSaITprhr+7ImsjkkCkMpoJY9O7c8RVDobKJR4YWL1Ew7zzmURI1NshV1NJRrIpuebBusuPczmfp/CH2YddwAu6f5Pop4ocUYDuvoepiOBKTlUWs3Q9FEmquX/9cWIEJsQNsii6cxqQKCQAXDvfFVygHA50SCSXiycpijmJbxD2/sE6YhDLDkajK1cmqYrw67EzhKk5WUB7tIYrZNYNQYqcSN1A5P1xgvtbIqmNDRd1QWPVOGu5PxCKxrBw/5adWNgxWqVxFZ1vdgNxWDUgk6U8PRh9QwO9U1cSBufFwYaLuy++VCYUi5siymiA5aW4+k8+ZdemkVyhkTX1/h9/cvUEe7AjITfAOoOb/g+LawlXc/crto+6hDgjRYszcF2OnKG9v7ODEO5x5RADcX96JO9ly7rZDwCHgEHAIOAQcAg4Bh8CeQMAJFnsCZdeGQ8AhcMAjAIH+iIjyXQECt06IBe94/0ev4hS/NI71b7/iw5+aPvOgg98v0n28WA+IBOsUI+L0l537Sk7/v+ScV74G10Vve93Ln3YyUnx+14te9vJX3fb3G2+YPnvOIRdd9l/v+8vvf/WL//32Vz9P/2YdfMhhfb3d3W9+x/s+eJpEkze+4gwbZNfc8Ntf/uyCSy59+1Vf+95PvvOl//kY8SDe+Pb3XInI8SMF1R7raumQw4+c/+iip1tqWByIN8H38dxf7QpW45V54K7bbyFexce/8M0fbJZrqDe+7b1Xfvx9b33jpKnTpuN2qkExQr743Z/9avFD99391z/+5pfU8bc//eb6l73igtd/4ktX/+jGP/zqumkzZ895zcWXvh18/vira/+3tB3wO3bhqWecfua5r+T6a9542Tuo950Xvwpf38WEhcWdt/79xhfLouPSd1/5kYnNk6ZcoPpWLl+65Dtf+jS+v4vpkre++/1XfPyzX6H86886ef7OhJsSsYLHi+QvJ6h3VxIhj9XG2cqnK7cqY+0AGcUnJGOnSL2EcrVcP/WZ8oOipu6lEiteEjXRhrysJvpNvFXUbsVGE67CkgLXShCjEJmcGrexJDgNDSmOMIA4ASGOkMAJfghpYg0gHND2SrGY1kIC9yTUAYkeHyU/qfsTxb41nP2Y8r0mn6yUBcawWfuN283AwzmTG6wx3X/rMOmhJlHXCBWQbBUiNCHjINYh3SGv6SPkLaAioECuUqZ1tAzPIlzcITJ5l1yIqfxembSWEGf4O5A5J/MbgtKetj9X3xGSyHcpM0fMC9gzHwSKhuk9bxQn8MC6AhwRLJYoI1RSpyWnwS/3LNcsfeX5/1M+1YJaVFrUC7mDuuEmuYNanzYSEIr9QrCwMS/ok3VBVGpJQjk7dkWaNn3lYS81vzbU+I4Z0ZqUwr7XR70o1hTJnEn3ZoPkNaszq+7qyj0uy4r7+7JFAQaXOAqs4h8rPWPzsImHJUy0PJI/YkhWE6sfzh9Zc2r49rsjJjdldaG1qturrZGgEZkTWh6e5G0MdwQTOjYVmkI65B+f4HVgJYGowrrfmVgBBGCCoIg1xQLthxcToyJWoe0ppl4un4quoODjQ9FoNhSOVkrIrdAFhEYr1mFJAzbsQ9b72NQtixLm8RgJCPxbEM5ntTe8otUN5VVf0RXVTpJG6BXbYC2wz8DOWomxx+gTfZksVAO5ofIlgoQUm0JCg8J+BN5EXE4hjEggyUqoKFPMjKzuyyIl8OS+6qUKzJ2qbBzcOBLPu/g+4UuMV2QkEfSFcuYJxbC4PdnlJRM12c8E64LmAoHB9X/FJVN8TELHSEwW9j/z4Em0OGAsLUomkf2D278fKPNOfsOYCUaEZC+yJ218mp0tAnffIeAQcAg4BBwCDgGHgEPAIbBLCDjBYpdgcoUcAg4Bh8CzRwAXRQSe/vYXr/rortbyPx9412VX//x3N/73p79yNc8QYPsdF73ypQ/cfft2XUpd/cWrPoIVBm6HOjs2tV9+6etf+fAD99w5ts3vf+3zn4LM/9/f33QH9xBACIpty8kgou3M8y648E1vf+8HPv/RK95Z+vxjix64F6uPN77tPVd+9lvX/IJ7qeHhoW99/pMf+sl3v/7F0rKKMV6HW6uuLduPDYFZCM/0dHc/LTj1rmI1ttzvf/nTH510+kvOeuWFb7wUK4cvf+pD7yOY9pWf/MLXKfvRz3/9e9/76uc++ZPvfO0LNm7G7f/8259v+8eNN5zz6gsvIVNuyeJFD1z5tksuuPnGP+Gzf2u67ppvfx1rjK9d88s/cBHLiC9+/Mp3j+3H1V+46iPz5h93IvPBPVxsXfGWi85PCzBb9sTTXnwm33GNhdXHjgSLEjdQhWdJ+O4QUpHwkHTnK2NdgRsdSCrIakhUiLs+EXqTlMOmTHG3qxYkTO0Z1bKoEKUn8SJUJiEjs0TBsyfKCkIigw+xDSlJXdQDmc2njSPA3yCcKMc1E6Qr3DMWHIgHEJjECaA8J+GtyxtOw/McBCvBvyFAIcchoSlHrJi5EisgPzeYqe8bce2UT20xg0vqJVxsMKv+e5kZWHKiohNEREGPkLU6Hq9PBBLatQQ7fcIChD4i2Nj4DPRrgvC6V6LFIn3flxPzw5gRacASDBgzc0aMCkhtCPQ/K2MtAdmMJQqfzAOCFEIFc8oa4WQ6ljgE4gYv5ov6t+bnuHatwMSaLKbiMXBdXZ8OchIcqtK6gNeg0f7RL9YTYow9Kc6Y+E7/ioIUBggNMS/80omR5nnVfuzUxnCF4lb43ZkAYj23crDQdf26TPuS/sKah3ryy1KFoF0up27RPd5bYAZe8kYl86LAn6b6Dlplph/WYtY/WOP1ZZYXZjfX+V1PrMxPP1TlFNuiP9cXVC/eEjQ+8bvsqzYdG3ognAiG03Il1V/r9YDj06wrxnEHxbuT/s8Dc7l6elM4XnZaoqq+GFzbkz+kSLzM5NLDWFbkQ5FoVpYXI0GvPVmDjBDNuEMDG9yhEaibfQVRX5rYGw8qI0qAHfMut2zF9wN9RRjYlQQBzn62rrmYOvClfdYRc7ZC4kg2m4o2SJQYrJ44sFKun9iHx0t0qSC2RrKnzETj2XWZVCSuMvX5TOgkrSlZkwSdXqiwIlqWpV5reWKDw/dKtNgog5MgVhGkWo/JTZGlxZJCxmzYsDS8IK+wOiUJXHE7hqUQrvtwZ3i78Ge9PM3aQC6jdmXs+2IZQOFdgDi51TVlyUDYg4i9B6L1yb44n67PDgGHgEPAIeAQcAg4BPYpBHbfscx9atiusw4Bh4BDYM8hgMuk81570Zv/oCDWzySwNEIHhDeCwKMSCsbGZRhvBFFF7Bb3XdMjlWCstUNp+UaO/E9tndGtcrhDKr1H0O0jFxx/EhYIuIYar53Zsow4SHE5Bvv7+4gNsT13RocffczxK2UtotjTEFtPS8TCUHzvoxEHngk2O5s9EVheqyxSUqmhIcSemQcdcui3JQDJ41P8/W+96PyxsTZsfViENEyY2LRm5VNP4v5qe+3gcmvmnEMOlQHM8Monly7Z3twgRMxbcNyJuOB64tGHIf22SVOnz5x94qlnnJnL53MILTsKxD0ab2C3WlTQGRHvkP0IBa9WhniFkIaEgnyGvCTQ9mLluYodkTbVx202dWfMNrHmrCk7VG6fahskEKRkYbHIhKqX6cw0xCfiAWQXRBfkNsQWFhW0xYl0SE9cwdjT7YgAEJmQmrRp/duX/p1iWUU+IYkhJiFs8ftPfyFbbZwKiHLWtXVjRF94ZpPEi26FGBgyW/44wWz6hdrzpprueyLqiRz8F/uFfEF5iFL6T5wLiF7aYh0jxHDiHLHj/yk/ppzZl9xEjQbaZjzMCaQ+2CNagD3xIV6qDEENHggSuIdjDRSDTStBdJ+mjEWMtVhBePqNMpZkYG3diEFSp7QlnxOxKZdQzC/uubD8uGq0H0YCxVC3VmJX1iz6wYbghkcG5BIq2OruiTFChDN/rDX6wNqi/+VaHLWJkJeWFcXQ+2bHGk6oD1UOKejBlITv10Y8+XcqDD3Yk+/766bcosf68ms3phTnIDCIwMTmoC7qpE+IfawXcFqr8/pnKpJDc6U38Fc5HOqW9cXkMjPcrxgX5Y3elvBQUL7QM4XwFH/Dre1B06LXR37dNddfOvRUYdaWd0a/n93ZWhJ5TrsITKzv/5IAcV4kVnZqokZbUa6fioKFYlUE8qQW5HMP+uHozFDIl8soHxdZRYsLJdYyJDxuzpjHhcqsA2uZgOiH2MMe+Kky64P3BHUwVhvngL2+swRWiFhY5WCl0zraPq7FeN/wrj1ptBLJ2IHibWRMvCKdkSVFqLqpX5YWISGYMBIoZEGSvjc1GDs+pd8aC4JaMlaeWXnI6csfbJjWXabniUOB9RZrkPEgLPE+KLqckwVHfz7rDQ12ex33XR9d17Ey9A5d3+q+b8xgLtPvn49e4/20jbqxvwkWJXEsGDL7B1y+pnyyMvum1O3XJ/UbMXOpYmBsFeLH4Od+OgQcAg4Bh4BDwCHgEHAIOASeMQJOsHjGkLkHHAIOAYeAQ2BfQuC811z05g9/9mvfQYj5zbXXfO9zH7niv/al/j+ffZVYAQmMmxdiEUBIIjbwCeGMEGBPKK8VPTvF1J080bR+uNpkOvolWKw0FfMlWFTK/VIUEg8CFIIb10EQofzmFDanqCGJqYtPyGNIZO4hDPC3CCQmZHmpKGHd03CfDOlpYw3wnWvUCYlIPXy3QXz5jjDCGBAWEBn4rdgaOjXvefSzV4F2N5j+h1rM0MpOs+aTG83wWvHMqZPVC8XZKOJA3RC2tMupdKwHIGsZE6II7pOwVCq6PxLRvE+QdhIswAmiuVWZuWB8uDTjtD5kOGNkPiB6IedtnAowZ7wrlV+vjFjzF2VIYeq7TRlimnkGC+apaLnyTIJsjyFN9XhxrjnpDam91RqMxVK0rkiZf3Zlg9zP24NbHh805RoM/aVPiGWsI2vVw9iyqsxTUO3aWRV+4qymSK4i7GXPbgo3YWUhYSIpEaNo+fX7Ddmuf23JDbQNFdbq3D7CFeua8bFvWA/WZRbCLusF4v8mZQjwCVpMbcoVCr69IVDk+TIz1BP10hVdQf1pgfEUjCW9RKLGP5u8zVtkZbFxwFQMfDf+3uGdxa6QYMH6ZWzM3Re1ni9MVNaZRE2jCcfiBcWusK6WUCcGjVfoj1Vk7g1Hg1PlVqk+J1sO3eiUxQKiBPsU0QLrJAhp9uU2wbeBQhkxBjdQCFn2/g5iVoDg1sRUISwggtJ3nqdtrllLKes2rPgQbpz8cH5YsTIKimmRl3BRJZdUtsJf6csrGITyX+UCKp6oSuVmnbj6qQkzOuskWPAes31knuw7gv3KeHskdDypp/1kj7f0b19N9A/3e7/fjhMu2vqwMuuYPT+uu679RbgYs/dYR4hUH1Fm/xXdII5JvDdwGZeUaLErbszGqcJdcgg4BBwCDgGHgEPAIeAQcAhsi4BzCeVWhEPAIeAQcAjslwjEpFB85HNf++655194yY+//ZXPveW9//3xJx59BLc2LgkBiRUQzG9ShjCE+ISghriGlCNB9EJgeqLq6kzjaRWm6ZIhk+3tkNunQVN94rBcP/F3BEQWZSGVISFhFTmFDfHJb6wRII9xIQKpO1/ZCgs2AK91Q2NPjds5shYSlgiDQOMa5WziGmQnhKK9R7v0AeKcDME+ElTb8yCeKTtXlGiLqT6mYKqO8Uz9SwfN5p8dZ9b/IGlS6ytNNtmv2hKi7xFgIDzpO2MAK+veBmIUQYPYGouF6f17e2yLUUsd8IPQBRPcFEG8MxcWV6wqsJRYowzhS1lEDESII5W5f4MyxD1WGsy5YgkUhRzWQ9GqQpl5e06WFXqexByzRiCptyYsBeSaiVSxYtg8siZl8lrA9BFxijmywhaWIc1aHNGIb9LTyvzGOZWh6HmTwuGTG8KVBOkWxR+SS6lgcyoY/PvmbHqJzuArTsUmWWuwlhgTxC17gxZxGQRZz9qGBAeri5SxTIH8L5LbBeO3SZh40XBQNhTxMltSJt5Qa3rasiZ6X5+pPrZgvJ5UEO9aHszKbQka8lXeQDbRz3Ia65Xp32OWWMEaR4BjHk5CrPB9X+R+GBdQgYJp/1usUAEpMxXyCLWiqnGoGzdLsbJMXe+mKoI2VOh/ZPli0iL4OxTY+knFc+jXJ/tlrGCwBkc6AAAgAElEQVTBWO01RED2NhYMO0qW2GcdsEbYo+wXRB8wZS+Rt+mvrVBzG0iguFEZMZP1RpBn6wqMuUCI7FLf74gmsnMnH9q+qW6KPD/5AWuStWzHwSeJ/iOYPKl8pMbdwv5WQO76uWdk73jqrvA3h3r89yo+h7VA4Zk1yq3KX1HmvUHMIyzlWFsHQuLfA6xgCEC+zd4rGTzXEWytQHkg4OLG6BBwCDgEHAIOAYeAQ8Ah8Dwj4ASL5xlgV71DwCHgEHAI7HkEps2YddCXf3DtbxsVYJvYH/RgRLB4ulumPd+7F75FEeu41Tld2QbExhUUpCxEK6QgJCMnyf0i5Vt3TGBaLu8wVccmTbwJIpIy1gUTZSGoISQRCSD0cQHFfchVTrvjZojT1NbdEwQoxC/EJyS5tZwAHCtSQGRSxlpYcK8YaHz0Gr/5bl1E0b59hnZ4DuIaYhdyk7asiyqI+mGVoD4CCHebaN1CM+XyR8zEN7eYDd/ZYrpvCUzPvzYronNEdDxkKeXABwEDgn6NMm2yvjh9Tp1zhO3NEi0epnN7Wxp1BQXeEN4IVswR8wUpjDUFxDvYcYoel13MK6IVliVYxkD6sk6wKMC9D2NmLsEXot7GdLBiwe5yYQYBLYGpKBQUkw2+wedQIbhn+ZBZPJjfaklhLYP4O5d10FYW8jKHVPmTz2uOTD2qJtQggSJfE/FiFSHP25wrZDvSQTpTMAOyqnj43u68n8wFmA2xXhg75DzrnvGyjtk3iDOMmWunKrMn+I4AyK4BY3mQ8hrTJlqZD/xfa6NMzphpA1p2D6aC2OyUiW3MmxD1N3UHdQyFbOK/f3rIgNT5NWZUrGBMEP+XKs/z5fopWlYpsaJc4oTsRsYmBaBWXI10KJIPWmZt2ZyoHi6kBuLtG55oGgzy/jK5W0okqlNrB7vKN/Wsry6X26XZEi4KEi7ohA1WjiDH/rH7lvEzRvbeeP8tgYiDCzHKgYndt8wLewXszhjtKiIQ68WKEdfpO2sUN1unKd+jzBotWnPImkIWI+ZRWYekQ6FCd3ldMjbtqPXrJszsrJA1BmuXdw9rljoQGYnFQrLvBuYR8Y13VZfgS886MRdtmFboWHlf+O8bHg8dmxr0aorh1EfK8G48Thk8/qTMvmGd75fWBLKSMGOsLMDrn8qITi8axbL0gz3J3kSEAneXHAIOAYeAQ8Ah4BBwCDgEHALPGQEnWDxnCF0FDgGHgEPAIbA3IXDKi1927ueu/vF1a1evWvGGc05ZQAyLS9767vcT7Hrl8qWcBD1gk8h0yGbIVVx72FPPNkCxPTUM8YQIUSNKLmb8yMNm6uWBaXhZnbzaQC5CTllrDIhkyGpECchJaD7IPEh9YhpAeFMvxL4tA9EJmQgZaq0imJNS0YLflhC0JGypUGED69o4AtRl67DP0S7jhRylL5Cl1hrDiinUTR/AoE9E6CQTqW0yrR8bNPVnr5C7qFrT9ed6037DItGycfVoispAymF1UOrz3rqcatX1E4QzZVZIuNgd1gWjQ9stH2DAvBctDpRtEGVIeAhZTlNDFFOGDE64hIKYh4jnFPUTypx4R7SAmOZvSe5DbLJuiuvombiA2snImKNwJOTVx8K+HxYn35/Om6ykAAkMhhDLnRnTviUTpHUq31qNMD/MaTSkOM2KSdF8VlO4/pSGcNPsCr+6OuqFZZlRWDdUyMuSInhyoJB/oCe/Zc1Qofu+7lxUdVr3YhDWYMDYWN+lcVgg8C0m4LdamXUOgWuDFbPXitZECsjNs+W5IIyFEaf1wYlrNtg1RDvtjFDlO06scSwVIopP0RmOJRoicRkDhWSzofgPEhuKGakmEpc9h3Lr/HV1FXXJSSL6vaqJA7Mr6pOLhvsSj1Q3950WCheOk0gxlOqPr1/1wLQtA53lh6YH43UFwpGPpFZlhBXbR27QTxvTZGxvER8YI9ixT8AF/Hi38Akm7EvuI4yyX6xggaXKT5SnaiwKfR4cpXGlwrHcOs1vp4Jrd5XXDT1YyPkb66b0VDcf3FEZTWRiKsseZE5Ym6xla5lxvb6frVwqnlKO8pR9IBoPKhqm51sS1cFQfUvh1uV3hs/q3ejH1V6pyyveee9X/j/lPyrv6lyNxWZf+81a473P+h4v8R5AzAxL6PCcW6h9bXpdfx0CDgGHgEPAIeAQcAjsnQg4wWLvnBfXK4eAQ8Ah4BB4Fgi85NxXvebzV//4l/feces/rnzbxRcQsBwXOF/90XUnLn/i8cX5XO5AceXxNPREokO4YVlB8FQIVchdLAEIGgy5a339c69M5HxKlOQqM+ezy0zjKxolVkDOIlYgAkDk8QzCBKevIf1xlcJ3GzuAMjaos3UbRL/sqXcIRIhMK2CUChLcs2KEvV56ork0hkXpd1sGwtmO0QbntvVBmELA0TYZ0pIx8T0yGng7ZqqObjJlB6VNvOVRiTanme5/RkwuudEUclWSPSBveQYLDhs4nDYh7kasMXSSXJjfKtECYnlvSUXyf7TvkMX0jSDSjIf5h2xH3OE7hDJlIZK5T7wK8EWwwC0Q90k2zof9vbusKixmRSuaKTXxmvJoqFE/8g25gr90y7CXKQTJzRnz66VJ09eRKZLVnH7HGgIyulAe9jxZUyQOqfQbT6oPl/flglyIkM6qpDMdZO/uymd6s0FEwkVasSoyXZmiVYW1IEF4Yw1BfNtYK5DUjBchAywh8C0Rf5u+W9dq1grDusfi97HK7AP6xsl/6gR/5gEinz1kXZ497fT+qHUFa4x1jPCKe6MhuTaaXchlFEbGJ0i1KasZNsmeMikkvimvHTLxyvTaysbBlASKBbJOmCIpgz1bo98n6P4GXavXSOao4lC4Pnn0tKPWmc419YOblk+IpAZiWb0+bcBy1gLiJOuBPUX/t5fY+1g2IXDxPrCuxhA4WEuLlFuVsV5AsIH0ZkxY9jDG2bII2aLx+LL+WNXQ2rVIYkpZKJqP1U7SLBa8+lA0t6SyIVktMWOByrOfmQvcmzE31q8WogmYgz994T57c6ky80db7fp2pCwtKivqCwONM01XtCz48b2/jB6fTXuIS6XpLP1gznCRhAu0AyWxtxEsvqFMEHLWBOsVsQmLGIKmB06sOFCWgxunQ8Ah4BBwCDgEHAIOgecfASdYPP8YuxYcAg4Bh4BDYA8gMPuQw474zDd/eO3ih+67+4rL3vCqTCYNSWVw6f7PRSsW3viHX1+HeLEbT37vgVHtniZEnEPanacM4QbhCLkHEQtJb90n+aKjIaCW6Jj2RJOY/pBpODdnpn0AEhvykfL83WCJeYhbiEmIXYhIyD3IW2vtACHIfa5ZN08QnZCy1kKCAULOUhflqAuyHFIWEheisxgoebSffOeavW5JR3sU3J785nnqs2IHpCmkJs9TP+NnrLZdyHjKQMIiQoy4SQpXpEz9izOmZuFaMyAPSGu/HJiBh+vM0Lpu1RTWqLAswHUS7VIXxJ7FA1KvXNjjZmntzgIpq8zznrT2M9oDVuChv5YoZuxY3XAann2zZhQ/cIekh0y+VRlxy1poEBcECxowtgHRd7dYASZgW57KFuaVx0LNspgIlUVDpqU6Zp7oSpVrQEcmQiYniwkCXtMfrD7yVRGven5NqPbc5khIHYw2xb1YLORHVDC/JBnk5PqpJyVfSfd359Mb5CVJBhvF4OCjc8hagfSG8Gbd8xuhhr3A+mfMrGHWDUIEwcCtZQTPWAsLhJ3TldkfuEJC1LN7BuEAbBkfa5K8o8TaZW8hNL5G+WP8ZjojZb6pbOyXYKEtHHj6PmCyqYhpPnjzQGV98lGR/sslTJwwWrm1iohIukHARGgpCnD6PaGqcTCdHoxtHOpLTCrk/SAzFLUxHXhvnDY6TtYDa4drrIfxEsLXMmXWmRUsGAPvEnJpYuxgBsYt6mt5TXP/9XJXVVnZMDihumngEFlUhCKJbK2EDDAgdkiHyoEd+w+h6t7RT/YgmX1sLTdYE+x5+kp/mCPeZYhbuHtCzOhVqPVcZWNhUybpZWOVJp9NF99pYxMCp3WlN24A7nGe2acujeMWin3B2ifzXiMxp+B3iTL/jnTIwmLQiRb71FS7zjoEHAIOAYeAQ8Ah4BDYaxFwgsVeOzWuYw4Bh4BDwCHwTBD47//50reymWzmw++69A1WrOD5gw874qi6hsYJCBn8PtBECxHmkMwQqpxE5sQ3p6QhmiwpWyf6lVgV/frftabi4KRpuWKRmXxZnfz6YDEB0WldKEFSQU6RrI94BA/+noCItS6QbBlL7hZPyStbYcEG2uWaPZlPnZSHEIRQhPjnNDqJ7/QBt1L0nfr5TR9KXUaNFi/WQ7ZxAay4Ql8hGbkH6QrRaf8WggTlhDdlIYVHXNZ4YbnCghE+LGemf6zS9NzeYTb+JG4GlnSo5SZlBfIujhuiH8IcfKmHOugbJ75v0zw8LtHiBbXw0dpn3IgxWCNAPIIhhDv9hcguurJSxjUUJK515wMxTcB65pg1wXjBjTIQ1/nnUQhkrdRuGkjHh7P5WHUibOQayshSwtTEw6atJ7v48UGzSfErSAMxlW4t9ysvmhqdPrPcr03lTbJgAq8vG5h0OiisShYGN6WC6O2dOa87E6SG8oECNmxdt7Rl1zBEOOO1sRwQLphP6/rMuhhiTVkXWwR0Bg+sBojbwn5jn4ETrrU4nc8pf57FbRXrGysn1h5lbKyH4mDGJPrGvGEhdblyQgS7icQyRUuK+ql9ppCvHu7dUJeomdxbiFdkBmRdMRAty8yQFYK1BsGioTRNkMBxRD7r/0JuoWZIsHiRHy7UKHj1QKHgZ/VQbWdbrclltvnPBfbFcmUEBsZ6ynidHR0Le2DcoNolz6zRd/bhLGXiUzyufqysa+l5onF6V4tcQZXJpdVcXc/JOqStuN9G1h5iAvjRBvgjyPI+sO7JEEF4b9BfBDneHYgYrHkwRKBCFKUu5qXoAi0cMbMTNcEdjdPzmcGucJveWsx7aXq3frDXb1LGOmlHliZjHt1nf/JeYP2C99j5Pk3XsL5A0ET42tvc4O2zoLuOOwQcAg4Bh4BDwCHgEDiQEXCCxYE8+27sDgGHgENgP0GgafKUqfOPX3jqb3/xvz/o2LQRsntrOv3Mc1+JK6j77/zXzZZUPVBEi1Gx4kyBAWEHUQ25BzFKEv9XJAkHTKi8YOpP9k3jy/Om4RVVJjb5BN2FBCQ4rQ2uba0jeNa6rLH+6K3bJYg/yFFr+UBZiEHK2785rIhgLScsoWljWNA/iEUSRNkaZUhfhADIQXzcl5KI9vS2PeVvg3jTpq0bghECE2IUoh6Cjbpokz6DEc/RVwhOCHobSLxRws2TJlwTNhXHeKZ87rBcRUXM8Koy0/aFAZPe1K3R5TViyGDEFghsXP6AAXhDfNM244LQfiET82WDQ9M/Tp7zm3FjLYDLLwhh+m/dvoAL5DoZIQMsEX3Ah0/EiudzTMyhYi+YCX3DOZOIhEyFVAnNhgnL3GJBOph7e0/uESlBhea43zSrwp+2sCE0PewZb/1wYWjjcDA8u9Ive2KgkLmnKycvUia0VrErdC+m79RtRRfWGPPE+Nkv1qUZ40do4p4lyO36Zx2y7livPGPFO7DjOX4TnJw1wLPzlFlviIisP9Y0dXHNCneeAmxv4xJq1B0Uz1MP+NcDeaJKoWVa6dqAiSW8nrLankHNRap2Un8oHM8GsbKMH4nnIrJKgNxnjhGjIOYR0UiB3Cs1SLR4QzYdrpZokffD+QE/UmhXrzy5XWqtbEzG+jZVxnSHtUNi3hFiXjJa1+jlp32wKMBkZ5YjrTwpUWUgVpG+vqwqtTJRMxxpbO3KKkB4j8a5UpYUWGvwXscCgxgr9N/GD8E9Ey6eWMfWWoX7iBWsWTuP9BmceaeAIfONuMGzfLJ/y1TDGuH68OyTci0dK0MfT3Z7Px9ngLhFQsBjjvd3wYK1yNoBL4S48RJCGoIQ68sJFtsByV12CDgEHAIOAYeAQ8Ah4BDYdQScYLHrWLmSDgGHgEPAIbCXIjB1+iwILfPU0iW4hdmaQuFw+OUXXPSmh+676/b+vl5LghcDAu/vooXECk5yv1kZQpZ/7zkNbYUL6yv/AQWZrjf1Z003k96aNtXHNZlQHGIU8o8MyWdJ/1L/+qVWDXy3J9MhasdaU1iXQZbwtIIG84QYYgkxrtNPiEMIMEgyTp7Tb57lZD8kJCferQhg66Z9cinRS302boVtxwosCDXvV/6VMqKCjclw8Gg9kJxYcXACWySmR/kn1YKuldeZhnN6zfDKQTknCpv2a28zfQ+0mEJqhu5DUNOGjWsBCc04ILbP1JxAsv6dfsnaYo8mrXewpX/ML7jAdCM4QEKCOXEFIHPpI/PIfQQWG8sCK4w1o9coB/lbeJ7FCjCybr6mMLkbB9LyWOaZhvKIqYqFzPyG6Kw3ZP2apq7C+gW1oaZH+vJlNREvVinFQpYW5TG/EFnan88kcya1MllQoO0gM5wP2BPUC9ls3UDhoglRj2YgvBEumH8wAweIevYPwo6NkwFmCHuWDLcCBcLOy0fb4DtkLriyFsAW/HhX8R0i3q5VxruNWMEFJdYT64q2SRU8oVgLpn6aIoQrhHh1cyFbVpPyKick1+pWVTianyhLhYRedRDN7CHWIAIdpH9SVhNbhvvilaqnIpsKT1DZkGJGBPGKQtz3C8kJMzvjNZP6vL7Nldl8riUY6KiI4m5KCWx4327PFdRoF7dia3/bT97DCIdbkwJpG8XUKNRO7jtR1h3Dajfj+YW07wW++kc79B9sL1Bm/+PeyQqPt+s7AttCITdVOou8ZHmPZFKRm6KJ7H/qelx1RSV80C4CAxjingv3Wf+QYPOgMDpI42c9M67GyEgQ7tbjX59ed+sP4psLeQm3284KfWE/HCj/HcXo2Q9jLXTsHHK91M3f2Dl3vx0CDgGHgEPAIeAQcAg4BBwCzwiBA+UP7WcEiivsEHAIOAQcAvsWAsPJQYhXU1Vdsw0R9ro3veWdWF9843Of+O+xI3oeXdi84OCJGId4xT89J6ttQGVEAIi/nMi3jGha35Q1H2xa3lNjGs/3TEJ8qh+ePEpKQZBCwkLmWrdOVrBgfKXkFIS2LQPJzfdSl082hgXPWXGCvz8gb63wYUUM7ttTy7SPhQfX8J3OM9zDigEiGcLSuuhBkKA+2iaVihVWQLGiCvcQI+gXpDLEsY2RAZFNvZDTtEWb1mc7Ln5G7nsKjBKf5pv6cypNuHamiV4/aLpu2WByvXIfVSRUWYeQqsR5sDFCIEOZAxu0t9QV1mi3d/+HhAoqZRw2yDinySGdId0RZphzRBsyfWcOwZP7iERYo0Cwgx/zbgNEp/fQHiqNGWHy6sGK7rTJ6HNSZcRMKg/XXjw99K5TJgYPKUJ0anVStgDqWEhU9+K+fPauzrzXniqYobxJrUkWwnoO3BERwAPxBgsAxoxABwaMkTKsATJYIGZQHvLcWs8ALOsBCwrWKusKQp3r4EhG4OB5AjS3jtbHNdbcYmXWlBXT6MP2TqezVm2cCyyMtAR1oTwwlQ2BYlcE7fHKQreIdpHo+Vnqwcg+GHFVxhiI10Lfme+/FwpeX297FfWdkx2OzPBChVgmGTMDWyqGmg7qKIQihSq5hqqKKUKIAlunJF74w30JxcXY+p8NkPU7S6VWVqVlt3lHSygw0UQmnahKhWQJ0jLUGw/kDioh0SSey4YlLATNEmQ6JCykim6hvADriHsRY0Yx4Td7a6oEiEw+F6oc7CqPty2a0jhp7qbl8fLMXI0lG4lnH1dm7XZIqGlLD8VmdqxqqOxaW3twy+Ebp06c3TFFAgf7k3lTm2behJmFuTXNhS/0rPe/PkZF4j1qhSoEIRu/ZGeY7Mv3GSMxSU4fZxDWlZl9/+7L43R9dwg4BBwCDgGHgEPAIeAQ2AsQcILFXjAJrgsOAYeAQ8Ah8NwQWPrY4kWdHZvaz73g9W/86x9//UsZU3Sfc/6FF7/vo5/+0srlS5f888Y//va5tbBvPC2hggQZjViBFYJ17wO5B1EOtUawaFHnLw+Z5ksqTO2ZNSZSBeEKaQ8xCsmJJQNWBaSx/n4sOQeHB3FnLRFs0OpS0spaX1DWPmfv26DYtg3KWHGD5yAiESzoG0Qyp+Et6U67VlCgrCWJbcwLfm/vbxzuWTKV+iGNqY9rnMJG4KEeyE1ISfoB2WvdXtEXxbaIhk20caWpe1G5iTZEjR+pNBt/1amedKsm8IMoRqwggS0EMaT4i5S7NFfL9lAgbmvtQf/Bkj5Z90bgzZjpH2Nk7IybE9NgwlghZLEwgJxHGCy6gRrNo8N7Xj+YRwSTNk3cPCYPv07Lu1OmMuqb6njIS4S8hpYyc/w/NufveNGEcLNux/+8Kdu5arAQXzZQ8GRRsSUXFPvP+rFug6y1CeIEGEHmM1aEA9oDD9Y05cED903MK+vQxkVYqO+sZ07t8wx9Je4HgiGiCOQ3bqDsXrFumcCZdcUn9bFW+F3Yjjso6rWWT6xZE2g2U4Oe6W33TfOcfCQcDaiHvmA1gasv2kR0Ys0huCCeMe+E9KgLhfMLFVh7csfKhlheMSoiiYxJ9SfKymqG84qJMSzxQMKmZxR0O5zPhlR/zuTSYRuAmy7sKFlhEhx2mCRGGLl+inmhICrRQoGvg2YF2H7QiwaVPRuqAwUAH6xp7uvuXl/bVsh7nfVTe8ryOb9N8TnWSVCRNhUgDJ4uQaNPViPtw/3x1g2PNx/d2159sqSr39dP605pDIlILDujfmrvJhlg9K5+cFpjx+r6N3mBmSM9b2DV/dN+qs+HmudsrpULLSxeEEWDUCSonnFsbvnDm6K35rPbEPW8T3Ejh7XKdcqsm/0qjRN4mzm1sYnGjrVNF+z6369wcINxCDgEHAIOAYeAQ8Ah4BB4YRBwgsULg7tr1SHgEHAIOAR2IwK5XDb7icvf/uavXXP9H/5892O4ESomhIuPvuctFxPDYjc2tzdXBal5sTKBsiGeIZ0hTY8RfQnB3y6XTxEz838KpvG8iSYiF+9+yGJjrRQgNTl1bwNal54ettYKYABpbS0ZLDEJ6WvL2JgU1hrDxsAotaawYoM9wMzfJZDHkMOcxKYP1tKD/nHPEv/2xL+tjz5Y90H2VL69R3/tOGwZrlEHAg9kG32gDTCjfYh8e+KeU/XUCVYQ2YqQgOVFOJCFxWpTsWCdaXlfk8kN95uOGwjEnVbNWCdAikNSP6jM6W3qoP9vUv6hRIvVe0C0AFMyfYcUZ/ysCdYHY+Q3cQEgwiG4wRuXOdcr40aIMUCoQ+IyFuohj+e6SJd3e2LesBAQPS8A9T9R5R71YGl3OpjflCjG0MCQ5OSG8Il/35zb8Of27ODSgUKuNxv0DuaChG5BtNJfiFXGybisOAcOCBEIeqxpxAmECu6DBfcg/CGleRYhEMHCCmhYWECaM9+sJzAC31uUbdwJ1gyWOqwn6uI7deOKjLVXjKcyVqzQNRJzp41qXjta7zSsK6IaVeP0gplyeG5z1cRgyA8Xx0Q/mFMEi5uVX69sLWkg4ov9F7mvOoKG/o7KqmwqYmSRQAyJ4kroXlsbkmDQIEEgp4DdhXAsm9W9QNYJmdRgLIqIsQuJ8bPedxa/otguQcPljkq+nCT7RXOMFeHPj8RyrRuWNIf6t1S0qJ+nSDip6Gyr60gnY0MzjmkzE2Zt2ShbpzpZVqyU9Ucs2V3eqM90sjdxuGJy1PdtrnrTUH9iSqw8bWRpMTGTiq7X9aHBrrLTVf88CRoMJZ5Ne2/uWNH4+4q6oRkKWF7v+wHrvU94VE+cnT8sXhksHurxTh8xViomHkTQtVZf9l20C9Dsk0UYH+9AxmsF39KBIGKyRw8ES5N9cgJdpx0CDgGHgEPAIeAQcAjsawg4wWJfmzHXX4eAQ8Ah4BAYF4F7br/l7695yfFHnP/6N13WPGXqtHVrVq749c9//D0sLw4EyER+Q4afp/xSZQhQSFJOlUPCrinSTKFwl2n90OGm6ZIGE6pRsO1IVPEZOIFNef4msAQ/wkMpwQ+ElqmkJhuw2lpFWBdQpdYXPFPqOsqSXfZaqVhhCT/bD+t2x4oipUSZ/dullDijztIypQRiKcNqv1OvDdZNWRt7g3ogmbkHYf2AMi6UIIvBxPrSH3Eb5Xmt+pxiIhUPmOrjQ2bWF6OmbGarWf+tm00+z0n3DcqUQUyBBIf8pt+Q3hcq/1Pz9rhEC0jr5ysxZsZo5xcxClKYtYEVAFiTKEM/wAaLCku4QzozL+DBM0VBag/ErrB40G9iQPQUG9b/KISFCet/ejOBebArd9+RdeEjI74XjfgmLKOLhFxBbdowHLSn8oGMLYriG3uBebWiF/MMyYoIAdGKAIGAwByzH7gP6c6YESDABkEAfKzQgXWEFfsQK04cxQlhAAzlY83cq8wawhKD51kDuC9CqEA8QCwpurNT2p4ARJ8hx7H24VT/ZD9kcuW1QbiqsWAqGoIBxYDoK7p5M+Z+rTfmk7rp5x3Kpyiz/mg3D7kv4WG1BIuJEiFCxKWAuJcYoOWsBdpWZ3TdyFohHM+EZMnhR+WeifuB2mC8u/LfDtu4fRodX+kH9YB9lSweIlhZhOO5lESLwWhZNiURo1rCQv/GZRPzctmUUb86ZPExTa6skkHeXyYLi1OX/ms28TVWTF+wrlYiRW6wszzcubauXp89yZ6yGyXKXKLrU7AKSQ/ETL4uWSuATxnqSUQ0/iorvBRFiMBrlCjyOo19TWXjYMyPZ8EbN15rwlHTLmuW6u1MDgIUOIPJHnHxNg6We+oS6/0mZQTxsQmRjD2631ma7ClwXTsOAYeAQ8Ah4BBwCDgEHALbIrAr/9HhMHMIOAQcAg4Bh8A+gcD6ttUrv/WFT314n+js7u/ki1XlAmX+bYdY54QzJ66hQlMmXF4wE84/wjS/ZbrEioLxowub43MAACAASURBVHJr5EG2QbRBikKyQk5D1iN+WIsIy9VZgYFyNhA2RC7kI/dKBYOxx7Ct1UWpdcVIz0bagRS2ZPJYqwtbV6lgUhojg3rsM3wvjbVR2vfSPpWKHrbf9MHGtuAaBDYkMflhZeJoQC5z+ppyYAVhiQiBG6B+U3HwWjP18m5TfUKrWfGBiBlaK5yCpHoHWc0zfEL+c5r/yNExQwSupuO7O43Gr6Ba2obIhlS0AYutqyjIbfoDGY/bIMhta3mCpQn9s5YhWGgULRr2YKJtyPYTIZfl2kkLxjPyBGVSkk06UoX1ywfyhfqYP60u6k08ri5U3xz3H1sxWHTtA3FuA2szV+DP2BgHggRrj30C4crcsgZZz8ypFbXYI9SBkMFzCBAAgOUJAsRxoxghPlBuqTJ4tiojTC1Rpm2wZ00hBtE3MmvJxg3R123T/IUX01frzo3vrEEJDOpsl/yOtflm4hwvXlZl1pfVBNPVq+N1G4GWsicrQ7rTf+pgDQyIyP+73CxNDEVzx5TXDEe61/2bigdfuYky7csnyuIhZSbM6DISDkz3+hojV0uygNgt8w6pjVBWtPjJZ0LNwwPxkFxRRdU3I9dNSbW5WfElyjtWNjZKTAGjKokUc0fHgVjYKwFlnqwv7pU7q/XpoWhnOhm9R32sUAyLw/RWwZJmNAUSh4KEBJhGCRee4mV0SsSYGoqm5FIrZgoSaiSESJjxFg/1JjZL5GiS+6uYBJ06LfPOsppC1bxzMu0P/i56WzblnTpmij6h3/coE3x9fxYsrBDN+h5vESDW3ae8fOwadr8dAg4Bh4BDwCHgEHAIOAQcAs8GASdYPBvU3DMOAYeAQ8Ah4BDYixDQKX1OkUNW2lgUNiB1VzGmQt7MNFPf0mparphgIo0Z+WFRSGLPumuByLQnxblmXR8xQita2NHyG9LW+jKHGLWWDqXWFJTnuhUP7D0rXNCGDZJNfZB9pf7R7bOlKI8VLuw9236pOMF4bNsQz1aUsM+Uih+lVheQ9vQLops+H6oMwUrdkHWQz/TdBtylXoQAcB8ReuIt/SbSUG9SbdVm3TeiJrmhQ1fLRPNZdz0IAogA1A+RfKjmr0dWFhDXuy2NihVW2LFiDFgQb4HfxygjBDAeyHprBQLhDsFOYGXmZJWyXR88t6cTa8NaphTbphP9Ui6i6nk2m6v80tLs3TKvWPqypsghx9WGWs5uCk9a2p+v7swEWFUgKtj1ZGNvgDViDHNn3ZkxH5D71joHTGwMEuYJnBAMyDaWBUIHiWf/pUyQe2JWcJ+2aQ8RkcTewloHYhcS3rrW4jprcDxsaZM5oB+4qiom4leITN847ah8UNUY+OFYcJBqYBx2LBDojI0+FAUREf8pLCkGtpSfkcuEoiLme3s2VqdF8CdKbTsQDRSU2igYt8kMR4vWFxI4sLSg6e25BKINi5Xt5vY+qQirFsazWe1netbX9EkkSJUpdoYCZA8qwHesq60upH4erDKITNYtGJZBWD9goeKrb4n2JycsLAqCgemVoNKrmBYpzeAEAbrCj+RnhaN5gnEbubkyqWR0pSJ7r4uWZxZUNQ6a/o6K4hjDkbzxw/kFFfXJf2r8vsrnJWHQroQNo3gZwSJZsvT2bhhxPVaSWC+IUwWJS95Dd/5ie1YyO8Nkb7/P+sR1HtY64yXGzZrfn0WbvX2OXP8cAg4Bh4BDwCHgEHAI7FcIOMFiv5pONxiHgEPAIeAQONAQENnNCfmzlSGfW5UhKjnt7Yvmm29C0U1m4qvzZuLFlRIrcvKnowPqntwVefwNYMUCSFNIWVz+QMLxm++kUiEB4gq3OTxnA0lDQELmc53vkLQQrVbMoA5rAWHFAevCyQoiY4O5jrXqKBU+qG+sSGGtPLhX6sqq1PLDPlfaH9tHSxbz25KQuBGCgGMsjIk2OTEPkW1dCEFY0za/IYcROtabUKLb1J+12qQ39JlNvxs0qXWyainiA3mOmMQnbUJgQ3BDwO5WwYJBKtnx2cDOCCsEGYdcZlzgQ7wDiG4EF4hkAgkjyFgXUswNayG3hy0rRodQxBfLD+JqHG0nPqVZHsgHZks6qJL7J39DbyH5uinR5qqIN/Hc5sgEfeY+9FhqcEAxLPQc65Vsg6pbgpU5Yc6Yc/YNlkNgBRbMOZYvzBVluAc5DR4IhKwznkHQAk+eg9QFY6w2EEQobwPJ27atlQ7ry4qFNrbIWMKbfkDaQ9JDoBdTSFenH5vraj4kH5NYUS4B4ybNJgIUlj60zzvBWgf1K+bDo/msf4JcPU2NVWRaZW3QLYuFJbJSuDEzFJGg4m2tm/oRKeSYSdl6TRtxxbWDtDOxAqsP+gMGrEncZWFpwtz0yqLizwNbKrZUTRisVbDsGamBWLJ3U1W3xAOsKsCVxPwjWJDAnzX7ZokLG7UzqyRUJMKxnCerkbbqpv718cqUp5gWl3l+IY7ViKwqhsqqh1M1k/vmKFZFkrgdyZ6EKQz6nV4sxxyXy+1UWnV0ywUW+5z+rlCO5XPe8vqphXUDHb5cZT0NhUt05TfK9yszj/tjsvGMwH28xNywRw+UWFH74xy7MTkEHAIOAYeAQ8Ah4BDYqxBwgsVeNR2uMw4Bh4BDwCHgENh1BCRWWJc0+NCHMMdCAGK1IBIvJEuKTWbChb5pfGWrxIqI8eNyBVUkNK3LJwhDCFVLR9qgyhBvNq6D7ZB13cQ9GxSba5CynMiH1IYAJvGdukuTFS2g/CCDIWvtSXRrgUEZvpe6pCq1hrD1lQogpSKI/T7WZRTPWa7bfi/9pD3+JkKosafI6aN1pWNdInEPEhsCliDUEJuMA0xoE/wgsfOm/JAu0/LuPhOuOsWs/nK3CYbzkgeYG+plnsAMopc+n6a5bJaVBT7id2eibvrHnEOUM445yhCQWHmAP+Og/5x4t+6TrMWFtYghZsULdXqcviIEvAhgiqYuEiqyQrFDMSyWJc1An6wtOjMm/5dN2c2t5X5DZ7qQP7spUpXOm8IHHxuWZlHEnTFi5cIn7p2YL/YM47finY0lQnusf+YaixPmmXVJ8PRWZQh++kV3WAu4e+IZvjOnpVYT7A/mAYIelznsN+YAoYPMfqDu8fDlGuvpVGUsXopJMStEtvtT+jf7bbVT8hWKacFY1igjbjAG3EFBHm9RrQgaGyLx3GCh4G+SGDBJMR6IXTEoV0rT5VJpG7HCtrEDgeKZ+oXC9ZUlum1sCwTVh5SJh8DYuwc6K25dfueMCerXPKHVbwreGn3yHgNbLFL+oExfCRDPOmZ+DlFm7th3lQrevW72iatTEiZaC4E3NNg5vFjLtlnjHpaFRaFuSi/zUi8hZL2sN56QlUpdWc1QgQDjim2xTLYV69R+TWC8OE6iqFtlprUckZsdjgbLNiwJ3ZfLeLgAK02X6gexSh5V3l8FC9Yhc8B+GC+xN3+kzPq3AtN2irrLDgGHgEPAIeAQcAg4BBwCDoGdI+AEi51j5Eo4BBwCDgGHgENgr0NABDf/hp+mzClkTs1DvJKPE8nXoxgVgWl6bbOpO2uSKZsxaMqmWldOkHZ854Q35CPkH4QU1+w9eyqd+zbOBaQobVoLA6wCIBAhxK1FhSVnLak5Elh3JFlXO7YsogZEuv2kjHXlVCoubA/70jLWkoKypa6pKGPFC1tPqdhhLTwYl30O8hPhxVqKcA9yH2w5dc3z9JlyWEXQhnUlZMUBcZ5+1MRbowpwvtgMr4mY9p9TnpPvPANhzSdkNXUWA3JrTnk+JeFidyT6SYZYZzzM25rR7xDHiBWQ8fSdE/wIFuAP6UhZnmE+ISBfKLECHJg/1tkUa6cT1agmqNdJzZCCbLeUhzyNI1j9y7XZqtkV/qT/aI1OKQt54TObwmU/bQv1PtqXh8Rn3UH+s7bBhLExLuaZ78yP3SPMuZ1TyoLH/2fvTYPtus4zvbXPfM6dJ+BivgA4TyIlmbIkyqJGykPsttRtOx3HncSVSndVKpV/qeRPVyo/8iuVTudXOq5K0kmV2t2Ou7tkd2Rbas2mBkoUKc6gwAuAAIjpzvfcM++8z7nnBTcOLwSCpCQMa7MW9zl7r73Wt9619gHwvuv7vgUVe9gsDvB5SWdEJjyc8Jb5igrkLZ4OeKvwjkDMs17AEa8ASHbeM647NFTa+PxkqrBCunT5YNzU4/3BY+PyoR3/EiySb7bqYSNfCAtJLnxCNyHNGQN2M1ZKSZgVRMTfqeTV35RY8YREisr5V+cOaOC/L7EixZviGt4T2a792e/e23lPd9qVj4C0oMK65/gPVX5HtkhESOfk6bArn++9pvBQP1Buioqu817w7gyLK8wHc0pekS2JMjWFdioqkfeWBI+vqJ17JF48qOu75U3S0vd8vtBtCZMz05X2ogSOY/KoGJf3Be/3JSX73q3wUKdkA+uAtnkvyjnNxMyh3tfGZntf3FrNI5hkxVhIfH7Hqpq/tVs4LJQFop3WA78dzA3h5uIREYgIRAQiAhGBiEBEICIQEXjXCETB4l1DGBuICEQEIgIRgYjALxYBEdscxMtnJ7VDyyBc7BIFS2mF2tFcmH5iJIw9+Hqo3uMk0ZDQ9hagDe/shth24uss4emBcQ/iFqKRHdPeiU9bkHcQ75B8ELOQmBCsnOnPooHP9qLAJq7RrkM++Uy/FhZsZ/Y8LEJwz6S624eI5rPDIlmcGBY6+O5CO9TPhrPi70rsnsdOCP0FFch+SGwT3Qf0mfbZXQ8OeE80JFrkQu2OJCz8N41w8S/qobWka9oFn/SFA+pAiDrhNUm4weTPVCCy3+1hHJgTh7qCdGR3O/PFnDJuRCWuQbqCGeMidI89QX6Z3hVgwBrDI2JDAxot6H/9xajzpL6MF9KVjW66JPCX5Xlx7J++2tr1d/YWx8dqycxMKcn//oFidbWdjpyo91jXDsFkjwsLdswZ88d9roGHk1Uzt04SDTnOdc89OCLwEA6IzzxLjgvWCdiCI88iPDw2GAtCBu8P/f0s7wrWHWsEscWiX78HCPSF93f+1dyR3qN9L4Q3w4yBFR4JPvgteCOnBNJvvLLrcRH/dyixdJBoIev6mqISaWdqv72PjJ21wZjo215Vb+/p7WfBEWGHNeejIaFgpFDpHJXIkIxMbb2vUG6fUS6Nb517de5xeUV8St4PO1nL7w9eD+eURPvMpZPT3fG59a6e/4BCQ21I+JCAEaYkfpyQ1wTvH0LE7nyht1eJvvuClQSNTfVdw7tCdQCG94S1wLrb5H2tLyevCUtEsytyfug+eW4QjE6ofEPlVvSyYM4Qda72u8SaACvWXzwiAhGBiEBEICIQEYgIRAQiAu8agZ3+wf+uG40NRAQiAhGBiEBEICLwc0UAQu0PVLzTF8IIEhRy+kIoTSyH+T86GkrzK6G0vyDiHCIdEQHiEyLUOSMg5yDYsnknhkkn+GH+vkAfEJSQsRCO7HiG+KVPdpfTDjv3IVkhYu2RYW+LLCC0w3P2VOA7BTssFtCPQ1QNCyu05b/DZO9lhQeIXoseWTGDZ+19YNtM7rtelhilH2OEPU4WDlHLrmLnurB3Cv3yDGQsnhRHwsh9rbDw33X6ni5pHx+Hm2IesR8xhITe7MB/SILUm8kDsqhd32fG4FBXFiIcBgrSnDFjP30yX4sqYO5k0YgyjAX7ftkHROmZrPq0oRFtybK1Tti6oDTy7V5fSDh5rtH70T851nx+qZW2dLsn8WL0t/cWyzkx0YNBMFbWMvXBmTHymfeDOUXAsfcF5D/h1sgzwlwxp6x9vAZY/7TDGn5aBSHvsyq8a7yX4Mr511V+TYW2eEd5Vyz62etoYNrlE9d5R+31saDPF5mxgiwememtj+/q3dNYT36swEXP6B7zi5cVYxvejET4p7ISSt+jMEhKMl1UsKPt5NHvQKzAQHBwEvLh3wpwu9bheUDMQew5Pnhgt8Iv1SqjzUQ5JtarE1tbElr2Eq6pOt74d8q90S3VWl+UFwSeKcOH3r3koPJxPLK5VLt7a63ygbULo/c21ion5epEfoVXJEicE35gxDvJ3DH3x1R+pHv/Vucf69xWHQu3iFD/XoUcL8sKv3W8uZVsahXt9D7QLqIm6+hWPFhf/B4QCnCngzX9XoistyJ2cUwRgYhARCAiEBGICEQEIgLvAIHoYfEOQIuPRAQiAhGBiEBE4JeMADuKISe9axwCsSYq7Xyo7JkIEx/aF3b9HkLFesiPEHYF8tTeCybn+W5yziGAIBPtiWBS36GiIOQ5Dqs4VJBD3dA/RK1D7NAu5Cxkvq85NwRt0DbtQZBTII0JucTOdnYs065Je4sqEMUWDHh2WIRwu9n2PVaumVzNem7QtwlI5+Iw6ej69OOd9xaIGIt3mTvcksMM0ZdFCJ7jmT1h/z96Oax970LYOP6CZuKQrK8IBeaQsdAnpCeCD3NBAlvI3Hd7OKwQtkEQMyeMC3IRzNkVDQGNDQ5xZTz6oaB+SYm2s+PGLuas3neN0ae8ijKChLpyWZxthtPtNDR1rapcFXmVrf/jRHtZ4aJe+MODxYmVdlquKceDyHnmN+vVwNyADxjYg8ieQ06WzVpnjvhuMQDRh3UNjtT/PRVEDghrxA3WBQUyHJypy/M8h+CBWAT2POskxcPhoJgvBBTs+lR//EmYVeinkC+nIVcIx2tT6aTECgj0Lw3apW3eddplPSE8NUTYFyRUrCuHw2xzoxwUGkmX3/Xhd4QpcRg3sESMu9YBjn+rwnpk3T3KAwpbFZJ8745iuRNIiN2sF0/tOnKpPn1g+QOHHn795PKZiQ0l5n70/E9nP1BfrW2LLX3RZVtz5LuShJeXX5+8pITbk8pbcd/KmYmndh29+OzkntVFtQ8eeFcwD0/quXlh8rS8Mr5WqrbG5GXhHDbgh22EbHtN5RGVWmVc0bNaCe/l36g8MTRI5or8KDmFhUpuwbBQLBrm7cdXmVyLw6zXeEQEIgIRgYhARCAiEBGICEQE3jUCUbB41xDGBiICEYGIQEQgIvCLQ0C77z+q3j6iAvlmEaItKrYQiiN3hr3/WTWMPlRUsuezoTizvXs8SRy2JetR4B34iAP8fcAkvEl0BgXBCwlpEYNrTijM8yb5IUsJiUI9Ev9Cujv0UvacDb/0quo4fwaELwfEn5NDQxxaNIFAxA7njEAEwF6LD8NeHHx3yCnatdeGvTJcH0IZG/gOCct4wMoeKAOz+n3ZC4RrTlTOeMCD+uCIuGNhxkIAhPhIyNeSsO8fboZzf/7D0OtuyqJHhFBNPVsIgvhFsGD3N8TzeyFYMJfg6NwajBNhCUIcDCFZne/AhD5kO+PIeqsYh1/G2cLaWRn/cH/R6kNVVo8rsXKjl77cUw5qFQjpfnJxhYa68Ffn2p1WL00VDuqBaj6ZViypnLJvM4fOyWLBDxzs6QNOCAyICnguQEwjREBy0zV9QFqzTvFOwXMC/Aj7BLasY+YNbwrmn3BSiBh4EbDTn/bZ4U97XLuahwVt8twRFZI6bws1WlmFolSZfHitPJLeUx0PtSSXnNSonuu0CovK33CXJCbsf1i5GkY67Xxj+fTksyL59+scmptearR43QeeBqydrCjhsGJ9EwflWg2TfLy/DuXRwM782cp4o1EsdRvKMXF+YvdaIq+KpfJoszO1d3VPvtSdV73Z6QMrjUKpO11frW61W4VqqdoOeIy0t0qh21EeDrxGVORB0jj70nxBosXc+K6NT+v7fokTxzV7S2rnL8FU36eVG+MZCRZ1hZz6PWE1li/2puS9gcfYd1QWVBBOj6oo0UeS21ob7TQ20umQ9OZ2cE1BTCXzDEnVb0VPA3vWkbOF32fWdvZgzdsT71rzH+9HBCICEYGIQEQgIhARiAhEBK6JQBQsrglRrBARiAhEBCICEYEbAwGJFYgUxMiHRIUkhdgcFxlXDfliJ+z+/V1h/P1LoXb/aihO9cRykgwVwjy7C9pkPcS0DwgpyDoIV7wxIGchcSHvh0OgeJe6d5JDwiKMQLY7jJN3K9M+/SE4cN+kJkQt/bALHSIXkp6dzNgKwQ4BBjkMOYodFjQglxk3fWKb823QT5Zgt0hCP9jpcFN4cODJQbsU59jAbuf2yIaDsv2cLXpkRZfsdUQAxui+ac/4sVN/V5j86Gj40A9+FE78Tw+EJW3Ubp5vDTJ8YB9EJ+PELkIOvdsEtvaWgZhnfBDZxotr2AvW2TBCfEes6BPRN4B3Bfg6KXY/HA0LqO82ov9VlCFkbzncq4EuCkCwJoE5IkzlYjMd+/5Sd1MeFhvKZTFyeCTXUPJtHmcNGQeHhQIbMOI+eNAnc8Fa411DCGGOEHUQK3ivIO/pk3n7CxWECPqnTdYxwh3rmO/gary95nTpzUO78i9/0S595o4wVL/bvyir8K5Qxol+/gqFhKqWa6Hd7RQmVt4YPSDiPVVuisfHZjfnk1yv01ivrCmkUli/OLp25vn5vLwLKi3lrbjeEFC5/PZS74sBIVnR/xBgskc2BBL4XevfFc+qDoJF35tI7X9pbG6jsfvO823Z/hPZd0Grrlebqu8rVtoTyj8hL7E+bsVCsTM5vnttVddf19im5IlxRuLFoxsXR4t67hmNuSdx4k7ZOsdY281CV7j8SLjcK3HiK3vuOn9Gz36afBa9btKVePPZXK63d/XcWPHUT/aemNy7+sLMgeVnFHrqKxIweI8XVdbVXl51S6//5OhkeWRFXi6bT3aa9fenvbdEhoLEdx6T4d+QIdhujq+PHLicOqX39Kk1ViCefcNiBYPh3eTdyP6ZcnMMMloZEYgIRAQiAhGBiEBEICJwQyJwrX9Y3JBGR6MiAhGBiEBEICJwuyEgsQKiCLECUtShg+oiEcUqJbtC7e6zYfLXuqF2z0gozq0qvgoiALu07S1gbwwLDhDqEKrsmIUUtEABQesY+lmY/Txnk/sQsewWh+hllzG70tl1jvhBm/aAQJzgsFiCcEBoFUKuPK4C+QvxS8GLAhtoDwKMa9iJfRDFjB3SmTYsalhEcH/Z7/QLmQqZSO6Akxm7IIUho2lrQcVjtK0mHoe9RLjPkRVJsh4f3HPSb4edGgu58r1h5H0jYf9/2QnVvXvD2T87HdoXc6G7vo2Pckjr/7RzVPMNBucT9m2/gwOxId1mqJ08mzlDiGC+ESXA3Pkc3AN1+wmjbxCxIovzZS8a5aMIJN+mDCacE6IZa66fg0PRoipKtF1U3UTJLJYfnEhyqk/YKEDpk+AqzLdzurC+WB+sO8QH1qFDNyEUghkYIog4nJHFMNY97yVCBeuVdrh3QgXxySIIuS6yHk0e3+UzIYUGdrEu++HGdGG0VFXyBLXYbiSnWvXkR/XVUnFrdfKRbjd5UGGeKgqHVFXYpJXN5Vpp/fxoe2SmjldBXgR8qrwOXUInycPgtM7Yc7UDbBhnRd4GoVRrKyF1O69QUhd7vaTVaf7MfzZc898UanNO4sl9suOA7JioTTR+d2R6c1aeFafUT7k80rogseBikk/3qQ5iCB4YCERjmug5eUE8MzJd39xTOH+m28qn83edPyahoqDnz0mgWHrl20dPa+z71PZjaSfXW7802k0upY+snB3/DeXD+J/33X92Ue3eLzwnKiPN++WRUh2ZqjfPvrT74Nr5sfzx7x86oWTcyYNPvHhC188K19bL3z46Xl+u7WtuVu+vjOUmK2PTz66+sSiPlsYDGQUIEZQ5v7xGfwbGN/Otq43Pv7s389ii7RGBiEBEICIQEYgIRAQiAjcQAtf8x8UNZGs0JSIQEYgIRAQiArclAiKvIVYfUvlVFYhRxIj9IiS3d8eX99XD1KdGQvXO+ZCrnA6FSepwENpmQcVhj7hmEt5eF5CoELSQg3g5IEDQfpaEMlEF4e38EtTj7xHsrIXcZTc6QgUkL4KCn8mGvXGb3P+YCqGtaAPhAgLZYgrXsBkikM+QlhDRXMNuxsUOeNrmusdiYcH9OJQJbVtc8N99IJ2xGWIZu2mHQtycbFgsfX0LEemx+Uw/2T6xy+IHfTtRd1Vb5WfkBfNsWPlmJ+z5j6th45lSWP1eITTf0O5yhRJK+smVCfuFiPL/qYDtOzokOkizSBkfc2aM+A4GjBFyuqV6OyUSfkd9/hwe2vYi2vbIuexhMQC43uyFJ0tJWGuK0FZYKNaex7sp0WJG13KKDLV0vpFOFHJhrNPtN0Gb1GXt8pnxO2cBAh+FdhAMwAqRB7x4L7jO2kGMQKBATGO+LLIt6PMbudB7WR0pN3gOu1m/CEQIbiRzRjTzbvSdPHq49qTKf6vSH3R5NA1FrczqRPpkZSyfnH1pZnRzeWpceR9q0qb2K1+DllavKVFgv/IxtBprZf2vuK7QSUu6hvDQbTcKJ9PuFYIFtu/RMiGHxEWVvveHPBMC3hUi9FMlwV5RuKZFhV8qbK2V5bnwtvLBE+4NkYcwUghA44S0kgjQHZ3dzJcq7Uur58dqsnNUCbU31FdDCbVLxXL7QY0VvB9UYV74jWFuEEZXZec+iRljI5P1dYkSzNe0wkTVZW9JIaQm5+88/9LWSlUDVyqTNFF28fAxjaws4eHwmZd2L8wpJ0Z5pLknV+gdpT+JMOnk3rX8gYfOhJPP7Lur3aj8TquX9L7/rx75N8LrfLeTn1PbzKtsIXxVWhKoClGVPJARBJkh1kX/N0CeMjfyu9RfTm/3kFeFq/o3/Lu6sFNIKNa487q83eZjvYhARCAiEBGICEQEIgIRgYjAVRGIgkVcHBGBiEBEICIQEbjxEWC3NWICxCcE4HbC4FREeHGiGUbuGwmzv74rlOZeD8U9dcWNMYHmxMIQ5tnwLfz5D0kPuXZYBWaKneNOgs05S/KbVLXwAYEIuY+gAOn/gsrDgwKaTk4NKZvNG2Fin7YhywklQsF7BLIUEYK4/RBg1EV4cT4FCGP6XxzUAwePCRLabWc/U9/922uE9v43FcLS0CZ9OCQQ98DFycIZY2A/6AAAIABJREFUt8WHLMGc9eDwjnjGvZNgYo8Uni8TkkZm58PM5y6E1tmFUN49Gap3KdPwD4ph+Vtr2kZ/UHVoE3HqlMSq78vLAjvf0TEQLZh/z4VDWzFWMLvRw9dgo0WrPgbksAAgJduu7SmHg8UkvDhgVFlLCyoOz/OGBjcq0WL8dCNNm92+0MC6pU3WGt+zyd0P0bwK7w15KDzPtAd5flGFNYd4eDEfuhfkx0J7f6cb8udEjh/X9yP50LtQSppnOmlRHk79JaEAQv2wSvQLmY+dJoGTxucns3PA0HjPr0w4wUBmemFiT7onpOWV+upobWO5pmBNYVweBk5AvR+hYXS6XqqvVmYlViTVsUZdiaW/WSk2EVeKQ6GhTqi+CPxukDBRLRS7HeW9GFdopX7OjG6r0O408+cK5e5SY6N0X7HWVr4Ija7rV6o/HdnDYaHAhErgCcH9jESTveO712vT+1cW1ddJeTS8IvFganxuo1CotNcV4mm3IAJzC5EOVUY7/D7xO8XvwgXVuyDxgmvT+aS7pvH3xcH9D56pba1V/tnp5wVRN/kVXUMcyqvuJXmH3Cvxgbnlt6kmsWIt7eZG9Wy+NrmVSPCYEU7zygUypYnaI48V5ulelb5YomtSWqqsg2WFg1Ky85TfZB9/pg9f4cstmnTbnkiEOdspJBTrlXf0lhFrrlzW8VtEICIQEYgIRAQiAhGBiMAvGoEoWPyiEY/9RQQiAhGBiEBE4DoQEGENgXmnComY+XMbYeGYCLQHQr4kz4pPdMPUJw+EkrwsinsrIV+BPKIOz3Cwu96kur0AIO44IGH7Mf9VEAosVDh5NHVM2puMMqHLc4TCcagqyEnad/Fz9kLwqE3U0if37lOBBKZPyESIQIdToi7ELX2wG5w2CQlFWBvqQTZDXJL3wc9YNKC/rCcEbQ12S/djsUPiI1YgXCyqgC1eDZCiFif896QsEWfsaD/rWWFhIxsmyuIAY6U/7NnOcVA9vKGAPQUxq42QnygpKff9ods8E5afXNYotV2+v0P9MRW8Twg3844PRAvGJG+Lvr14VOgz5xtdrGDMFhSyBHGfUC8JXeWxuE+TpTzbfTHhG4M5/ITOFi0KGmRVFWgHjwoIaHBwjhF7wDDneEBwcI81RX0EOeYCwpz1wRy2ZpJL6+PJ2lfPp7vH6mn18WJoH9ufO/3ymd6ePVIR97fTUjUJvaQQOkqckV7ohMIrKvZQcv6XdEiscN/YDun/5qFB9DqJkkyH9cZ6/oe5YuUR5XgYRWDo1jUETaU8F4LCKrWn9q0Ux+dzIwp7RP4J8kD0lMdh/cLx2e9LjHhIAb/6HljyqKhWxrdWCoXepESDkdpYY00JrVulWqHU3ChtKaH1cmOj8lqp1zqlvBLTxWrnbLteXJFg8ZkrbHvzi98XxEQfeJY8F3LpMdlyUMJEW4m0m2O71p+UsHL/yMzmgoQVJQ9PHSrLYbnAGQxo84OD+aAOXhtOJD/H2PSd345dCudUO/IrJ7+2dGrq68pdUdUS//e6TjisZ5v10ugbr841Dr//5Ct6Zlp1J+VgkQiPRB4Y0njTU7LjiIQNfo8oP1ZB+KVPvY+JPDzCSrfT3khyuZGhFwcin3cVrxi8v/gdvZUO1iu/W4jSOx1+N9+W+82tBEwcS0QgIhARiAhEBCICEYGIwM8HgShY/Hxwja1GBCICEYGIQETgvUIAoeIPVODIIM8oijgjQm36o/vC5Mf2hamPV0J1YVWkd0PEGkms8cZg9zgkE+Qnu5wh/vFigAikDXZ58/cA7kP4OcOqPSsgqRzKKOulAJmLFwJtIopA7PKsd+FC8nLNO24tGpjId5uQgdi07XmwbRd9Z3M/QPzxnT4dDgpBhv4ddop2IS1to4USXbrs8cBnh31i5/bnVV5UYUd3PyySClhBvCEuIMY4OTO2OR+HvTeGRRzaz3p48N2HRSLaZ+wKC6Ud9IWxH4V0dzEUlveGXq8Wxh7JScRQmK92L6w+xdx1VG9BZ3bzvyvB4rIh2wJFn2u9ScQKm876Yq76hzwm+kW5KUJVYZ7mFPxnoxO68rhwaCfwQ5xCRPP6cA4P7nnNsiYQOixS2UOANcw78lMVQg/xmd32Z+Ul0a2GRnU9HSutpJO/Is+K47TRCqX7FnuH7qwkjYoCcY3Lo6KZC9rFr5BEQpuQa4SB4p2DhPc7eDXPGexz3pf+mFuNJGzK8lwh7J493Nvf624qB0NvXl4RYe3CqHSvXJjav9KuTdaL8lpIESMkEDTlEZETCX+HBIuqvAkeladD2kvz/fQLqvO+kYnGqUK1LeEsJGPz65fkhdBRHog98jTohLRTKtZa+/V5s1pqLPXaua1eL/87nofrOD8oceU5hW96SqGYlsu1Vnr0Q4uH1P+UhIJJnRFQEB4RIwjVxbvi36ZsN8wvAgjnV1T828CzzNFosdq+Z+7wpeMK8XRGXhYIUP1/62gMh078aH9v9uDSlxSW6qca70e67cKMPCkmhUV35tBSKvHiWJJUDkrgwIYDKnil+JjWS7NSKFfSQqms9lrC8LIugejJnCFW3IpeBrw7/DmUxSM7L7yblzN0X8e6iFUjAhGBiEBEICIQEYgIRAQiAjsiEAWLuDAiAhGBiEBEICJwgyIg7wqIcghrk+eIBHMi2/aJnm+H8Y+MheLMhPJWtENhFA8EyHXIUQg/Cs8TtgnCyaE8IHAhavk7gEMzQfZxeGc07VCP52hn2JMA0hVyn53OFgJozwm+qZ8NB0Xb9qzw5mR7PEAIU6jvUFK0A5FsIcO5MrCPz04YbW8He0Q4ZJW9LHzGHsg2CGJ2yXN+fDAuxkf4GM70BwsJOeeQQQ49ZbLfAgRjsoDhM3Y4F4dzI1i44XnjvajPj0q02AzVI1URw3WRobM6txXWKxdqdxRC/VWI9Sn18JjWwV8rLJTHSL+308G4HTasP24rEEqgHaaKobSrlBQXt/qkN15CzDXiAHPod4D3xmGY+Ozd+wh44MxapK7zmfCZ9vAg+jcqf6yCsHVU3hJ5vWwl8fuFXsixDjnwVPpVfe810sqSvCrWFKrojGK2ybEjRx8XpRW92EkL9M1BP1fbhc89J0ZHONvFgPsJt2WBQjgVx+a2kvpK+3l5PJTLtWahUO5MjO9a7yjvQk6JqTsKudSVSPFat5O7sPS6TEwTiQ75XSpyDkg35I3S91CQR8aFysRWQ7kjTqnOhbST1/uXjiv3xbIQ2tLzI/lO/oH2VnH3xqWR1+WJ8IhEkMEQruvU0nP7JJbwW7QsgWJE4gVeTszVsyr8lvAbxFxA/iMY+HcF4YnfNjyNwJnfHsQEzgh5zBPh06jzNeG8S8m4l06/MH9OniAIqtvvYRrmlH9j+tm/uvfVX/nCj5+XN8VEvtjZX66FAxJpxtcvjFYk6pySWIEQwto5mhnhQBBNKrlCcVWhoV7OFbfu7javmEKeY75uBq+l65q8AYb9XCRXeZA/W3i/btffqOvFM9aPCEQEIgIRgYhARCAiEBG4BgJRsIhLJCIQEYgIRAQiAjcuApCdd6h45z879NkN3Qujd4vc3p2Ekfs7omwhySCUIO8gUZ27AeIPss27+xECIALtrQAJS7JtCCdCLdEPfXCY/OdzNmg9f3egXQ4IfupBgHr3rUUEiwXUy4Zm4nmLIVxnjNgH4YWt7LJ2kmIIQO5DThIGyjZB6GIDxCIiR9arYrg/Cw2c6duiDM/RnnMF9OPgq3A28QYj6TBCEKcWJrK7qB0Cy8/Tv8fu+rbJXiSEkBGpnnsxFKaOhOLkgdA4cVJixXyY+/xEmG1Nhtf+h92hdU673NOWev2MRIuvSrTw3NDe7XKA9QkVQjP1QzblhCITB8j1XnhN2bU7CtdDngHmK+udwM571jTriDXK3FN43MIXuQp+osL6xyMDzwbWHFgTBsrJ3pnfEUUgaiiLw2YrFFkXDleGbX2RRKLFOYkaL1VC88xYsiY3hUKuESpFXVc0pyrrNhu+7PIcKvdBdj4R8HgnWHN9b4i2PCx6Gl2hnC6Pz3XGipW1V+Q1IAI5mVIYqHRkakv5UdJ1JZ1elxhQ7XWTY6d+su+4Em0fndi9fmZzubogb4JEIsRl0lnCRLq1Vt3qVvJjCqGUlwfGxtjcZrU82lJ/xQkJHHgDKW9Fbq63UVZS82RV7V4Zqipr9dU/X1AgqMbFE9N3KYfG9w69/9RFiSv3D6o7zw5Ygw3CBWIlBRGAcFzghrcLAgTzZ68wRAye4TvLAbyWlJPig3d8+LXnfvrdwyc0/g2JEH9X1z+kGhvCZ/9LX7/zew8+8eKSxJvH9aK/vLVeSVfOjo+1tkqEguLdZC2wBnz0f/8ERU5tFZJc/m6BpYBfCrnF5GwfrAV+e1lnt6JowRzglfabGVz8kfXPO3orepfsMNx4KSIQEYgIRAQiAhGBiEBE4OeNQBQsft4Ix/YjAhGBiEBEICLwzhGAPCNuuHM71AZpgBWJZlQ86P6ZULtbnOgYRC1iBaQZBKDDOiFIQMBClFukgFDjoN52eKkQHlSB2EUEMFHn8DjU5RmHjaI+JCGEroUM7jlfg8WIrJcDbXhjfJbg5zq2OjQUNhJehPFCfmE73hCEWsFWPmMfJCZ16DfrVUF72RBUfKcdCxoIERZWnDPDooLHYrEHm5yXwrlDICQhkrNjMzmZ9SrJYuHPxoAz9iu1dvKvg7bEh1ztcEhb3dBe7ykXyUzobuTDrt97I5z9583QFnedBMLwLEq0gMBNJVzcioQouOx0sM4QHMhH8EeuUBaqU/2/xSZzs8XwSiFJlzWhzCWEPAQ2zy0O5svJ5FlrkNomvC1GIdqxxiHNmS+epeCxgShGfZ6VZ0Wu3A4JngAcrEHIbbwFuMYazWtCv92U+tRMZx+TJ0ZNybm5N6+cF421dJx3B0GC9Xe1gzVIIntI+v5Of8QKhTgKS6/n64317iWFPXpIIs37lDy60FivnJC4UKqON5r52c1UJP1zCm80Nb1/+Xfl2ZDI22IMsULEvHJavKk9qr1d9eXqliSZVOIHYaDyhVJnTPkdxokeVqq1C/I+WJNnxTgrTmQ9797LKnhxvZ0DDBEeFLNK61ZhqkZnN/5InhZf1/cTmq3P6d6jKqxnh2RDuAQbrjE/hNziNwEvCn6jEKH4HQBH7DmmwrzxDHZ9S8LL1O47Lh7YuDjaOvvKrqMaP+8bv3cnNYZw/vjs4Se/+MHvLLz/1A/kWbF+7tW5XcLnQYkxrIOPq4B5lnzHli2lgDnWaW5OKun2rIouXXa2stcO838rvpt+r8B5p4N3k3f0dhRUrwJJvBwRiAhEBCICEYGIQEQgIvBuEIiCxbtBLz4bEYgIRAQiAhGBnxMCIqch4wgHBQG7nech1edUokJxNAlzX7gjjH1gVkm2V6C+B/WyYZkgzyxccN+JUf1nP6QohOtHVSBmIQezng8m+WHmIAlpw7kenFPCxD22OgTUcOinbNgkk3lu2+IFzyIGbHuQbIsQEJ14g0AWIx5gK9eo41wXg1Atfbv4bOGDNixcZAUDzxbXsNn3hgUGCG6T0eDv/sz2ZnF1P1zjvhMC01fWM8VYYRtlQeUjKkq4PfZ8yE/Nhval0VCY7oXeejmMvr8Qxl54PVz4ymsayb0qnx6MCQ8UhxbyeG7lM1hBIBMqqH+wqZ1wUCTeXu2kl9a7YXSr1/dEgsQm5BfCjnOdsLYIIcQa5z5zC37OkwAJy856CFfWOWuPuaQw9xDokN2sL4Qz1hgkOuXxwXXmBLIbgW2/km7/ZjfNf0uhoSD3F4pJZ/lAcupcM5RTCRasX2zo7ZBwW5f7/bDOOa4IwcO4Ny7multr8uFIw6g8BEZy+VCXUHFcAsOd8rCY1nm5k8vvKVY69yoEUmnl7ERja61SWzs/JtEjuxz7AkQQmb+qUEgFiRwkqd7KFSoHi6WunAjSkC90t5obZf3m9PvjABNwfbsH9fsJvnkdG+vlF9XepMJLHaqMNb8h4eKTusE88P46wTm48pnnwBSvGkQm5gzhhza5xu8C9cATEZI6vNN8PqMwWcmhR07h2VFaOjn1tAScdY0P8WlKIs5nNpdqDz7/lbvx0GBk5CfBcwRPgT9VYb3we+ScP7zjfJ4XMO1U8bl6XZyfLmsTCFDMlX8L9PGWOsCYwV4tlw7vJu8o8xWPiEBEICIQEYgIRAQiAhGBiMC7RiAKFu8awthARCAiEBGICEQE3lsEJFbALH5K5TEViDBIUv7MfkFZdyfDrt8uhulPjYd8VUm2i9uJnLcJPYjOQ4O6TjzsxNUQoXw2CQeR653jEG32PICYynoNcA/C1qFbGKzrZL0ZLD7Yo8HfDY5DJnnnstvI9kVdE//Yg60ILQ5pxdl5A5wUnDNEM9chnSGceYaxWoDBdj5nhQa+2xaPg+8U6oEr2NMewonzaViY8RZrRyeiP4cayiYKH+7DIbMQNr6g8lwoz50MnX2K+dOsqpRDYbwZirtHwtxvz4fO+XJYVZj/fD/PBvP1Jyq3k2DBnEM0X0EGFwey2LF6+ImSMnQ1u4gRkM6Q38wXa8ckMmKFw/zgRUR+Eu5RzyQ87xfCA+sCUp55Q6ygf3bvQ0rTdkteE9ShPa8v5t7rfVGf75GXxYSEi4vyrsh1Q27vcjp1Ry2pk68BIbFft/LnK2EH0YI26Yf3GDsdwkwfZchmMvP6c9U3xneH/dWJ1hvyhpBo0ZtO8umKvCdmGxvlWYVdQoxIV8+OF87/dLYpgv7HykPxcQSeNzn2fnOvyjPjaNqr1JXvYUz1KpvtfFB+h1AsdyQwVBRaSpk4rvQZ4D1AuMkKFxZ6TOz3G88efZGpWdivsFD1bjc3PrVvdUJ2P6864A+23xjgwrgRH2h/t4qFQ+aHdcDh/DsIC4T0AlM+039flJJw05WHyEnlsxhRTo+9bxybOytcHpJoc8cgqTaeGQgVzl3DHDOPvGO+dqUAoYzcymHRS/JKWn75J7BvD2uN3x9+sxjLreZlwXj4bf2myn81mIPsCZycM2aH2/FSRCAiEBGICEQEIgIRgYhAROD6EIiCxfXhFWtHBCICEYGIQETg546AQv70JFpA1kGifV8FYk3bnEVbT35gd6jcNansu0q2PSEiKZVIkbDjGNKMXa7eDQ55BnFO4c97yDjIQQ4IJuduyIY+MQmfJeq45p3eWbHBBG3Wa4K2h9sYJvizHheum/V0cLvYanLfhHDWDp5xQmtIypMqjJnrP1Y5ocLOeUhsyDSLFtzPJoelP3s/eNycIbN5xjk3IJEtejBOPnvLup83gW3cB3C/pS71IEUZF2G/dofS/GsSK36scFAfCOnWNvFbPXx/mP2t9bD87DEhgcDBOCa1Ni5qjdwuB1hCLv+tyiP9QQ9mTIsjreYk7+STS/kkvdjDA2mb6Hd+E4d/4t2ASPZcI0axXiC6eQ8QgJgTdogTVoh6ELS0A3GO1wbkOuIB4YV4N/EAYP75zLojoTRtIXLQ7pSEjYqEi7VWWiqsJuMH19NR2kCE6K+lrFjxw2//P7q0fSifBWPGvu+p4Dly+UiSfGPp1Px9rz5ZmhiZahV2Hb0wJW+KcnVi67S8IhQOqlhbOj3ZU06GXKdR3JJIcEGhju4u1loKB5WEbqsg74DLIsSoPishdm7usijR00KTJ4a8LvoeGENiBXbwztpby3ZdLRlz1nR9Tsbw9uidmH5hbmGpO7twCYzxanB4J+cNcdg15sMeFAgXzskDjnizUMht87QKggUHQm0/P0mu0KsrGfmahJEHVXZtLo2Ul89MFCRcjGlcC6rD+0S4KfDGe4C+sIXyln8jyaOi2WnUi91WQ+G5rki4vaj6/E7fimIFmPp3zr+hw54kvJu8ozHp9mARxlNEICIQEYgIRAQiAhGBiMC7QyAKFu8Ov/h0RCAiEBGICEQE3nMEREhDskPaQaQSNgixYjTkSo2w+x/MiMiW9HBAoYRKY7pD2CjqOVyTE2LzHaKJdiD/TdYOCwzYnyXt/d3jGibluW6CHkEFEguiargNixFZfNy3RYkrY9S8uUt9uJ6/W9jgeYeNAqunVCA0IXjZIX1BxTvT2f1t4cHiDTbZM8LjsceHQ1r570gOOwWZaQHFz1t8cRseK7hk84dkvU48FufeoF2FghothuqRg2Hr2MmQlI+Exut1ec+UQ+VwPhQK64rnUxLCe1Ug1NlVfrscMMMQ13g09A+HhMoL/T3l8JFCLvxAlyGc7XkC4eycLWf1GeECIhvRh/XBAVmO6AD57t31EO98R1Tgea8h1hhriHeKNrDnNZUPqLBeECgscNEXYgNr46JEi+eV92JvJy1uKq+Fn79WrH+LNF9VGx9WwUOkHwMrly9+ottOZlfPjbR6veKR8mizO7lntaSE0a1CsXNJORnmz7wwvynBoSTBgbHcr5wOven9K3q2FxSO6bRCM+W77UJeybRfVJ0J4Wkvpn43unZJ+S3scbWN1ptHNscNuIEjgg5Y/MyjL370ko68QFae/+pdr9z7iWM/npxf21Ostj+nH7g5YfWiPCOeGYwXjwWEWOaoH0JLBZwpiEgWoLCH3zxswGYECH7vttTWw/IWuXdifn2iNtG4uLlc+/b6xZGKvEoOKi8Hc8Ec0R5rg3whCCB3qVjMzY6nzsJT7orydiioYc7+cmJ3/w5eC46b7T7vwhNXMZp3k3fiChXnZhtgtDciEBGICEQEIgIRgYhARODGQSAKFjfOXERLIgIRgYhARCAiYAQg3iBWIey0HVokaZq0wszjhTDx4fFQRqwYL4gzgyQ1oe5d/RCIkHDsBIc8c4gl2s56BbivrGiQ9X5wfSff3inPA6QhO8wtQGSfob4TWGfFgCzT588eg8MqDbOBJgFdj35on/GzSxoPlCdVnlOBwCSJOAIGpDIEpp93mCjI5+xYs2KL2UjqOJmuQ8RAVlsE8lg58zxtQ3RC4hJbn532zAVkMCQ29mSFnaygo7mUl0y+2pP3TCW0z6uNcyJUcyUJFe0w89kDYenLtdDrPaueSPD8bRVI9dvhAG8IagsNl9WySi4kI/mkUe+m5wUsaw18WRMWN5gD1qhDpoGXBTx25lOP+oSCon3Wsr1o6NfJt3mH8NaBFKewzu5UYW055wprxR5MiCSIJosi4SUTJErWnWd9eN35fdkxdJC8LXryskD0oD7eBNuChY4e+RM6rSOdRmgoqfSUck8siYh/rVRpN9RYffn1yV0SBPbImyKPviGRIh2f22jtvuPCmsj7rkIibSjp9KZyO6Rbq5VXV8+NH5eIcFoc/EEJFQg2ziXjLq92di4W1jf4vq1DfZCLJ1GIqvlX//bwsfm7z3cm51dfHJvbIIn4Ea3vLeXOaCtBt9tjDnifeK/AnjnFTkRJvJMcsg3Rwr+bPIsI0Q/5pfYKudGesnKETQkVRSUWf4l8HrKF95MwXST//jUV/14O//5shxlL041up70L4aIfXuvNESOWsX6yIujbwuMmqcRvFXjb023YbMbOO+pk9DfJsKKZEYGIQEQgIhARiAhEBCICNyoCUbC4UWcm2hURiAhEBCICtyUC8q6A/LtfBfKTnfR3ixnbF8qz9bDrCwoHta8WctWitktDHkHkQcBCKEFuEpbmhyqQd+wWhtjjM4TSsFhhYt6hoiwqmKwzH+ewS3gqOPk1RCB2QsRbRHB7EIpcgzzMigJOqM28mliG7HS+Affjs8MrZUUNnnVYKtqDNKYtRIsPZvp02CfvlreHgzFw4m7n1ciGdKIPvpMPBOwgtamPCASekKaMG7ss9kBoQoxjhxOAQ/AhcBCmC7LVXi4WgOjHniLbJHmSKCdJSUm366+F2sL+oFMoCPKxh3aH9adOhcZ55nhB5YjWyTOEDqORW/xw3pVDHqcnTckkwlg+bMwWw5KAZI4g28HdB3PnOWEOwJs1wVw4TBrrh7XsHfzMObvJuc893iPWPnNJHwgdeFywPsjlAEnN+0XdF1RIQMwz1O3n3lBYKN4b1ocFL+zrkcPCh8JDXf48+ODwOogpl48kp9EnyYiEi5GekGmsVaf7ibFpP5FA0k2KIuL5TXjzmSRdr01uLUq8aChkVHHu8KWVfKl7TqR9qpwSFxQ26osbS7Xq2rmxWYWI+s/14BVhqIYNG/rOu+ADTyfEw+GQUcNN/KZs/HB9pfrTE0/vf2llfvyk8k0sj8+t39Pt5N9Q/oxjtYmtp5R74ru1qToeZqx7xCTahRQn/NAJFX4nwZ5wTL816IR5ZL6YQ/++LMvbolwst7dmDi6f2bhUqwuHSWGFEPQJFch25ps5G/b6oll5q6Sh02qcbzfqR4YSbnOfNcocNCU27ShCDQNwo39/+hQQXnHw7rB+dzp4NxGKo4fFjT6x0b6IQEQgIhARiAhEBCICNwkCUbC4SSYqmhkRiAhEBCICtw0CEP2HVSDcDok6nxIRuRImP1YIIw/sU5igXkgLIrYTiHNIU8hTyCSIVr5z/WEVduCzy9u7vs3zDocnsucEAGfFgazXAZ8h4p0fgzYsQFiU8AQ5OXfWg8DtQvrzdw++ZwlChBfIRe9AHyYN+8FkBh04lJKveTwwvu9XgXzGVg5YN0pWWLEnhMfrdj1e+uZ5E+BZkhlBCJaZZyBKHSbKnhXssuezRSJIPMhjbKB9x/rPeoyYmObaaMjnRkP1DiUSeLkj4UJ9K8Mvm/QL41oP55lPSGGEGmL/Z8n5wZBvuZO9Ui6vCXa3tzUDl4T+aifcO5IPX9Ilh2ViXiC1mQc8IJhv5gkRgblgfbB2WHMcCBkmwnkOQYJ3kDmmDhizE//fqeDdggjCNXbVYxPrAcKbuTVx7TBR1MVTgpwqLw36415WKBtcfssJG7GH/AzbRz8kUTd02w3loeiwxmpEJ0q7OSekvuLv9VSXp8KaxIlmodidU+il0VKttS7yfkv5LiCZL07uXR2RN0Yib4u1l75xZ0E5Hr61sra4AAAgAElEQVRK8u3BmNyeQ2Q5tNpONoMxouHbOfhN2i3RoiaxZHTl9ORp2bRr+dQkQkmp10teKddaqwcfPn1vsdqqFMrdhu5jA3PInPKbhweZvWEQBW0r2PZDQqmwBrjHe3tSobFqR3/1tYuvfOvot9cvjDHn/Mbye8IasMfIsHdFfzxac+VCqdLLF4uLnWZ9YTssVP+wcOWk7G9n/DdjHXDFo2Wnw+s55rC4GWc22hwRiAhEBCICEYGIQETgBkQgChY34KREkyICEYGIQETg9kRAu+Y5IFXZpQ1xyp/TEyE/MhWmHt8K5YNVMZZrojtbYtAg1akDcQmBx45jyPVHVYjDzgFx593WZtgcjob7FhXsYZAF3mS860PK0hcELAQffUIgWkAwoQxJb8Eg257DKtmTwzvYsRk7hv9OkvX0gAizJwf9OKa9xRjuQ0DaZoeicogbCyROAO6+dho317Dfnh60ZQwhu18e9MM12of0tOgBSWpxh/t4j0B2I0B5Fz/t2w76cSgj7ieaVwXyKc6Fwu5LodrbChvP5zX/JSXlVr1XGTekLvNAzPjbQbCwVwwCDaG+tt1S9D/O3ZC+UVQYoVyiNZH28QBb8GaNQlQj8rA2jDuPcY+5Yq0yd/bScX4GhAruE/qJuswzuRQgzREEaYM+IP3xKMI2+iB8E/eYJ657DWCXPY92ejd0+y0HdjHP2P3XKp+lBoJFp9UMIs1rhWJZnhJl3gF7NNA3fXr9KuVFF4+KVELFlMQLRD3/VkC0vywhYDzJpw/LA+O5Bz770uK5V2f/z59+b+GvJCQ8pvu/PWjvuzp/XuVq/25AWHGorZ3Gkr1mTxN+T8C5olwa/6nOXQkYo5XxxoGJmc1NJcuelEfI3NqFsa3qWOM71YnGkmxlzTMH2IJo598c3kHn7qEvvnPPuWSYn7/Qm9UulJRlfKv0qkSRBV0Du6xnwI5iBbDzn0SisW67tUCUtkw2crDmN5F58m/atTC42e5vv2rb63yng+tZ4ftmG1+0NyIQEYgIRAQiAhGBiEBE4AZDYCe35xvMxGhORCAiEBGICEQEbhsE+HP5V1UcE165K0TEleZqoTi7T3krRI5VSiFX4D4hUhAM8B6ADCUcjcPQQJxBIJpoYud/NtFvVrwA3Kw4YBIfWyBNIf0gJInL7/jxtA1BCCGP4GBRw+1wHxuyO8mzf+fwLnMIQ8awU4Jf28gZ203gQiR7FzW2Z5NXmzB03w79Qz33zy7xbNiW7Nipx3ioAwnsHd2Q3hCbFIhc2u/vcB/Ud1gtPClMVNMWuFOPtuxZwnXGAnYm+bCH75C55CZph6I25xcmR0K+kg/dRiWUdhH7H7IZrNi5z/zfDgdYQVQTfunyUdKsVYVeJw0/fUA+FbVcX8MAF+YPMp4zQgFz6dwGrCM8I5z/g3nlmmJv9dcEa50QTIhSJGHmGnUhwHkvOf9A5bgKc8+zzPe/VvnR4HmuMd/YTUHsIBcNQhPvKt/9Xujjzgd5LHQHQp92/0Slnx9ASZ/7pdPYEmfec5JwN2JvK6+rhsIgLckZ4IIIeoQWDt6XXxnYQ5us/zGJGR8tjzQ/f+DBMw/c9dhPV/KFHmPFQ4FxIqD+rPBj4P52/02BBwzeJrSHtwQeEOBzUDY2KyPN3tjsxp2tevGDZ1/affjC8Zk7l16furfXTdqaDdbAt1WYJ/fHGJgDwkQtqrBWOJjnV1QQDBnzQxJGgtrb2Fyp8u5gB78PrIGdkmwPmumLP1vCerNZXz/Y3tqQd8sVjgSsNfolfF/2N9bP3+xn1gc4sbZ4L3Y6mBdwvx1C1N3s8xntjwhEBCICEYGIQEQgInBTIBA9LG6KaYpGRgQiAhGBiMBtggDkGaQmpOkREXQKB6T/5v+wqB32JcV+0ZURvCsg7KgLSYQ4wA5Xe1xwHUbNpL3Jfs6QT9mQNIbVRFOWdOR5SF+ECggpiFt2aEPOs7McAtQhYhy2x+S/27H4YfLW/WXFCNvE2fX92d8hzByGCnLR4ajcT9ZjIrvT1/dtl9vxd/eDXb5mYQGi1rvx7eEBHggmCBm0Za8Jh7JCdLCwwzxQIPp4HvKZ7+6T5ylmPz3W7dBbSUGeFmNroTBWC61zuTD6QDkkf44XQUctMAcleeTsVx6Lq+16NtY3xFkhdLJrApuuEI3kWJL9nrWZeYeUJhQWXg2PcxN1oqwWlXT7Y9qav6YE3Ce1QL3TnvUJ1g7R5TBQFqOoB87ON8LZuSyYQ+cuQRBgbh0G7IQ+k9yd9hASIP7JsfBJFch3clYgVvCe8B4TzgnPDNpnPbF2HG6MYVzrYJ4RUxAMsKN/pN12aDfr8rLYyhXKb8l3DUEP1mWJDudmDi3nJufllJVP/Y7w7jA+bH1cxbkhaGhFwsXGriOXiieePrBSX6625fXAfer6ACcEAA7aspeTPQ0I1XStJNxgwW8Y9dxWohVRXDs/ttJuFSaUGLvTWCeteigq5NX7xudGTo7ObrQ0Dp6xMIBwBEaEwPsXKl9S+SMVBBQEIuaSQoLtvWrv7Knn9jblPfIZXWIuETUcVm8nbyse5fe1Le+Ki63N1TEl3aa1y2DoA2NhvsHhams4W/9m/MwYWet9L5+h4+v6zrvJOxoFi5txdqPNEYGIQEQgIhARiAhEBG5ABKJgcQNOSjQpIhARiAhEBG5bBCDaIMje10cgFTFXu6MSRu4rhuqRkZCriLQmMXM/qS7kKwUinDPhoSAXIfQg8ShvkoFvhmmCWPN1A20PCYdrMrnMmd3p7FRHKEC4gDglye3jg774DjHMjuXhwyGnssIAdbKCgZ8ZDilCHRNg/H2F8Thhsu3l2WGiMTsW3/eZcXuM7jebI8G7ibM7pbnvZyDBwRdyzmQteGIb9jMP7OrmHgQuYW9MNNO2E27z2USpQw4xpw5JRMwZEqtfCuUD+0PlQDfkJ4ohXyqEXgvBAsGkv/P7rZD/4q9IjMjO57DHCgbZC8aeKGAFrlns+5gPhI00I2CkSgAM6czOeicxn5d0p2QuYXOlnb78k42wKAED/Nwm9SDZwZjCunHYMHshMIf2RGKN+33BDp63R4d38FOHMESsBTxp6I/vvBefGzxP3Z+oUJf38csDOxga7wfvyfD6496OB14WH3jsD7EFUQoPqg9QMUXFzMt0xTgilwJRxDIHgoGI/d6Fqf0r53YduVgsjzY70oNYixyInNiJwAKpz5rjNwQvBTB7WF4Ze+786PHv/OSv7v1/u638P9A1J9bGftadhaCslw848C4g2CEYDf/G2EQwP6KCWIB3hX8belpGhU4rP7J+YbQmwSIonNXJjYsjqfJrjM3ffe6Qhunk5rSNzdhrLxl+OyHUmRsEJkQEbF1Vu6cb6+X8xcXpQ0r0fb7bzhPqin4RXa8lroBxvdtuX+w0Gw9lQkF5PKwbRCLe41vi2CHhNngj0DFf5Aly/h7ekf9bBcFi85ED47eqYHNLzGscREQgIhARiAhEBCICEYGbCYG36759M40p2hoRiAhEBCICEYGbFQHIL0i29X74k552B09+fDTU7q71vSt6TRHUqQlDSCNISAg3yDknCjYBaA8LCwEQk9TlOkKAidOdzuAHAWfPiH6SXBWIY/pcUHEy42yuC+NuoWHYUyLrQUHdLMF1tc/Uc3uQxA6nY6+HYW+N7Hh49jIhOjAu69FBu9kk3rafa86DARFLcR4L+gV7iFLjwxm7wOjjKvepICpwHdyxybv53T9tOBk396jjfBkSJZSjpDh+WMm2m2HkHgWJekPeNVV2xlMHotAksm3+uZ8hx4dKou/GyvkAEGgoYAYmrDfIZIdlor7JbbDg85jaKamwPin9v58ihIg8tQAFuf4fqRxQKQKWcleM3D2S/H2FhJoczffXK3ODVwTkO+uSOSKMDYIb9kFw0zY4Yhd28hlBYFEFcQN78CaCeEcQQuxAmFhQYe0TEgxPD4QPJ9qmb0h85pz8MX723kE9CHzmi/54xh4f+njNg7WBCPatQR/EhQq9disQnijt8hq+5ShIsGjmC92zuULvy/JKAAPWjN9VxsP4Ifa57oTR3G/qjVmf2rtSHJ2qgxuY+AA7/4ZkvS64z9gYJxiwrq+2256pY14WVJgvsGOOWRcdTfmikn7Le6QYmhuV/c3N0nS7URzdWq/cqXNeYsPfqh52MUc8i3CBAENCaN415svJ7llzRTzV5DnS3rg0UtXzjwz6w2Zsddi2K1SfN4ccemmv88rm8rl8r7Nj+pGvqi65S1YlMN2qhD2/faz5/1rFwjTvE+8i7yTvpt/VDHTxY0QgIhARiAhEBCICEYGIQETgnSEQBYt3hlt8KiIQEYgIRAQiAj8PBCD5IPGI114JxZFJEdaToSyusyDON21DJnrnsklwwkdBNLJjGkbNu/2HwyHxnAl2hyHKeirYG4Ln3A5kLmQgfUFqQgC6X/qBLKSOvQiy3g5ZccJEXtb2LH7Du/L5bhuxx3b7elZoyI5zmHS0DRY5siSqRQYLHFkbqG+hx23YdntUWGAwAd8PHaOCeASxDSnMmfvOmcCY2DHPsxaUwNA77x3Chr5prxpy1V6o3ZcTe9/uixiECNsmZwlD9JDCQl2NaM3i+159ttjicFgOCeYE5BDAkNEIN9gIoQmBDMnJ5/tVCG9ksYXnCM9EfdYvXgkIBnmJFf3QXA/vH7NnChg5ufR2zCP9T4Gzwlon3DNdTCragQ+5zrwiCnBAXNurhu88Rhv0D+FuUYp1jR2MxyQ6dR1eDYKc7xYlGEff20EHc07+BArCAu+LBQxCFTEexA3OCCDMP2OzUDZoZufTIJcF/X9D5c+p1ReNlHy73aiH7pUkOmMfeIckr1Qnti6K8H9FHgqEsbJHECGqwIV3HLy+p/KMisOl9XPT5Iu93Qcffv18qdp+GfFDhL8cfvqvDx4aYIEoMXwwJtb/z8ppYZGKZ8Eh6+1NB8zFcQ1xRYVQToqAlWstn5oal3eEQjLlnAPjNdXD6wTbF1V4x06qIKiANaIV79Zir5t7ViLImgSLhgSLR4eMZt5fVOnnCNnhuNDeqn+/XV+/D3uGDnKX/LXK9YT5uko3N+xl5ov1i2Cx08H7xHvRiR4WN+wcRsMiAhGBiEBEICIQEYgI3HQIxJBQN92URYMjAhGBiEBE4BZGAKJzVHR2rx/2p7znQph+/I6QGxfBWFJYIN3dDv8CgQRBCsFr4hOy1XklIGxNyNMmBB5/5me9EWhnmKT3fee9oI5j75/TZyepZSc1fZjk9HMWF7LCRVYUGZ667L2sLdnnsyIL/Q3b7LBCtO3nhr01suLJcL2dPDB8jboWb8DQggekKdez3hmIDZDg4O3QVQ6/BQkLOU99t4fdzmlgMhyy17v2t/vKT8i75sRSWHtyMzRXWAOMhbmG4L9b5WvDoL7b70MhnvpWDNo01s7v0dcNBvcRK7wGqY5YgxBBMmJIcL5DluPNwDqlDRPWtA92EPOsPfBjDniuNVrOtzaaXchpwtJ8qG+L7raF0KpkM50+fFRp6Y/Vw9cubgfzAkPw5j1x8miHi7LQxDxQsJm+sQ2CmzljfrGNZyDoecYhoqhD299R+bEKIZjwpECQgbhFDOH9wHbCHhHKyvPv+d7RLaJveeZQOCh/o/7xQXu0uQ/Boisvi55yKuBtkeTzG/pteD1Jcn0PIBH746tvjOeVt+HXRmc2TyxMnSIsFCID65Q5o95zKosqeIVgO+84IkZVdXO777iwUCh3nlfy6z6Ora3i6Y2Lo0+p7aPdTn5aqDwxbPN1fEd8+Xsq2dBRFome1fUl2fBbEkpq8hK5FHLpyXypq0hYPfDF2wTcPaeIE4wL3HlvGAsFEaKrNrCfuQZD5oCwXQhnTpyO2eCK0HLF0et0vtLYWNkvhUjr6C2KBWvBv4/XMfQbt+oO4aB4Fz6t8omrWM07ybt5y4TEunFnJ1oWEYgIRAQiAhGBiEBE4PZBIAoWt89cx5FGBCICEYGIwA2MgHbKcxAjnN3bkIbtMPlYOZT3NUN3LR9yUyoFhQrKQV46LIc9IAhTA4nqBLpZIQBSD1J2WKzIehZYBPAOepN+TjYMgUyBlIYA5rO9QfxsNjwSn51ToJ8getB/dre7P2ftsrcE19weuFioyAoZnk17W/DdY+Jz1vNgWAyx0ACJ6RBZ1Bn2AMEedqzTh8Mxseuefpz8m754ziGisBWCGsKU63yn2GODz/YegV6nOIQOApSFJuyRcCWFqtdSSCi40X4f2APhT72jSrr9nh2ZxNheP8bEHgHOjeL5gOjHk4Trthtc8PoBL0hhsGDnO2IM68ChzCx0gBGEMmFlCKUEiW7PDd6Dpfnxcji13Fhrdnr/Vt//UX/AmoGeitIyh6lCWG6WwtH9lfD8pXaY0GX6oX0IaLDGPghVrzXGxZicBB1wESSYB9b2fhXIbj7zToE5dnKG7KZ9yH28SNixf0QFLCDN6YP+GL8zNLu/D+oaQgeijdeAPl7zoE36Q6T8rsoXLntZbG2KS5f3Q6GQ01J5plAZkadJMiIr6ptLI4dyuXRGZVoeBotJXrGktkUZxkT/vMuQ/LznX1dBDGCeWKsQ/UdnDi7Vpvaubsgzoacy1tgsTa6cmfjT15/b+5HmRumJN9OXXHMMwxV+a4AV17GJdcE4EZs+JbHirPpPR2c3+0nDJZ6cr4w1duv6jPps6sz8YDvzimDBOmM+mCdEIoQExrmHdtTyKT3HvCFYMG7ni2Etk1Ca81sOebCMKRSUxrnj+BBWvqmycouGg2Id8C6wxnfyqAEU3kn/ObEjSPFiRCAiEBGICEQEIgIRgYhAROB6EYiCxfUiFutHBCICEYGIQETg54MA5BCEG8TZ/pAUL4WRB+8La0+3wuxviDjVNuq8wgNtE3Ts+obcpS6hOiBnIVezgoCJUyeVdax46kKoZgn6bXJ8mzCkngla5xOA3HxIBVIxS2ZnhQ6ehaAlNAtJaCGybS92QuBDTEMYOoRUNiwT17GNXfaQlvTpnfxZIcW2eqzZv8tkPTx43oIDNlEf+xmfCXefh/8+5D4YDzZDqFIguGnLZLeFGF26TIbTJlhwD5zB0GSoBRWHImJXP2Q+Y4ZctajhEFaqr1BQxbFymPpIElafYhc4mNAeZClk4rs6BiIF46VNizcWabAdchd7wI3vJt+pS/+Q3IwLEQXMIe45IwBAKEN2giF5FBwL3+Q+8w/Jz1rmzE5/5ghyHkKaddCWh0VdGZnBEpz+sTr77xl0TpZIsNjaV05+7VwrfUlZXuYUIiptp/1nEaOYL+OFTRYdnJOEa17j7L5nbA5pZW8P6vqdQYSA0Of7R1XwGnGIIvKWsF4IC4VXCWPn/q+rMG8c9vqwR4A9dga3rzyJBPeFVN4WrLsfMmyVL/hGc3NNYaHaYXR2Ty3t9T6rGEqXJHLdIXL+UrtZeF65H0Kp1lrQd8QfxsuaA3+H4kJcAqu/O2gT26jT9zJBLlPy67yKlJHQqYw3HqtNbH1nYn7t+8/85f3/rNMq/LHqgavf5R3HcpWLYMzvlufAgqVwSg6FJF0tVVtteXlM1lernZHp+ppmqCLZJZ/kL3uM8VuI2MVvCmuYNcM8gRfzebLdKPxo5ezEHnmbIBjt5Emxo1ihd6OV5HIPypOlnPa1niuOf6FvfzXAdNuv59Y7wIX3B2+Wjw1wtdDDaP+xCnPYjeGgbr3JjyOKCEQEIgIRgYhARCAi8MtEIAoWv0z0Y98RgYhARCAiEBF4EwF2CM+LFNwO3zT+aCGMPTIVRu4fCblSLiSVaugl9YEPAEQc5C4ksZP40pJZNe8HzuaBMEnuOhDATk7sJMmcHbKIeg77BIFNn7SXDY2U3bHuXezfVx3qY59FE2yDmESUgAj1jnzb4rwBfOdZ6nqXfdYTxPVNrNMu9ppEN2nKGcKcMVOXNjmcKBxiNBv6h+eze6jt3WFxBgL0p4Pxs2sf8h5PGHtb0HY2JwHPZwUACyDUs8hjm7AFMhnvFcYCqc21QW4Q5XIozBZD4401XWWneDrIYwLpPCbPnDF5WfTdL97uMUiUbc8UCz/Y5bm1hwt9EHYqm2gZwt4eCcwldRBdaAfbCY30PhXWAWNwKCzapx3nlWAuII9ZY1xDsGDOEUAQMMCEdQDGW+1uX7B4SeU1NfSFNAkPKa1CqOZCdUs9KzTU6/kkbCmvxbFON9ylW8wRRDJrCxsQzHhfvLue72BgQYNxWIjiusUZPlOXwx5GPMOO89cG7TGX7OpnbbDGIcZpz14W9lqgPuKN14Y9MAbN/8wT46FPRBDGMd0j4bYUhXyhGLrddihVRunfYY2m5FWRE9F//uwru54vjza7k3vWdikPBfgyDuaa3xzWHPYgMIKVwxxhP2MHE/C7oHVXlx5UKI+0npDXwjdGZ+rHV98YOy0xhPBk1/tvCotg9O35cSgwXUrrxXKnWx1vrBdKnYrCUO1r1kvt6lijnSukkOf2JuM9pH/Wj0NEIZIh7pzR2/K9TrMwqXBWgivH3CCmnlCxxw1ix46Hwm41lLtis6fUQTsc9LUwaO9nCk9Xa/9Guz4UDsq/fYwTryIwz4oVCKb/6wDH6/EWutGGHe2JCEQEIgIRgYhARCAiEBG4ARHwTqYb0LRoUkQgIhARiAhEBG4rBAjjMqui0E+Vehh9UIRhux26omKT3pb2ja/081psE5KQqZCgeFdwjcO78g2aPQxMSHOfAklqMtfhVExQZ0Mk2TMDEtk78E3s2+PB33metiEESUZMbHsIZ++85jp1ICch9ywy2G4IS8ZFHYhI+uSaiUD3Rx8WBty2wyrRBwSxiWl22bN7nPjqtMt3iHAIcMZtTwsLFdkz5Ljb2w7PtU2KQnZDztMGBCnXszH4aQPcLVgwBofGYqwc1LFowWfsZcwQvrRH31zfzjmSkGQ4vx56W0q4XmB9QDJDkCMkgMeRQTgxt7/jGZFCpaQC6YjQwPyCM9/tccC4WFeEpiKcE8ID3xm7hQRsfFDl/SqQ3FxnBzZt8gxrkuc5E/roByp4YnxGBTGDPsAMwnNRhd38JKdmzJDJJIEGc3sE9b1gyop4NHiO/i71F4T+B9Alne8dCZ1aLjkxWQgKF9Qn3VljTrxMW7RJgma8H/DgwDYLWLxDeEhgN/0xh+BMN9RD/AIn+uY+ggH24hEF4Q0OjBNRi3HznXnnO+OBIGf9YZfFOgtxunTtYxByiDFwXCaOES3arS1FDdO0XBm3iLVRIhTS0qmpkVe+fTTf2CjjRQL5jPDhd5e194gK6wGbvNadgJxxcDh8FPY/pDBTn6qObykR/FVDBV1rUM4dgoBDH+DK+8vB3K0UK+3TlbHmqkSL0uhU/ajElhlya6iwjpj6RRV2+HMwDtYRQot/a+b0At3X3CyfPPfq3Bu6irjBe8N6RhzZ+d9BaarwUb2X5VmxUl+5mOv13qJH8O7zDrKWmNes2Hmtcd8s91kfzBFj5Tdg+ODd4n3I/v7dLGOLdkYEIgIRgYhARCAiEBGICNzgCETB4gafoGheRCAiEBGICNw2CGwnIU5EwJX3KvDJoTQUxOUVRnrKYbEa0tUVMbRO9GzvABPPEKwmQE2IU8fhiQAR1o169jggZAr3LWg4ZA73KbTtkEx8znovZAk6E7C04wIx63ZpA0IyuwOba7bTYonDUHn3efY+9lsU8YLgO32YvGU8CBR/qUKs/6MqToAM4QbxRqx1SHFsQSCxNwNtekexhR/GxY74p1UQFSD1ITohpCHgnZjc4bXAzyKGx2RxhjrMHd9NktMfxDF20653+DN+b+mmzUbIleuhdndDgsWmrIQghfSnPeyCeL3q0c91kKa0ST2wgpjmM4Q8BP0hFch68jBAStM2BeEJghdyGDKYOYXoh7wHCxJN0w4YgSUkPeKDyVxEAMhhCz54BvAcz4MB2FOfuWEciyqIA/ZA4HlsxJbKnokymGL7H3DNig95LJpCdaqYfO7XZ8NnPz2dlMbzfZEAcYIzXhzY7udNjjsXC98hZimsJ+x3OCGHlUKQsVDEGPAKQagAT4jb7wzGAAYcCGOMEXxYb2DE2JhXE7xZj5zBY9c8YQ9Cz1Mq9tDpj6y1taGyHjqtxkXNN2GSIP9ZX5+Rp8UnmpulS+1GcUPeEIgszDsH2DpBOd+xyevQ94eNqqmNr8pjQWR+tay+FwfjYm1fL3Fvbxv6cFg7PktYS/YqlFOiwvtYzhW7o/K4SLT+mR9wxduG95j3nLnhMyIj7/7/pcKcb2nsS5tLtUT5Nx4tVdsliR1f13VETNq12Jsd42av113vtpobm0vnDnaaW7wbV9zXl3+i8tcqjJ15vhUP8GSN/xcqf3+HAbJ2eBd5J29VDG7FeY1jighEBCICEYGIQEQgInBTIHC97ts3xaCikRGBiEBEICIQEbgJEYDsU+6KZHco7aqF4kg1tC52Q0G8am+zFKp3Q645/4PJTp6B6LNgwbC55tBCDjkDGQtBx3V2h3Md4ps2+buAd1dz323am8FtOFyQRRBscSgnnof4RdjgOchZ7nM4sTGfszkmIDizHhsOwTO889zfXZd2TI5ClGEDZ0hv+v21wXeuQcY6LBRCw5dVII0/khmzhRHapQ/bRbsQvowXoQMcIPchpamDGOKcExY7PAa3Y68Wh+OCRLWnAIQzeEP8Q9p7TrnvnAncr4dCrafk6/K0KdgTgjrsLId4vbRT4m2EioF92M/8g4V3lfM89iMO0AfEMUQv7dujwvlUuMfYmU+IYZ4bhKvq1+Ua6wi86Aey3yGqEHY+pAJ+7O6nDdri+odVMJJnnECZ78wb7UKcgwntFierhW3xZlvw+K4qEnapf8ijIhRVDlWSrdVOmlceC3CH2GZNIB7QFqIQWDBHrFPGQH9es17v2O4Ew/QPDtjoRPNeL9gCZvTDeCB3EXZYG4yXfriO8MPYOXgWzBFvEH/A/noOsMGT46JbZ+cAACAASURBVIsqjIVk0TmFLlJYKEUOK1WVfLvIWH18evDhBxIrfuvk0/tevufxV0/Kc+G7uo6HDHZkDzCwmMF1i5TZOtMaxYIujOdL3SUJC3+jz5D6CFvv6b8r2o3SA0uvT52pjjfTUq3d6HWTbi6fTGhV8JvCO4zoxDzg9UQIMoQz1g4eI16TH5rct/qpxma52KoXNy+dnK431suIc4yVdceZd6N/KA/IhVZ9/bmNC6c/3pWD2w65KxCnWOOIUMO/VVmcbvbP4OK8SDuNhTXEu+h8Nzf7eKP9EYGIQEQgIhARiAhEBCICNxAC7+k/LG6gcUVTIgIRgYhARCAicNMgoJA+kEPkfCDsTy2M3N0Nudq0PotU7aShtLsYcjmIIQg2dqVDVnKY0DVhzjWIWBPnji0OMUpxaCaIJsg+iFXagtiFmLaXA58dUgohgmftNUEddpXzdwjagLSzRwD1IHEhYyFrbYt3lVOX57Lhquz5MRjS5XBJfLcwYWIwu4ObPukP8pBx2D6weE4F4cLEOvfxvoCMNX7epO8zbTucE31Dfi6oIIJQB7KYnetOCG7hIWu358GiB9+dJ8R5GiBUsZkCTrTHDn57YRgriyGd0Nm4EJqnNkN+fE/objisl8NO7db6WZNoATGPNwUnk+8WBJhjxsP4Id95ljViDxBELLD6VRVEGeejgIzHLnvYUId+CHUEjhDV7HBnPRH2iDYXB/1A4PMdEp/nINoh6/HaQBiBZAYLiGXWGFiBL7jwLPfwTmDunG+A849U+ju6+0BppLDXhIU62QgPPLkaTrfScMdAGWMNUiBewYA5oI03vRNoY9tO1hJ1EDb4jsiA3XwHR7Dy+0NdMCFklsUJzqxtugZDDp5nHNRDBOE9Y869Xt8Sa2jw3NVOYEQfYIpwpqwmaSAslDwB+l4WxepIL19Qzpsrjz0awV3tZnGP8jh8uZAmz8jTgNBQn1Jh/pz3wp4mjBMMdvLErmmmHte9s7XJrYm1c+PHOq288bGY4/WPFXhCMKfMAXNtQcSeElcdsgSKs/KOePri4vSkhlmSt8Wm8nAcVwJwhBba433lNxGxgveUpfDbgzFh+3E9V1Ti7pm5hUsvXlyceUr5MMaTpKT2EtYB6wsB7bJg0eu2a5vL597XaTd3D4XYwk7W3f+iAk6LKtcrOF11rL/sG0P5K8CO+QdfwrztdPxYF/H22THBxy97PLH/iEBEICIQEYgIRAQiAhGBmxuBKFjc3PMXrY8IRAQiAhGBWwcBdgwr/M/oT0P1zrlQmNeO+kSJtsUdJpMV5TKAkEcgsIBggt2hl0wSWhBgBz51TLBDljp0B2QUoXogqiFenTOCurRjrwR7AdAnxB5tQMJCONMGxCt17REA0QlpyO5j71SH0KIuZCWEsb0OTMjb+2CnmaSOvRUgz/jMGfEBYQRimDjyXIfE5Qx5jp2Mn+/Y7pBQkKV4BICLxR57fVgIgIQ08YxNiAkQm4zDNpvcBhOLR9S1F4iFFc70B9YQ7RyESeJ5bMJmMLaXCPdN/lpIafa3eVcPi1RuNnS3rF6YM9rFNsjbvx20zQkbmQ/OTmBOXex0CCDmEIEBbwmIbz5zpl3mDXvAD4z5DoYIDOBNfxZEwJD1QqEN1oNDISFOgDdzRXgmsGL3P2uMfhAljLlFJ+457JRDFTEGC120QXt4bazKs2Kiv3iE1Jp6faOVHt5bDp862wznNruyWyT3YCz2KrJ3B7ZZtGCt2LMDjBgLOHmHPvMAXtgDOU4bXgdc5zPvJaGnuAc+9lRiLXKf8SL0gCVt0z82eb3o49s6sBMbvq0CMX85pFGzvh7yRS2NJJfLjxQlfCasAR/7RdCHtXNj6woNdVGhleSJ0Tsm0eIhVbjsqZKp77W3o1EKs7TW6+SeU26MvASQPx7YgQBhby17J/HegAvrnNBqeKuwBrDNwtlOooj73aN+PrJ8ZqKWL/TC3nvfmJcAAabYx/whKvEO4FEBsc512mPtFjSrc71OfkkXS8VqeyZf7KwUyp09IzP1b7S3ivvkcfFJ4cI7wCu2kna7y82NtbVeu/2+HcQKqv1LFd4D1uutmruCcfIe4Bn0eRUEreGD8fObzrvImo9HRCAiEBGICEQEIgIRgYhAROA9ReBn/SPhPe0oNhYRiAhEBCICEYGIwFsR0O54iB8Iz3kRbFuhducZsYm5UKi0taMe4qijLdTapZzag4A/u73hIBtGiMZNpEKGbufE2CaQHbaDM8Qyz0GamqjFhu2+roxDDwHofBPUgWSkHl4DPGtBgfZM9rJbG++GRRVIfshqPtMW5LC9GLLhVOyZwBg4sl4PJsSxHfvYqQ7hCREKIUrdIyoQ7tgHiezcCvQHuUvMeQhj7+bHVtvhvB70C/nmMFN8pz7jhmSFuINkB1Png7CwwXNZmz0GY+QEw95t7jBNkJ6Mx3PqcFsWobbnTomGQ2F8PCSVMfXSFfJg4vj/hOLpCyQD7wpssgDFZ5O4VIE4Bzvax/MAAYK1h7AAvi+qgCuCE6FvXlEBY3CEbIbcJpQQWICJk2ND0n9S5TdUII5pE0EGnBgDa5d+ESPIK8GBiGKhxoLEYV0zmQ8pik2IYAgAvUcOjDNuyOg/1aD+IY30GX89nU/6IsVTGlhzbznpKkSUBQREFOcW4TN9sS55R7DNni1gz3XatwiBLfSPKEYbjIG1D/nODnOuOQ8HWPJuURgnzzEe506xgEc/jN2hqH6mOMAYfSjxNuPHxpdVvpW91+u0Q2OD5dQ/smLF5Wqddn5CIkOl181pvtKHdYNwZNkDzxkO1s+Oh8SKU1trlcXn/uae+a3Vym/qO+sCMcfJ7C12csZjhnUKjqwP1oZtA2PWmEN9OYwYc4Qo0T8kKEx1moWw9PpkWL84Qh+7ZT/vuD1m+L1hLYMp2DBXzH1OCbenlaj7Ho17XGLNlJJv3zM6szkvb4tHZw4ufaxUaymnxaCfTqfZWF9+vbm5hoiz04FHCu85/fHOXq93zFWaveEugwi/G/yu8N59WYV5zB68e3+qwrtyq+Jww01MNCgiEBGICEQEIgIRgYjA7YRA9LC4nWY7jjUiEBGICEQEbkQEIC6fUIHA2698FcpjkYN8gyhXrJf1C6E4vxSSPOSwEwRbKPAObXtXQDBBkDokFEQiRCAkoEMQQS6bdKMd57Uw8U2b9pgwcc4ZYtceEuBo8QKb6JPv3skPCfmfqEB0LapANEIUO+GxRQgLLLRn0cLeCb7G2aILdewp8PcGfXLfdZ0gFyKNZ6iPTY+rQJZiI7ZBPEKmWzRxbgWHoHKb/D2JMYOX4/lDilrcoX17WTgcjsfkObEYAQlrDwOeBxuIf9vk8WfD6UDYV0K33gjd9Xbo1W2Dx4ZdtI+NzDOfwRi8+WxvAch06ljEsjACQe38FKwvnkO8WFDBEwSRx145YOKQRtjFuoWsp02EHXuLIFaw1iCjuc936jJe+oJVR9DCPueX8I576rFmue7EyPTFc1liFML4qwKsraTbRZJuKwjS7ntHkgOdNN281A5Pl3NhRddrmhRwoU3EAz4jNEBwc81Cib1SLCYwF/TnnB8WF7iP/YyVMdqrh3fI4doQz7AfrOiTd4d+aYs+v54Zi4UzXXrbx1UJYlHuobm5EnL5vPTOkWZypZeF8jMk5QvHZ4/O33W+my90m0mh9yfq9T9QwWOFg/m62rEm8eBfnj8++6rKR5UT4tcHY0M8YV0zFuaaAzwRKRgzuQ54H53fg/VloZX1iwCEl4NFEoQuBAkf3J9Rku9w+oU9ExIr7pTo8MLMweVRhYbCK431DtYIa30BU3aOyTNjrdMqtOrL1VEJHdLycucrY81xha9SAu7crJ69VBlr/KSxjnBVfEK/FGP5QvGRfLGYdJrZn6C+GVxAeP26CqIe/d3KRD2/e/weMFf8dhAWzQfv4ldVnOclcyt+jAhEBCICEYGIQEQgIhARiAi8NwhED4v3BsfYSkQgIhARiAhEBN4pAhBAkHRF0WK5UNyVhoL4v54i8adkfW2fDIXq84M6JgTpy2S7ifIseQ75B6lG+BKIVEhFdpRDPiEuQDZBBPOZYpId4tghimgv68EBIQkxS91+2oDBZ2zxLn4LHRBeDi3FDmzshvg2KZkl5bO4ZZlChAWEBIeyguylbwslFg2ww885Bj9EKPchTckNYoHHHhRZTwr34TwftIfgw9m5FRymyaIL4+Ue4wQjig/bYgHC+ToeVAUSTWMb7Zsw5352Lo2nr2k+klrIT3ZCcWZRNTeFtueNuT2ua1ncHJbH5D+kMbaChb1cINvZie61B5kMuU54HXtdQLwvDHBkfTLnCCxcx4MAQpOx0AYEs3f9s37AnhBYfzm47kTI9s7ADrfH+Hmews542mVOIKoh+oe9fhgr6wySnBA9oajZragcroYHHhlLDss/aWV3KZQlWhAqi3fAHkZg4WIRzeKZRSvsAB/WjD2P6It6Fia4B072pAAD8IXwt+iFkON1gsiFaEif4Idg4hwRb9vDgrEOvCwQAP53lS+qXJFDQCGN5GmxEpobq2eUjPtJ3Uf48VHaXKl+Vh4Sk7IMbxmEUjD3wTrOigW+zvjOyNPhwukX5meWTk6V9bkgYQDbeb932gDFtY+qEDIKrFjvCFv89tAnv0dgsBPxDXaEG2LuERz7h+wObxzbNSnBZI8+0z7rmgMx8J/Srmxa6yqnhvJdrK6eGzu1uVzrlUbatSTXm1Ky8UPVia2ZXD49nS+0f1CbOH8mTVvn5Z1yst2o1xqbq6M693OCDB0Q9F9XYT0xj84NNFzvVvgOrqxj1gG/VyR2zx68cw7r9RZl51YAII4hIhARiAhEBCICEYGIQETgl49A9LD45c9BtCAiEBGICEQEbm8EIH2c9Loe2hfOKyTUnpAfySnxtsjIbi8koxB9/JkNuQdJ7DwVWa8E776HxFtUgYSG/OU6O77xoIC8hcAn5A+EFEQkZCJ1YOkgP50M1yKEE1dD0jrEj3fvY7s9DLzr32GIuAchCfkLWUnb2A+xSx0T8tkxcC3rdWEPD8ZkYcB9Ik7wLOQh92jf4gX9QXrSN8l4GWM2JwF4c9CWc144ATTtut+s+GBRIuvVgq0WTjwmzwPtU9e4YBPz4QTP2ONnaXvYa8beDJdC2lUuk+aaPC0Yo8M62eskr9mDbPfBfGA343ffzCn9IQA4YTTiA2uC6+AEiW6Bimepx/PMOTutOTMeyEo+QySDN/1Rl3nledYa4swnVLCX+WHsrEfWLp4WDlkGcY3owjOsswUVcAQX49wXdOQt0J8LwkIpQbCTuVfIX6FwUKEh1En9vKcUpuVZ8aNdpaS60U1fP9Ps20u72GahiLlmjLRtYcoCHt2AMWMENzDDXtYuWOENwDyCH3P95yrE+6eOk0HTJ+Pg2WMqXxq09UmdEVvoExsQZTg81sHXa57Ae1Hlf1Rh7j8+sCd0283QWFsmTNbhYqV6Npfk8sLucoNpNzcnEn9KyasRTyCmmXfPISHLwDmb14Jk6RI/krryX4xLqHhZ3g7ZHffXMpZx8puDEeDPmqAfREzmkTmgPebDB/j+UIV38VMqrAc8RMLWajWMTNVrSsZdVtLvEwr5RDtg8Jvb9dLJbju/2dioXMrl0v3j8+sznUahVF+pViujzY68M1YKpXavvZWOK5/FdGW08sqF1zrdrrThbkvpYnqKuNa7wnmCOWRt8JuJQHUrixXAzLp1aC3e2eGDOWEembtb2ctkh6HHSxGBiEBEICIQEYgIRAQiAr8oBKJg8YtCOvYTEYgIRAQiAhGBnRGA9IHsrYvSuyc0Tq6F9vJaKO2dCflqKRTHJFwkznUAYQqRygEBC1FnLwAIQXtHQLRC+LFL2ST5dnihbXIYApl8DJBxEM8Q0xDJTowNKeewQd6BTr98tldBdnetd5U7fr3FCIhfiEgTW45X75BVFiuMjIlbb3HGhix5TT17bvDZnhL2doB4dyx974jHbghkDuzDBoe2csgniHOwyYotjMH1edYeLJyd78AEP9jyGTLa3iM8bzGFtiGZEQio1ydgBwdChQUSixZvijlp2lUoqEbYeLoats4VJGs49BMEeV70ci15InQV88YeMRaz3I/DdUG4Q0SCh0UvJ0XGHuyGXKZd7KUOXhf2qmGMEM3sqF9QQcRgLfEcuS54hvk2kcma/rqK80ZAqjM3iyrYiqcB69pJvekHG223BbRhDwtVuYxxnzwuq7VET3VBLQmF35gJYy/Vw9gr9TCrWwVdpm2LOrwTFvBY+/RnbwiaY60wD6wtRCNEBd4hRC9CjkFaHx88R10IfdpjnIyJtc1zeEGwLhkjeRF4t1gf2IHXA/fA7AoPCQy41iEvi+4HHvtDcAZ3vCwQHRBQ+ke33Qrtxkbo9WbukFrBnPjYkJAxunZ+7EO7j148rkTUl6QDsSYtnDFnrBe8b/iNYG4beC20G8VUCbaXFWYJb6/PXcvGzP1saC0ug8OdKsw1aw37eG+ZAzB0Pgwwe0rlayqsnX7ui143CcunJ76nkE7pxJ61k+Va6+Ekl7JWP6534aySbL8k74vDW+uVPQr/VFT9rsJDpeOzG7l8uXOi20mXO41mrrGeVv5/9t4EyLLrvO/73tKvt+nZF2wDDDaSIAiQIEiK4iou2hdSlCVZiRVHUiVKyeXYVhK7KiWlKuXK4iQlu8KK7UihVNpiO7ZY4gKRokmBJEiCC0AABAiCAAYzAwxmn+m9++0v/9/r9x/eafQMZume9bvk4b3v3nPP8j/n3Gn+/+f7vnajvXlx+ujPNOZ6O7ttzRKEHQKi/ODgu/CU0l8o8T210HlK9zUe5wDHZZ3VohKWVv6mLm8wa458KVZc1kOZjUsEEoFEIBFIBBKBRODKRiAFiyt7/LL1iUAikAgkAlc+AhCjkL8d0UAHo9vaFnPfW4zadQsxtLkTlVtEnkLHniRVITxh1ez331YJjkUAAQrRZlEAVz3slIWEhSyENCY57gDlQRjyNwFlQFSZlAJd7tuljl09mby3ZYZdPXEfcpiDcixk2BKB921BsdyyoihWUD/9s+tK2sVzSNoiFt4dT30m/n0NLpDzEKJuH/e8g5j8lMfZogr99M577ns3tdvG2S6eKMfucyiXflvAMAbkN662vLDowzsm422l4veWRKGe2t9r74j29ExUJoZlaTE7CO1NGZDtEOXHe587uUPfW+khgi1+QJzbSoZxhxS2CAQJy+52dtojHGAhwOFg5s5HWeww50ybeYcy9w76TVwIyPy7lRC+cKHDnMJ6pRjTwrv5aQNEvvtLefuU6I9jVjCP+/gULQQG7eOEkPBHApE2v8eTaVHIiHf+wNahmN40FOVjrRgSB41IgaUDefskvBJtYP7QRgha8DRm9A1hAoIazCDYeQ6hz31IbHDFkuTtSrQVscfWLwgStJ24KW9UshhjUQkcwIc57vmhy7M/BqIF7aU9Dlg9KKAXbbk2qk8fHypv2r6vMlSj/dTTFy8ULLu2MD26aWKoMynin77SR74XtIs+I9Awji1ZNTx7+Lltjyro9R3Th9cTE4JgyxYAz6bBXsPOCwbgTUwIsH+tEmPBurMAyRjxfQJvRAtEkn/kAiSe/NzRPVuekVjx+I47j3xr/ba5H9EKaElYqckV1A5ZgGzSebg+O9JoLtSmxjcu3Lg4Nzx79Mnrnlm3+dh4tzN9U3O+e9viTOn6xlw7KtVSdNuvECuY03+qhDhFoHhwudqtK/h+IVIyr1eyovmy7v+Rki2Dzmb8M08ikAgkAolAIpAIJAKJQCJwzgikYHHOkOULiUAikAgkAonAqiIAUbjkYqanHfi97mxUxkQIVqYUcLspkhrxAVIRctVuUyCWfM+79SFITbZDErNTGvc1S8G7f+D+BlKQ9yEFuSbZfZCtKiyKsAua9yFjyWeS165+7H4Igpud0fZtDrHnHbgm8h3Dwq6VANHbmZf2xi/9tlUC7YdgtcVC0YqDsiwOuAyI0eXkKIQw5RbdLVkwsOUIfYbIpp/kp15bYDiPhQALLrTRLpl8D8zs7om+0W9bpVgAMgbF8iDP/Zu+0B5wRXQYj077cLQnq7H4wqR6bGsaXHuRb1xvkq9P6svKwoKMg68zD5gDCBKMD/UzbzhTFjEluG+LGvoPkQ5ZjaAA/u6H40xAMtNXrC2YB9w3Ee92M2ctqJGHNiIaUC7toc97lcjHO+DG3GK+Qb73BSq7gdL18oN+OsZFnzz1lm9cQ0224mYJFS/cMlI6unuhN6xbjCdiCGMLOY+1BO2DhKZex+iwyzPygQMYO3YKeUn0BfECERBXR+BE+ZRBPyjjPiVwQYi0+xzWCNe0HZGBvhfHnm6c68E47lb6mNK7lcC2f+DWqD47ualUqXTGN+2YKpXLWzEgkEAxN7q+3pbbpOG5E2Mvbtgxyzqy6x+EPXBhDP5SAsAukf4vvvDILROyWril1yn9qu6di1jRb4qS53exf8wrYmggTCBWMZ8gy8Hc64t56zGx4NcvQ+1/3eyxdb97w12HEGTBflGzf//UoQ0PHnp2+zub87U7ZV3RU7yK2dZitR7lzlCn2X2D4lVsknXFnbNHyzF3XCpHXWKFrDYGB+PBt/hLSsxbxApEPebYihYFV5F1BRDwncRahTGzeFkcs+KaO8UUpZgprxOBRCARSAQSgUQgEUgEEoELRSAFiwtFMN9PBBKBRCARSAQuDAEIO8iwMdF6i9FujMglFETkhGJYnJBxxXW6DyHqXdTsOia/XRCZEITY4991CFiIJ8hRSGlcxbA7HiIK0hZSGGIT8tX+9G1VYUKdZxCxnLnHGRIX0hUXMg64DCkLeQuR5UDMtANSmHbyHm2F/IW8hbSGHLXrJLtcMt9sIr0ft0CJXeyQkbZ2cCwLb6jXoz6hbpKT395BbxdP3CtaSJid5Gx3OdRLGbQXDHkX8pLD1g+2LqE+3vU74MzYgCt1Fy1DKA/C2+8Oijx5sphCHSbTEQOWiOySzr2FmWge2RFTX2Q8aBd1QOQiHIDLiJCifIs4XIMTfQM7cGTsGScEAw7npUyIWbvjob3ggCDCGDNW9MvxDsj7FSXGZUkwWaoLDPYq4UqI+xZMTMhTPvXbqoLxtQUQZdl6xkLYmcSKQRf6dbysF/tWJ/1BVU8Jvn3baOnH5CNrt2JZfFW/982rNj0CV4t8DgxO29ntD1YWXVg/dhVmF2NgiFDBnGZ8OYOJ1wUYWRzjmnFh3Omb1y5r0AciA+V5Hnt+FrKc9SVzB2uFLyr9UvGtbrsZzbmprdXayL7hdRtHS+VYmNg29zUJFm+sjcptVKP6mPLvWlaT5+RTsqZ4+PsP3b6uPjPyXyr2xXtP9ZZ01u1bSazgZcQecORgTjNHOTOuzA0OXGwxB7FoeVIJa5X+gfhSrcnXU6+0Q6kp11ZodrdVh9rPbbxuZqusQqZnj48tlMvtzc36euk1zeHF2faNR56v3FhVlPZFjVyniViBm6mTfWF9YVUBnvuVvqfUD/wuYeJqJ+gZJ3DHuuJXlJYH2wYksEBos2XUSeDyIhFIBBKBRCARSAQSgUQgEVhNBFKwWE00s6xEIBFIBBKBRODcEYDYhDRdL/pyA65NYu7Jaqx/y3jUdkggaEMuIzB4RzgCh11CUVuR7ITwg4S1KIDAgJseCFRIWQQL3mc3M4F1KdMWGBDN/F1g9zU+Q8wiLEB2Q/hCKls84V3c37CTH3IWMosYB5DdvE9ehArEDEhidu3SJvJz8D51QvJSNqSl++PgrhYreJ+8RRdLtNlWB7bM4H3HJCiSpWBWJB1toWGrAvpEfu8wBy9IbuNu90gOfO24CPy2uxj6A4HsshBy6BMY0m7KsFslW5pQJ+Q1Y2Y3SEsWML3eXDSPbYumtoN3O7iIooW0izo4eG++IFiAgeOa+Nouv6iH98DfcTwYO7C6Q4m5QZ8YPwQRdpdblEAcYQx5zzEpaAfXtt5BjKCvjBtzgblIfvpkd0vMC9pMueBKjxAFPC6mjlckhxVsW1n7B8/pC+X9mTq2X4G3/3uAJZ7FeiG9tRa3v9yIR68bjn17F2O/QhQgruDmxq6PWHOMG1gzhxCMqMAWQbYMoe3MV7si4zcWAfSRMQNf1gbzE5dKzGNbZ/DbfcF6AAxpN3gjJiHw8B5NX3EHv+6f9oBEVywL8Kc+gn9D6ONiqX9gcNOqL8b8sYO39KL34PDoiIJnd09IsCiNbli8aV21CynNmkU84KANjPtBiQATslQ4PHVww/sUu+JNZ2rHeT6zWMHruBOzdQ798XfJAgb4n2I9hXjSXKyFLD+OKfD2NxSA+4OKZbF9801T/4nEmP1H94y/3G7Ella9MdKYH5LFSWtduzmztTnHsJaijVihYPW9bowq+cDd1d8oIZAwbszvcx6X88TjUr/G94E1wvdgJbHif9b9Lyqx5mxZd6nbnPUnAolAIpAIJAKJQCKQCFylCKRgcZUObHYrEUgEEoFE4IpBAKIUghsiF3crlWgfa0freDvKQ70oj0KMQuhB8pqIN9ltMtQWCuTxTuU+f6sEQ/cBJXYMs2PZhDZ/A0DYukz/TQDhDClrN1EQ07QP4QGiijY6dgR5sOCApPVOcghfW1jQBu9M57kJbdflgMO28OBdx68wwU7ZtiCgDL9rt1buu90+KUv/8H0wIq/PFjbsYoq6aZfJajDkWTFYtXd8O7g2ZYEJO7FpE20EazBmh7ItDHBXA5bcs8UL77oN9J8EXhC1JvkZo0p0exujM9uO+aenFXib/lA+hCHPCUqMn/3vqafe8WzxgP67P9RLuxEnEIzon2NvQJqDDe+DH/kg38GD92xBAKntHdiMJ/nJi/hhF1vMDfoCDg6eTV9pE0Q95ds6hTop21jYSqg/n08Ts4JHxcMCFP3ZQuE1/U9TramppbeOlOL6Wjy2vRZP/T8v91pTtGKprYgMjBnv4WBoSAAAIABJREFUM9fBFGEJkQYSHXKcvmINZIXEYh5zjzysI1sfsT6wSEHEACfG8ttKtygZ6zsH9YEDZZOP90h9l14jH586rZVF/SMM08rHQLRgLIgbQlk/q/T3nbsnNr7VXIzZQ/uGm+PDx2+8uzO1ddf0hFxDXS+LBIRQ+sk3hn7Rv00SA56qzw6PTh7Y0O52yghRjC1j97ASrqf2KoETfV2toz+OSog44MUcsdAK3tRPYr1KgCjJLVT5eLtRrTYWatslwLCmpjWotcpQe2Rk3fRCa7G3rtNsb28uzm3B2oS4Ht12RwMvqJe+nF7XXH9ViXXBPeYJ/b5WxAr6D970HfFrpYOxYYyWC7+rNf5ZTiKQCCQCiUAikAgkAolAInASgRQscjIkAolAIpAIJAKXCIHe5/sVQzayu51drXPi0jZqV/2sYle0o3b9hijXsMCAHIVshiA0ibaSqxXu2W0QBB7XkOUQ3JCluHNitzwHRC3PIaft3oj7EFJYYUA+Q2LyDKIQIpv3IS95DnHI3xEWA3hmd0YwrLQFQpvyIbogZ+2qivJ41+5nqKsYK8GxIOgr/Yekh+SFDKc9EM4Qa+QrihH62T+8G9tEOPeoC0yKO7VdP+XRRrt/shhCG8GIfHajZGsT2kVQZXZjewc+/UXoAB92Z3Pf41HEysSf2+u/xyzYDHaWN8ejOzcW80+diPZCQ62gPJ6xE7ofuLr0wVcQjI4/QpkWZajHlhYWCxx7wsIGc8xCBCS23XmBF33iPRLl2HrD7bXFh9+3ENEn4SVA+Dnt4NlKRPD5uNyhfOblHyp9QLGT7+iptTWV1N+iX4m7R8sxua4Sz0mwsChBXxCawJKEqET7WCee02CHMIfrJu86tzDDGfEO3KifvAiCCCHMR+Yy47tH6d8rsW7BmvqfVXKcCQhx8oPlBRHjgwDclIegQHtPCha6xtRCBjqddzQWFl979IX2H93w+t4LGyXPlCp9axpw5737lbBAWVicHv3c8w/f2pg5PHG7hAHPObB5b7+8JcFmLQ6wpE3Fw+Io30kw78fQkAsoWY8Mbel2S6PqwaJiWnymXO7KcqJ3b7nS2j0y0Xy+01x8b7db3oJQ0Wm3ottaUq1WOP6J7hHcm7Fj3BB+fuAoai16evmVyZK5S4m4NssPRCTWmAXHU57ft5NPYR6JQCKQCCQCiUAikAgkAonA6iGQgsXqYZklJQKJQCKQCCQC54oAhCckMDu08Zd+vyjQanTma9FdFJHYVdDt3l1i5+xCCdLOu5otWJgAtoUBpBv3IPog9SHMuYZEt9slxAtIae5BACJM8L5JY7/Pe5CpELCIBhYgyGuLDxOuvAMBa0GA9lE+RJjFAIQBu9YxmU6fuLYlBuQxv21xAElJHoQPyETaACnr3z9ZaLcu+0eRALb1AThwFK1SaKPFE7uIclvpF8muoOiXy2A3Pm1iXN6n5N3xPPfObFwA2XIEXKgXsh8M7ObKdXinN22g3yJhe3X1Yi46CyMx/ThiTU212PKB/kMyI5YUD/fNliveDe2xLQoMtNniA+XxDNzssqoloaErt0L8rWjy1v2kXPrv+roFq4gi9ucjQizr0ml/UjZtRoDD2uUB3fgHff9O6kFbrZjrROmlRt8dFHhg8cC4sQa8ZshuiyGLZFhHsMOf+xDzntMIHZRjKxtwYQwQjn5ZiXFjfvLee5QIvP2tQX7yWtBjp/oHlR5Usssx8D0tm35aBAoPBqIF5UEu/7HS313+Xq/T23Lk+fJvPv35oX98/883x0YmejfJymJI84q+0fb9cgV19PiLm78zPzl2h6wrsNZAcDkZzHuFtrA+qdeBu8+mueeaB3z4LoAj37Sm2rmtPjc8O31o3bPrt09X5epqR1R6Vc3D8VYjNj7/te6vyh3U9o486nWajb57LB22AHL9X9IF8/U5pa8PnhdFvnNt55WcH4yZAysJNQ/o/neV+LeHNbeW6/pKxjDbnggkAolAIpAIJAKJQCKwSgikYLFKQGYxiUAikAgkAonAuSKg3fEQP3tkaQG5acK8GaXeYozdtl1Bt0W99kR0liBkeQ6xzMF7RRLZ4oUJ5cEO/b51gne9QzbxDtYPXFOmA0Iv/3uA8osulSCx8XMPMQm5SX52n1POzYPfkPOQrjyHtGWHvgUZSH/HmjBZzNkujLAw4YDsJ58Jd8oiDzvTET94DkEN6Y/FBuQveW0FURQj6Dd9BAsHUoZ8dTtom9vnc1FsMVG/5PR+KdnSgLot5nDPO+2JWcB7JIs+dmcF4cp7FhFsDUM53OO5Seu2fN6MRa+5MSqbZqMld1BD/bFDaGIXPCQx5WIdcPIYiAbiZvte+Y2hXevwflFwKFqc0IciUes2UnZ/nqns4j1uXZBVQLHdZ3vNTu5CHAteAy/GGFFhsr8I9D8VtXQwaBM3DsfzG4di2+Fm3K3bzEMsi+gTogSCEzgigmEBwfggzNn6gvlC+UV3Y8w9xgqRD3dolMcY0gasPQhkjbWUrZuYe4gk1M1YsGbIy052REPmvgO86/L8DsWy4EX6BfmOZQdr8KeLpcHZt+qliRcfr/6KZsi6176nPTO6obdYGeodr1TjaQXl3iGLBK2x9gQuoSQKMNewIlp+UA/ri36AGaLk+R6UY7dkFu78/aFM5hl4m0xfL3FiUuNc6zRah/d8szQ1f3x09x0/3DzUksQ3d6K0Sf374amDjU3tpoo+NVK424kLrP9NCfwZbzBjylxrVhX9MdOaYukwh/m+rmQuYWugfgDy4kCndcX5Tvt8LxFIBBKBRCARSAQSgUTgTAikYJHzIxFIBBKBRCARuIQISKyALGL3N7u5S/pPI1qiDqOs69Gb5FAHl+sQbRCDjqtgQtxEuol6yCQT8ggGEKF2O8N9dkFDEELOQgTiAgQhoOhmykKFRRDQgWy1GyPaAYG1SwnBwLvybTUA+QjBSJstKFAW73O4zZxpr/8WYec0BDFEMP20/39EEghk2m0SnvewSiHAsMl5uyyCdKRM+o+oYusG8HUsApPvvGsS32Rl0VKFcvhNWbxLfoho2odogGsgE/92J0TfyVN0S0XbOGw1wpn3IACJLbFLyZhBGGrsy4ej1ByN5oGX5JW/K58+ErL6xO6TSpDmWF3QPluQDKpYEhd0dBAwOFPeQHDo59G9k2Or+2fc2V9872QFl8+FhR7mARj2D3U7hpSGy/Fzrx8vPb5vIp59qd6bmu/0MUP0IYg0c405avdf4M8YMqYed7BhXjInuU99WAIxBjzD4oV7lImgR7m2VKFc1goWG1haIGIgOJIoA+GQdcT8tqi1GoQ5a4R4DBYV/2tdnzzg77vteM/+J6txbG8lJrZ1P66vzVNzx0rN7bd35YiuXG3MN7udVutIqVJFbDldnApbD9HPCxEsLNj5+2FrIM/RvmVTt9PuC6ClcmVrp1U/1m42NC6lZn22/trnvtZdv++xkbFet3c3Up2CacuqgpF5hSEAwue/GGCD2PfNwXjVZaFy0QW44rhc4mu+kQh471P6pRXaskv3EKYdjPwSNzerTwQSgUQgEUgEEoFEIBG42hFIweJqH+HsXyKQCCQCicDljgCEn60dmqLEK7Fup0SE8pACLYuYHhdpWLIVgYlvyDwT6ybc7UYJgpXd1RCqkKEm2k08YqEAWcvuaZOCRXLQxJ13Obt8x46wlQFtgsCiHLtK4h5tRCjhbwzOkLC2RrBAYVLSMSXsG52zgxmz65385KUsSGGLEd7VDZHsfkPic9it0l5dQwxDxt0xaKPFGPK5X4PXTlq48Ju+0ye76oGYpm0Qs46d4f55TOg7dXlsKMP9pI22eqGdYGgRih3sLsNWEIsiWxW7Ys9z0T6xIYZ2bIz6gbpKpkzGljIYR8b2FYJFv3Ow9j84n8LcXuYihMfjbM620mGnfH/e0uvKkljRB6tdiQ+9cSL+8PnF0v7HZnvHGrIs0G3cMzGmtmxgbSBAMU8R2Rgfxg7LCIQMB9+2yASRzxpCXEL8g/jeNXiX37xnqx/WIGN8qxJjRVkIJ3YvRbOLFhz8vtCDOr6stFcJoeUXigXC4ysGdcyfkC+oE5WP6NlbdW9y9phEsl5srNRKN224vjc6VIkfW6EhrE/a6/XmLLac8pynj3ZHxzo90wGuRdHDllesB7mp6o21m/XRrqKHD42OPy2xYmtzfrbUqs/Xut3ObQqkfVu9P0I/0FhfqVX0hUEsYGgXZ6wsGNtrWqyQdYXdovGNXEmsAFjWFmuMcXmFCvQqY5uPE4FEIBFIBBKBRCARSAQSgXNGIAWLc4YsX0gEEoFEIBFIBFYPAbmFasvKAjJoQVTQ0ShVb4uR2+ai16hEe3I8hrZDSrMTmx3ZuC9BILD7Hhg6SFBIwqI4AbkP+Qohx3MIWUhYyFq7U4J4osyiQGGLAzpYJNxPxjXQ/X1KtAkLB0hfCFqeQ3zxjl0xYc3BrlxIS1s0+O8O2k17yUu7OEMkEsfjHUqQoog4kMLefQ7pSV2USf2Qzg5oTb8sCrhs2sNz8rufjkehWyfbRNvcdos0/IZ0RpxgRzx0KJjaagJy1dhbbKEN3Ctav7ge98GCBuNB2YxP351RoY3US+wSCVZz26KyrhW1HcOxeIB6wIz2gIPfp45r+WDcwQVXTB9T+o0++6+RqC2l5vFWPDJeiaqEjK269ToNMmuDNYf4A/524wUhy9hSJnPQ8UYQKGz1wxy5VwmrH/JjueP1h4hEO3YpsTYYS9yEIb5BkjOvmEdYVNFmEhZOPF/Ng/YzP1hPBJRmHZziHorKCqQ+a2ln35GYjm6n+03hp/Unm4We5n6vt1AqlxE+sM6ZEoazAvgu/ZjSGeEFkcdrnzWwoHyPSxjbqDzX68GirsEZbNWWniwdStRpi6flfR/Sey2V3ZL7p+c67eZUY3bqHRIobompY892Wo3XyARErSsaSJ0Rvk/oKS6lsKp4XAkhsy+myrLimiXgB66gbBGHJRDfo+UHawrMmKvXshXKGSdYPkwEEoFEIBFIBBKBRCARWF0EUrBYXTyztEQgEUgEEoFE4HwQeKFPFmmXc1SHSzF686iCbovTq5YUd7salWGCBUMEOtgz/347NgFkJ8S+SXvIechWyFPegShl9ywkLbuMcV1TtB7w7u7lxJ0tEEzie+c071In9eNiheu7lSAtyYOwQDs5Fy0awMVluC4Tw5CJX1F64+Ad2g8RausQzhDE7Limr5BnHPSROAKOYwCBTILQ5x1EE3AxEW23PxZQLMpQFs/s9spbtblnt1IEM0YsggimfMr0Tn3HMFgu+FAuZZHIY+GnGF+CNkBs8y7kNX2Zjs7cYpQrE9E8XI5ybaI/N5aIdfreF1Akdq1oXUGl19jBvHhCifn9GwZdqyeUbjnQiMWXG72ZkXLUFjonhQgLS3Ypxvh4HCHXwZjxR1xCKGSN7hqMkYU28jNXEfEQkhAvGE/egxSnTawDu49iPvLb65f5y/usJe7Rj1cQ6CMfn4r6R1jW53TQL9qBMEO8BvqAAPOLr1ZKt936e1MH9sTYxq3toZHxXqU2slmzU8YMrbqEiM0SCo5UayMLvW6n2mm3ZitDtUa5XBlRhqZ8NkmQ6VW67fZNrcbCYfJ22839w+s2yZtThQDfEkQ6L0nAmJQIcnOpVJnQmTV6ykFlEi269dkT71icObFB5ek9RIqeMC5C9Aq4nlFBr1MiLgWusTg+qcT4OVZJ61oWKgy04k/0JFrwTeLbwjeK+bv8+H8H82g13JW92tTL54lAIpAIJAKJQCKQCCQCiUAfgRQsciIkAolAIpAIJAKXHgGIy7Yoo9cp0PKJWH+/rCxuKku0ELHd7kavNjLw8QPRTZBfCFWIVIg+dnLbdRIkJQQUzyErH1ZiNzfuTyBXBzuc+0S3gwcvd0djMt+CBehQLu9DrNoNk13AQKBD4lMeQoX99EPCc8+iha0wqJvdzbSP3eYIILSfqMH8hlilDMQDnvGb/lAe15BqEGw8h8WlPK4pk+R4G/yN47gf9NuxJSzAuH8+F60/7KrKQcl5166Y6AeiiftWdI1joaMo1Lh8u6pC7KDN1GdLC132D9p/MLqtR6N15P5oL3RjaPNw1LYfEIr0nzYQP4HxgCTPYwkBxgvi/4eKgCgKTIxWYvuvXFf6H39sS+lff+zl3u4vTfWiq/8qH3OIeYaIYIsExCJEKeYQVhXkIT4G1gW2ZHJw5uL85pp5xVokmDZrlHusGdYf9zlsYYOYwUH5jKktOIrNX41rWz0QQ8OiCd+E33u1wjvNetRnJiVItDcPDavrMrloLsyNlQRqp9V88+j6LQqzUiaoRLPTbES3UqnIZdNoeajWViCMyYWpY7c2F2bukGBxSJlulOjwcrk69AkJDi932437JYLsGF2/uVStjTaqI2NjEjD61kv9ePEy65BFxZgEj6jPTkqk0PDqnsQSxvgV4kahL6wf+vpFJQRU+ox1xdeV/H24pq0qiuNeCLbNnCXWCWth+YHA/Q2lFCxebdHk80QgEUgEEoFEIBFIBBKBVUMgBYtVgzILSgQSgUQgEUgEzhsBiDURe3GP2MChWNg/HWN3Km7Bnvmo3SKSs2R3NJClEKqQ1napYiIe0tUBpikPYg/LCuJMkCBdIaYgZRECIGDtCslWAJwdR6FI6FsIsWBBPRyQjFg+QMxi6WCXIRC+FjiKflvYte42Hhy0BcL/nkFbIYdpK32D1KUtlI+ViK/BgrIhhOkL/bCbJMfPoO+0wZYV5HfQb9ptYcHt9W+eWdDgHQtBiDL8pv2IDIg27p/FDWPoMhzM2eWRD8GFxD0HO7fYQn6EpVntZVf/y8NR3bgpTvxNIxqHxA6fFGPo2xdkXYG4c80d2hUeIlqX95txwhKGefAZpZ90hr5fsHK8c30lnvj1G0vVJ+Z6e0+0+iIEYhdzkHEAU0QG3kdcYJ0xxoyT5xBCE27LKJJ3vYYQtXBjRhnMR8aZfIwla4LfCBLMNbvfsXUHa5L54ODf5D0vYlgWA+7ySufF+9/1dx4Z9Akrg99RepfST5zuJYkD0azPB6IBWoKsKBSsW16aJFJ05YpJ4oSi7GgJyOKCMsqVKiYYIxIX3qB4E8e7rZYEA4kMrBeVpXfvjMbif+v6FES7X54sM2Jkw5aQcKFsHYkieKIiVy9ai/KM1+kslbLkv+p0YgVjhBUFc4Bv0gNKjCHfRqxu+iJTWlW8YrSZh29TervSe1aYC6wlvsfgCsanHKzFPBKBRCARSAQSgUQgEUgEEoG1QCAFi7VANctMBBKBRCARSATODQHITPzNbxOtqR3XzYo87/eiun5ccQxE1o0p4HIVMhXCE8IektBuaWCNIOb4N91BgskHeQpRCuEP2QrBahEA0t2BuSHeIfQgWMnPs76/+kF9lGsyHtbQRD7ubiB+IVsRISifdlj0KLpX8j3KtDsn6qCdELS0xZYR9+vawV25R79tBcJv2kmf6T/XtN3uoiDxHecCLBzHAnx5h75xbT8yxXY5iDbtsXst+sp7DqDswMyUa5dcjmthyxT6uJKFBfVSNmNH/yxYgJ0xoP30a3u0DonB7ZZj6wcnYvKzuNJRLAH1rdR/l7gnZYkW16RP+RWI0q5EDMYbYvVBpbuUiB1RJZaFBmp+pBI3KobF3FvXl5796+M9LJqYM4wd84WxZF4yDhbAmHeOL8I9W0LYOgjrCA7mFGUx/sxHxDV29zO/yUv5lEs+yqSNjBuCCNZCCAnMMfIiJpyXYDFoy2lPIuubEi0QR+gnawYi+uNKrDd21iNm3nxKAUtWDdErKTUUB56H7aWl05TYEPXSQPlb0jaXdIb+/9L/Mx7En+hbZkgAWZw6KkFkuG9d0Y9LgcAhqwpZcixZXJz++JoeIQ7970q4laP9vECsCgtE9LWbYsWKIDIfEYvBjX9XPG58YxDwWEvM1wWtuWvyW/Nq8zifJwKJQCKQCCQCiUAikAisDQIpWKwNrllqIpAIJAKJQCJw1giIeG6IgH5IL5TE+v1wzD+9I0ZvKUVZNGt3SgTmJpFJVQSI7UoQjogEEEyOu0BdkEyQSib+IaOwxsB1EOQT4gLPIaUcNNqWBZB6EH/4fOfZBwZ1OXA3xC2EKofJfNrCtX3vWyDgHY6i1QLlkw+/8nYZZV/+triA6bTAgDBA+ZC3tNmBu+kj19TB+Q1KuIkBC55ByFLurUr47kcEoj4wu1OJdtiVFe2BsPbfQtSFayvHzqAPtsygLg523y+3yrAFBc8tWtAPDpOmrgeRgvGhDtrsmBTUjZhE/tnozIzFzDe3xvCNlSiPK/h2m7EBX/I70Dht85gMqrumT2DPXGLOEyQY8e11moQjimOxc7QcvyYe/B+9bX2MPzwdB2fa/bHFuof14MDpjBP42jqHMll3jCfrgjIZi/cqMZbMPe4x5xAA3qQE+c9YIVjwLuvA1hfMQ7tCQ9jwPPb8tfi1JgMJaS/Rgrq+q0T8Gfr0l0q40vp3g/PP6IxlFsd3lLYNAme/sk2IGf271v/Ordl9gaLTD44R7Yam8uCLgUhiK4tlJfKNZCxYhx9VYn0jBLEOeJvfFgY5M67n17hz68oVl1sCH3Pcc/+/KHQALIkDsleJteTv8xXXx2xwIpAIJAKJQCKQCCQCicCVi0AKFlfu2GXLE4FEIBFIBK4SBCRWLFlO9HSuaCd351gn6vtEuJWaSzEMrpOlxVAjqlUT/3ZDBLEP6chucgdjhsxj9zdkFMQTJDw7v4sxHCBqTcJD6EGU8vytSuzyZocyO8q5Z8KPXeAm4iG7HMvCwaAd0NrWHnZvw/sWFV7UNbvKKRuy1qKGXVOR17vR3S7y0F7u03+EDFtJQAiTD1GCfkKuUTb3wAH/63ZDZTc8WDHYKsXWJWDomBfktxugouhSdJelLCePouus5fdps90AWbxgx73xtpUI4opjWmyVK7Bq1G4ajsqGWnRmO1GqyB+P8K7089g9WP4NV0R7aU440DVEK4Hg+27AGCDiWei/tY3VGL55JKrPzMe8jAUYd+YU44HQwG8O1gD3PO+YZ+SzBQzzBrdQCIE8w6KDZ4wJ85OYCeRn5zpn5hPzijKZk8RAgXxnfZIHot0B1MmzZrvZB5YG/bUp8YI66cs3lcDqr5QQAghazRoCj7+txIGIydpa/aMvfFik6K9jMAXf3x+0g13+DCPfEa/3z+qatcTBN6dveTTIlyLFGUZpEGgbEY3vpee83+DfBdYOghZWdBZSV3/cs8REIBFIBBKBRCARSAQSgUTgNAjk/9nNqZEIJAKJQCKQCFx6BPj3eMlCoiRxYfbp66KyrRHr3lyLxX29qG2Vo3d4ziqkJ7u3cUEDgcduWAhOfPEXd2vTI8g8fOizE/xeJYgoCwXepU+d1A1Byo5wRA92jGOhgIsVdlojBnDwzHEgqMtBtCH/bVVBeeQrEv2OL/BF3YdYREiApLVLpUHx/XeKRCNtKrqGgmQ1icp973qHdCUvZUMW0zdIfchmSGjIZH5DdtIXsPOOet7hgCT17nbaRj/dnqIFxfI2FsUKt91to1zKcbnkdYBwxpB8jBFn7i+1odsgfy2Gb1AQgZe70Xi5E7Ud1eg9Bcbs7ofkBmPKyOMHCIA/64EAwYz9LxXB6asPlXjXa8dLvTdPxNefW+jNSrBgLkDIskufdYC4QMICARGQRQdxzjiCPXMXoY7iwJ/7zH/KYG4hYDAHmUPEmbELJuYfAsUHlVhTzEXmL3UxropZ0h9Tu0vT5dofEi9YN/WBcGE3ZrQVwQYy+3qlP1EiH2IGWNDvHx08+7LOfF+wOAGf9w/O3P8xJcqkj2DJAQGOCyKviX+ra8RU4ijwPvXwDvfAlLnONXXyjHHFYoz2gaG/D1GI4ZFixQDsM5zAmLFEhGLslh/M6y8psZZYU4npq2OaORKBRCARSAQSgUQgEUgEVhGBFCxWEcwsKhFIBBKBRCAROB8EBi6h9oqqkwsoEYW9Zima+xvRPq499VvkzH2+Hq2jzajcJNK+tFP57M4I4g8iH7KUHbN2OeOA0OyehYyFHHWcB+5BkFNG0a0QxCM7/SH8IdIhtSAKIascnwLSkHds4WHrB86OX2ErDOIEQNqym5xyeQ/iEkIXch5SrOiayqSYxQ4TqI4fQV7qN6lJ33kHEpN2QiTTV37zjAQu9BNSGWyol3LYwU1/6Qftgpz1bvqiWx5beRTbZgGjaHHhtvIMHDwuujwlXgZ9cUwQ3GO5LohhnPgPRWdhU1RGh+UGakQO/TVyY6NyDQVp6x38u3RNUOE124VPo6/QA+wtBjDeDg7f746sLO4YLscnbhuN4ztq0Xix3p8ziHi4c2JN+DfuwyyYMXc8nsxj5g3jbFdlCHusPcQMyH7WDu3gPvMdUt3iErvWER0dgwVrI9xXkY+5saYuoU43pggXEi38mDVBPyCqWSeIBl6rxoe1zTPEA74rxJKA3EboZP2zlr6oxNpCTPWc5xkiIhYc3P/WoB7OiDzMcUQf1qkD1Jsw97ovCpmn61LePzMCjAPzEnGaub78YO2Qh7VkUTcxTQQSgUQgEUgEEoFEIBFIBC4aAilYXDSos6JEIBFIBBKBROCMCECYHpBMoJ3FvaMx8/RwbNpTiU231qK+fzJKw8NR3fyICOwfjVIJwtPEJ2QpRCfkkv23QyZCOiEOQKSaMKQBJqAgXclnVyoQlZD57Ly15YDdD5GHeux6xYKF3ddYPIDkchBpk7AQjpSJtQf5uE87uaae5ZYMFixoH5g4CDZthwgt7vblmlQUHCBXi7EdKIN2gRn9gAx1LAm3g+d7lcCLOnyYmHY+ixW+b6GC/BZtLPZgsWK3WM5Hn2kPpKxjH9jaYoMEi9HolurRnh2JhefKimOyGIsz1Zj6Sk9o0S/GlLgCT0rkyuOVCDBOrAvGBxECF2cnDw3CXSPluOPedaWXJyo93J6ZGCcPBDnuzXij3Yt6AAAgAElEQVSfnefM9b1KzFdEDcQvBAvIesYWcewLSswr5jfPIfS9nhy8njnwFSVbFiE+YVHxxkFex7lgDl+yv8sLFgpgAX7uB78J2M23gDn7opLXKPOZ/iBqMI/Bh28I64n5ynjYEsIiIv3EXR33WafkfXSQ3wS5yz8ZgHxZ+2hTHuePAGOBpQ9xjbBAW36wdpgDrIUURs8f53wzEUgEEoFEIBFIBBKBROA8Ebhk/8foPNubryUCiUAikAgkAlclAhDQimXxiKhASM/1Ot8W80/OxPBNE1Hbvi460+PROnZ7lK+fil5tnZ5DIDoINP+ekyD8SJCFkKjLd20XrRNsLYHLFohbSES/A6FOOZCxFjUgKyH0KdtEosUACEa7mbLQQD6EAYhPXLjYlY6tKkzmW0yxeMH40jYIUEhk2gBJzE5uRBNbcBSJNIseFlBcpl1F0UeLH34G+W8f/pDTlE/bIFFpM+23+OKd7z7b8oJyHRvE7zkuxpKLr6Xnxp0d6Qg3xoZd+JCGS8RtSfV3FxSvYlF9747H4vPzGvNW9NozenZIFOIRncGSsvN4JQKMC2NCTAbmySmCBdllZfEhTZbnhsslYd8j8DVzh+DtzDfEKuYbB78RGnBtxLzzHIfEZe2RD1ECd2tYFjA3LJZRN+MEmU8+YgIQp4IDUYT1hqUBsRkg+Rl/5vplG0R9IBisRF479gZ9Y02v2IeCBQfPwcBrlvcsBPp6AFWe1ggB5idWXR8+Tfl/rvusIdZSuoNao0HIYhOBRCARSAQSgUQgEUgETo9AChY5OxKBRCARSAQSgcsHAQjMH1aqi87bHdNfv16Blxux5UfXR/2l6Wgeno3SO+QiaGdDVhbs+ob0s3sPCFYLFPz7bssKE04+k98EIaQ9rlkgItkhDukKwYqrGtyzQOg60DeunXDbYndSLsPWFbbuoG4T/5D3kL2cIXMdxLvo9gn0i1YV/LY7GuqmDbSNdhJM2TE1bKGx3G2Tf1v0cOwN6qBddttDO8nr2BgINGBGfu4hVvDcQWndRpO27i/tdWwRiFj6yI7x1yshTjhWB+/TZsp/QentSow3pPeSW69erxrNl+Y01s0o1+aiXN0a7akFBV4/EY39+6LbnRNSlJ0kIqivfDA/EQcQAHA99F8NxsRCVQ3Xax/cHOv21OPYZKs/Fo5NwRxHtGD+MS6ISZTHuDKPES/sTox5+B4lrC1Ye3sH7zI21IVYYeELsY61iQBCbAbcgf28EnORfHbNdtXuZl8hxsTyOZxzWhNhrQ8F3OZ7hPDM2bGHbFHDN/pfK31qMC+LYtRaNy3LTwQSgUQgEUgEEoFEIBFIBE4icEl85Sb+iUAikAgkAonA1YZAr9cT33xKKvH7XA5ZWUAQEfAX11Cj0ap3Y+abx+LEgzPR2NuN4VteF6Xaluh1IE0hRdmdbVdEEKgQTpBQkK52/eR4FzSlKBTwN4ADdbMbHPKc9GUl2sHufwQD6oJYhXS1tQD3uWfRgt8ONm33SdRrawgLK5C+tJH7CAHFjRPeHU+5JtMgkukLJK8FBwfa5XfRkqLoYsriAKQzVh7kg4R24G3EHrvLou0mpMkHJryHCEHffba44b7wm+e0DcKacrjeOyjb/bGwQR5w5jfl2zKD+4pb0huLTmNY7qA0ibrDEimEU28uGgdnFM9ia5TKiEVYvryU7qCEwukPj9MtyoLFEIeDqKMYndhQjZF3bCxt/u2bSwuvHeuPCcnWSowfODMPEO5sCcA8YtwQHpi7dqHGnGHsER6YKzzjXWIDcMY6CIsKhCrcUOFSiTmOUMKZeeDzVStYLA1DHpcSAYkVfCP5d4JvCXOZ7xUHc5w1wsGaYe1YyL2UTc66E4FEIBFIBBKBRCARSASuUQTSwuIaHfjsdiKQCCQCicBFQaDo9uRsK4TIxCf8HWJXX4zGodGYfGhWBPaGGPpeOzoinda/Y0uU1jXk38akvQMDm7SHnLcPebehePaGBYhW7uPuCSILshXXSBC4b1OCnCVQMGQuB77NdymZpOUMaU/cBghdynDA76JYYasIynA7rObw20Qt7fLfJhBq5KFvuM/hvkUYk2t2tbS8TOqxeyieObA29ykT6wlEGfI47gZlQSzbdz8kMjv16T+uhbCYoF7ag9UHQgpn7mH5ASHNO+zsx90KIgixCrzL3iQ2BPYuJYQK+gUxOCQRSjmPd6I0NBHVjd1ozYxGqSN3UK1GdOtyB9U9vhTfJIPgCoMzHYwvY4HgxnxlPSE8MHcYq7cOl6JcKcX/sXsxRnQGf1vVYMXDnMA9GvMG8haRizEtCguIE8x7DltSMP8RwXifMj03WUOsM+4x3hYUESYZT+aJ3alRXooWA2DztOoI+N8H5vevK90/qMFrg7XCmmHtsCbOTXFf9eZmgYlAIpAIJAKJQCKQCCQC1yoCKVhcqyOf/U4EEoFEIBG4XBGAwESweK8o05J23m+I1pFSHP2ERAsZBkx/Xa6C1lVj3X0bojS6Ta6h6AckKKIDJLiDZkPOQjiZACWjE/lM+kO03qMEaQr5Cunu3eO4yMEtjuMyIDxAsvL3A7vJbSnwpK4h8iHAED0sBFB3kfQqCgtuC+13HrvGQQCBVKOdlEXbHDcDfCy4kN+unSinKBC537YwIS/EHIIBIgXXtqjgGrGCciGnwYG+IUj4fe6DGUIH7aUM8OG5rT4s2DhQOKQ24oVJbKxUEEsgA7leclHV7dWiM9eOXmNDVEY70a0tRKlyLLoN3Z99RrEs9vXzlqIu64qMX8FIn/lgfBAfPq6ENc1vDnDvv6Ulc/9oOX5o10jsPtAozeyr947Od/qWTawFxhTiFrdNBMZGmOL6cSUCcDPHmB8czHnGhjlF8GK7j3pZ11gTMX8tfnBmzFmnPLf1EvOU93JcB6DmafURKFhXIKrhdtBiBZXxXeOb9Ekl1gxrJ8WK1R+GLDERSAQSgUQgEUgEEoFE4CwRSMHiLIHKbIlAIpAIJAKJwDki0I+lILdQJuZPigelJZHhdAfEJYQoO7tHRI8eE3V0PBpHOvHyvxqPnf/N2+U6SO6DTlSifN2M9or3xMDaNRI7/Tkg4CHNIdU5F8UKnlvMQNzgXYh2CFTIdIhVCFiuyQepbhdOkPoQ/5Bb7gTvv0aJ3eO26uj3ffAe9RWtKPyez3Yr5fZSPiQz74MFYoUDZttaAgsQE8KQzC7DdRWtN7hnN0H0A9IZkhiMIZR9DZEMfmDnYLP0h/wc5HMMDEi/pUDZS/cQM0i0C9wQKfhN+X4XnOgLZws+EOG3qpsjCrRd1rgei/Z8NTrNjsQL4dAbjxN/Dcl9pxDE2oO4InmcHQLMHcb0icE4MC79o+//phTH7xov3bCt1qssdErf/cpUD1dNzH3mNqIYY6Sx6QtXzAHmJ/Oc8cbqhvJYN6xT8hNbhHFn7rBLnfeZP9ynDK4RQjynvUb4zfxmfqV1BQOUx1ogwPcUiy++cczX5QffKtYKaybFs7UYgSwzEUgEEoFEIBFIBBKBROCsEUjB4qyhyoyJQCKQCCQCicA5IwBJZHHAFgIQlafdvUp8gt7n+4TS7yn9d0qHxbAuxTloTl0fL/zut+O6//yGuPHXdsnSYjxK68sDwcJujvi3nbpIDujs+rhnwtztsFDBfZOwkOTsLLeIQB/oC66hEAogbXkPstYxGhxc2m5HAKsoSlhUcFuWn53X7nP4TRsg+blGSMBiAUIZCwyLIOxyL7q/ol6TwVzTPltAmBCmXwgKxof+0GdieIAB9ZKXoM3suOfalhw897hSvoUIiD7G7Q2DtlE+cQyo23ENaJfdWiEKqaUKdNJabEVnapMCbFd0VgyLdlexK7rRWTwY9YPsxkcc+YzmBkR5HmeHAGOGtRAWQb+l9O+Kr1VL8eFaOSrHmvH1F+u9dfpdbUv6Ux7WGrEmcAPG3OIec8Dzk/HE6ohxZFwQKRDYGG/WA2OMZQ5zlPeZrwhNtqigHOZMMaBxt/4RuQHLIxFYJQRkUVEsyXOX79B9Sh9ZoRrWCPOZNZNzcZXGIYtJBBKBRCARSAQSgUQgETg/BDLo9vnhlm8lAolAIpAIJAJng4BdIkGQmzQ/G1cbR0ROQ5o+qATZpGDb2t1d0o7+rsjRyQcW4sj/tzvmH5fboDplP68E2e76HHzbxBN1QkbRBspze+iD/e3bbZEtLngXcQLBwPEoyGOXT5x5DiFMEFd2p0P02y2T63GbLGT4bMHEZBr3uUd9kPS01VYaFiQgeSF+IZUd4Jg+FN1L8bsYy8O4Y7lBmznoDzEpHAScM+Qy9+gHvzkjOIAbzxwk3DEJjCcEH/UjePAeGJD/jsG7tB2Rg77ZBRXixo398ns9xSU5Wo/2TCvK1XaUh4Zi5PpWVNZ149gnl9xf9fqENy6J8jgNAvftBPJTDlvVME9wWXaKdUpZbqE2VuM9G4di0+2jpc0SLIpiEkIV4+cYLYwX44yrNq49x21hg5CH9QWWN4gWtythceRg9I6TYeENcQNrJeZQWlbkrF5VBJaJFZTNvOPbhLAmSfwUd1A8Z22wRlgrGWx7VUcjC0sEEoFEIBFIBBKBRCAROB8E0sLifFDLdxKBRCARSAQSgbNDoE+aygVUi430A+LoVd+UWGGh4QvKDFFO0OAx0U6Loq9fjvrRauz5v+Zj9vFq3PZPx2LT+xAzIE0d08EEvsknKrcAAIkK0eq/AcjLM1tT2JLAAkLRWsHl2lqCtt0yaCNl2LqjuCGi+A59d6Bv2lAUK9xnBz0mL3kggDlD/GOVwM52RAOsLSB86TNEcdFyxeXyzG21eybKo50Okk157IYn2LhFF8egwOUPbrNs5UEfeY+2eoc9beM+v9l5z2/EC+oAHwQM2g5JzW/EJXbs7+/n7c5tl0XFYrSmFvuiReNwKcZfo7gWjXos7lkK7lyO/6iz26/LPM4SAceUeNcAf0QExq/vHkoixftvHint+/EtvYONXmn316Z6uPTaNUjMQ0QFxhHsmbeMO3OB8WXuIdZ5PiBkMCd5xlzg2R4l5ptdtDk+TIoUZzmAmW1VEPB3+kMqDcHCh9cC3ybWyDeVipY/q1J5FpIIJAKJQCKQCCQCiUAikAicKwJpYXGuiGX+RCARSAQSgasSAWJNICqcLl1Ap1Vkzy6Biu6SXrVICRcQ9A8p7VPCzcxuUfzrRWCvF426Mya/Wonn/8lstCYhT02KUq53i0PEQ5LaYgFi3eKE/ZTzvNgux7ygPLtdWm4VUvzt2AAWRSyEWChwe4oWFctdRbm93pHu7fL27w9hDJnsmBJ2A2VBxlYixSDf3mEPcQyZTIKMQ4SgHNxBIXRA2jmmxJKbplOtKsjvg3ZDWDuAN2XwLlghVNythOUE1+BC+bZIsYstBB7euSG6ndFozY1H82A1WsebMXzDxhjaJPdQs+2Y+dq+aJ5gXF9SOpjBtgujcPaXzB/iRmCt9PXBaydjWcjKIjZU496NQ6Xbtw/F1kqpv1aYG8xDYk9g1YKwxJm5QywLxo6gxCTHnuA9dqmzi525gLUT881rgHyMpV21pcudsx/DzHmWCGBZcRrrCr5TWP28ZVlRXgusDdaIY6yckm0F66WzbFFmSwQSgUQgEUgEEoFEIBFIBM4PgRQszg+3fCsRSAQSgUTgKkFgIFSs1b+HJrghub2r+mxcQhXR3asf7HyljVgBUKbiVvT/MxEzj5Ri9tETUlqeU7K7JEhTiHjIckhbiHPOEFSOpeE+Y1VgV092/UQbuTbh6jbbFQ7tW27RYFHGbS/2s3hNXY574bz8Lo4B1xD8tgRhl7pdNCEgmFjGZZLjUBTFCvrKbncCKT+mBJlMWQ6m7TN5ED8I3A1ejtWBqMBhgtnt9+5j8KVexhUimvferoSQYZGH+rz7nvdNhA9rnOoSK+aiNT0SnRlZU7RV7pDcsZSOx8hNCzH//ek49gXteu5MqjSI8b2D9uTp3BAAd8bgaaU/V7JjfyxX+gM1XI57dw7HvbeNxo7raiHNoj/mjCNz4ytKn1dCvGD8WH8ESv+sEgGKGfvvKiEmMh9wGfUJJQKkO2YFVhq0wbFZznX9n1uPM3ci8AME/O8PFl18n95UAKe/BnSwJlgbrBHmac7PnEGJQCKQCCQCiUAikAgkApccgXQJdcmHIBuQCCQCiUAicKkQQKxQ3f3d/nLbtBZEDaQ1BDsEd5/gVz3n1F3trG8pCPe39RLBUokVQQEQ9bfqSoGZVez0Q40YvW1rjNzSjFIF4p48DqJNfXadZIsFSFnHh0Bo8DtcF/3tQ9LadZNdRPXhGvTHnfFvY1h0J+X+WqgwiQzBa3KfM3XZHZXFEs52BwWZxg52frs/tgbhnvvg9ll8+bRuICzg8uTWQf9oA+INZVoo2alrSDxc+jgQ+cn5MegEbYTg433Glec3LOsHdYEz9eNOisMxQ2j3QvS63WjNlqLxYi/ak90Y2jwm64odcgs1H80jR+UKqiy3Xy2hgUuhT6R1xQDF8ztZKGQMvqT0s0oID57EQxOKZXHDcHz6retL7c+d6B1c6PQFvnuUiGXBnGCssZxhvBEjsKBA1GIO7y3MAdx9IZJ5HfWtejKg9vkNXL51wQjwPUWQRYD7gBLfLx/9NaCDNVG0ULvgSrOARCARSAQSgUQgEUgEEoFE4EIRSMHiQhHM9xOBRCARSASuSAQGYkWfWJeIsBYuWvobuClfCcHCQa3PBy8IUtx2QKZ7pzeuajoq/fpoHR2N+d3TUdnwYtS23NwXMpbIfQhyiHMIKdwqcZ9/+y0ecMZaAQsGiHYLArTd7/lvBYsDRcVlJYsL+lsMsF0M/G2LDbcBLCxOLBc7XA95HQ/CwgYEHH7XIeOKlhEOKk655MVK4/sa3y9qvJ/V9S8rERzZwcEZH94nGC19t8sf2rQ8DgdlWngoWp8YH4sm7ofzYJXBNW2el3VFJTrNcRlPdKO3OKpA2wr33BiKhQOLUaoOx8LuiZh/4vBAJmI3P+JUHmeBAK5rVnCJw/zDWoL5gqXSu5UsJHmQ77tuuNS6Z11v4dHZmJdgQX7mD6LW+5UsrrGGmCPsWOc5ljtY53APUcPPcONlN21r8W05CzQyy9WEQGFe97+5Z+mmyTGN+Ja9eQU8ENRYE6wN5vwr5upZ1nM1QZ19SQQSgUQgEUgEEoFEIBG4DBBYKxcYl0HXsgmJQCKQCCQCicDKCBQsK9ZKrKBiiGxIcAjxfnyJc7WucOu1w55d/Q8rQbpDLkGcQqLeINp0Wyzs1U79ozfKvdBO7d6nPruhYXc45KkDYkOek7Ag4KBcfjuYNGWTEDDstqloReHr5dYoy11G2T2TBQrvcufvDlsfIJRQv2Np0B7yF107GQLOFhHIT6wIfuMmCtGBg/dclq1H2PF+m8abcSAWCNYW7ICHqANDCD0CMYMl5DRj5ra6HRYpqAOxiLLAgTHlfccFKbr84h36B7bko58Sl3rtaDf2RevwwWgerUR5uBTlito/pHOtEq0jC1F/4Xic+NazYtLxJ/+Exj6PC0eA8cC11jeU/nR5ccSykFuo19y9rrT53RtL7dFy7Ne9R5SPhEUFMWDw8Y/7J8QuLC8QDxl7r3HWGYmYKdTH2HdkXXHhrc8SEoElBJZbfJ0OFwu7iGmIa1gLrXSwFlgTrA27CkysE4FEIBFIBBKBRCARSAQSgUuOQFpYXPIhyAYkAolAIpAIXCwEBkKFq0OsWAs3UCaWILMh09m52loFK469KudTSri0wTUUFhGjorB6Mfv4UKy7azRGbxXxPTYbIzsgS3FrA5lq0YAA3By0h7ZtGjy3FQbPeA8i1j73IfEdq8JWGRDzdhPlvhaFieWxL5b7wLLwAEGGOALpy+502lS0Thg09xUnW2e8od//JUsIyrBLKOrjHkIBiTxvVCKgNjvgb1OCxEN8QLRwUGyuwdSupKiY9vi3A4Lz2+8UXWM5XgX9AncLQZS7JAyVSmpL75aojJdjeHsp6rv1vlx4VWpzGscjMfvNxXj5D76vGhFVvqjEDv48LhwBxpF5jvBA7AlcrJ2y43yoHO/aXI3qW9bH7m/NxPEXFvvjx7ghVCDg7VXCjQ5ihQUv5i3zysG5Eal4Rl3tFCsufOCyhFcg0P9G2uLCFhArWBbxLbteiW8f7vCWH6wB1gJrgvm6Vv8W5hAmAolAIpAIJAKJQCKQCCQC54xAChbnDFm+kAgkAolAInCFI9AnmddQrAAe74SFvHSw3QuCTTvtO4plwa57CCbiJrB1G8uAjXIJVY6ZJ9oxevtcVKqVqK7bE9VxXB9B1kO6QqTi9uhJ+q5k10mQ7JCuEFYc3GeHOK6I3jn4XQwkTR6LFUWCy4KFxYKiG6iikGABwC6nKBtRwRYgRQuO5deujz5RJv3pW64M2mT3W36P37cr/ajSLypB0N01eJd+2EKC8jggqBEX+NvIcSgQPo4MnhHDgHod34J3LOyQz4KG41zwjB3O1AP+aum82ro4HPW9cto1M6rf7aism4/FF6aj/uKxOPapA6phUghjSfO0xjxJxMHgnO3pNC5seiJ0GR/EBVzg3KHErvOiT/97hyvxQ7eOlv7PN66Lr++v96qLvf46Y57hlot5hsjHgYjBmmHOUCbCG/OEMUfcsMh3ts3OfInAGREYzOuz/R7wPeK7jqj724O5Wiyfb9LnBmuB+dtQ+Wdbdo5UIpAIJAKJQCKQCCQCiUAisOYIpGCx5hBnBYlAIpAIJAKXGoFicG3assZihbsLCd8XK87XFdQKuEGo43bmrUq4MqpKGhmOXlte9x+tx5YPiICt1qL+0m0xdtsjURp6ozoLecW/95CpEPEQ+pCruLd5vRKkLYQsu8e5RkRA7LCFCM0wAcu7RT/nFirsYrIY08KiTdFdlLvkMhAL7CKKM3UWj6I7Kpdj10tul11CWfTwffqMyOA4F/xG7LHwgNhj11GUaWsSx+6AjLbYwj2EHOezOynGAlGCcQZD8KOdvIu4BGm4Ua6gJFA0R6KzuE5unzQGrY5KUt+GqtFpNeXGazRmv70+Fl98eeAK6mGJFRaRlkGSP88HARGyXYkWWBcRD+YTSh9SQsDqHxqMN8kxV2wZijf/ynWl5w81Y983pnuTrV5/nbx2MMZP6YwISTm4XWP8WVde6whT3bSsOJ8RyndWCQHH7mHOvl0Ji6DlB67yWAOshRZrY5XqzmISgUQgEUgEEoFEIBFIBBKBVUEgBYtVgTELSQQSgUQgEbhcEZBY4ab1Ly6SWNEP5q3EruzV3LkKMYrYgHsn0o1iWmdVw1C0pjbHwrPdKI9UYsO7N0fzyPeidv31Uaqw+xthApIVEoszVheIAxDte5SwRGAnOX8X2KWR/0YoCg5FCwqTXEVhoihgLBc5LD44CDUigAl+l9F3paNkV1bLp5UFEQf1Zqcw/SGuAH1BhCjibfdNPKdftBlhZsmd1pJ4Y1GiGL+CMmgbIgWH83KfuhEsIKcpC3wh/hxY21YfuORqS6yoRrdzg8QKiRRzE9HWa+V1qneuHu0ZOSGSB67mwUNx6AHcCu1Tiz4rsYLYI3msPgKOcbJPRf+R0j9WYt73DyaDQqC/bvNQVP/+ztKG6XZvz5NzJ12oMd7MT/z9M2ewpGB+MJ95lfnXS7Fi9QctSzwnBPiO4faObxbf/eUH3yvmPmvA1m3nVEFmTgQSgUQgEUgEEoFEIBFIBNYagQy6vdYIZ/mJQCKQCCQClwyBgljRb8NFEitMzPfjKqyidUUMAjCzOxaXQV9XQrxYEF2qHfy66iyc0E7+WjQOVGPhuRuidRBy6oASJCuWCBBUiAEQ7ez+hxg30e5YCxD1JHaO++8ECwQeS4sCxfsWHchzOpc4dkVFO9ip7jp4F0KYXesIMVhCFAN3WwhZLojQTtrAmf5RPnmKYgpiBc92Kd2vRIwOW1Msd11FWW6XBRUIQPL7HQhqykP04BkiCa5XKNeiCFjeIrHiNdHtbo1ua110FzdF4zBBtiViLA5FSa9WN5SjeWg+XvyXB6I3o3vR0BhDJOaxBggM3N4wRsw/hLo/UGINEJC9f2givnOkHLftqEVVAbjrm4aiot8WCLGiQZwixghrj/nKvF2QUNFSyp3qazBuWeRZIeDvL98wvlW4PcOtnw/mOHOdOc/c7wur6QrqrLDNTIlAIpAIJAKJQCKQCCQCFxmBtLC4yIBndYlAIpAIJAIXD4GCWLCaVg5n04G+26LVFCsKlUKQQj79PSWI+qVd42W5JJr8m7noNI5EaUR7xMcQJtjOX4nhG+zGZovuQbBD4nOPA+Idt0Ym6rEMsGWIrQ98djMci8LChJ/TFgizopBhSxPv5nUMClw1UQ871fl7BCGAPPTJlhIWKIqY28qCZ7xHP3nPh2NaWDjyfdpYDOxdFDWK/UJ4cMBuB8/GIoV2I2IgsnCNZQdCEHhBBO4d3L9z0JdRCRaV6HUqilWhns72ZFnRk1ixFCi8NTUVPYlLh/5sNuaff1E9of8fK3Y0r9cEAeaNLWQY53+udO+ymj46XI6f+9XrS4s/sqlU+c5cb+rPD/W6exb7Qhjrj/ndXyMDi4oUKtZkqLLQlRBYIcB23zhIiTPzEkH6o8veRQT+jBLf+77IxvxNhBOBRCARSAQSgUQgEUgEEoHLEYEULC7HUck2JQKJQCKQCFxxCCwTR9aMCMLKQsG32SELIfURJXbSsitfFhWTSkeJkaAICTUEgXEFcx6L6sZWlEc3yMQEwh7CHcGCNkKeI2JAckFkYXXBLnJbLVhAYDyWWzlYGPBYWahwUG6TupTHDnVIXeog9gaihMumLZD1fYsUJQQDCDVbOLi8olBBnUXrD8rjud3zWDApWlsUrUpPNz7OTzlgQZtItBuXP5B81MPOeuPIGSzIB5a4GKIfS/ExOnObozvVjG5DsSqaZVlVtGL28a7G5KU4/lfb4+gXHhPViCXMpwdl0rc81h/cWKsAACAASURBVAgBdpSL8MW1E2uGcWVNvGeF6lhbn985Eht3jpQWZWUx+zu7eyctctKaYo0GKIs9HwT4JvG94nuO8MzcXX5s1A3i6vBtY+7X07rifKDOdxKBRCARSAQSgUQgEUgELgYCKVhcDJSzjkQgEUgEEoFEYBURGIgWkOYQUJDsN4tGH1eshMmYe+KQYlfcHJs/WFP4X1kI9DZH/WApRm6ZkbFFS6IF72HBALEOYYt7I8h4EmKBLRMQFPx3gu/5DBlf3FXOtQMP01N+Q4zZ/Q67e3GhQ8Bru1dy/IjlVhm8B7nG2aIKZTr+wHL3VEaWOu0iqhh3w/FEitYay11L2VKENoEHJDaiiQOB2woEPHCxhcXF9YN2QhAiDv3CoL+Q4WPRbh6K7vTmKHWbEi3mZGkxEu1pBUTf04j6vk6c+JNuHP30Hkkajyn/k0rfH7j8cn/yvHYIMN7MR+Y4gtnTSj8xGG/P+Zv0+11KCGbf+8Dm0pyS51UvXmIKLB0ifteupVlyIjBAYAXLCmPDN45vN0Hk+eYyd33wDWNOM8efUUJ0RUReM1E9BywRSAQSgUQgEUgEEoFEIBG4UARSsLhQBPP9RCARSAQSgUTgEiAgchui/BOytvjxPkFV6sd9uE3uhypx/DONGNt1OCrVTky8eTzaxw/H9IFWbHy7xIKh55R3k/IiWODOCJIfgQBiFuILwt5unOzqiWc+fM9CACQ/z7mPGEIgYlwkYVVh6wieUa5jANwyKIxdwRBoPENEgQVGhCE/1grcdxtdFq8ud1FlAaVoEWKLDPt2tyhhsaIYcJsync9lkw9BB8IPkQUBBeGCNoEf7aU+sIOxRvBRgG0F2e51W3IWtCE6k/VozcsCozMevXY5Fp4/Ecc/3Ynpr9ejcbShGhkLSMRHNJ4QjXlcPAQQpJhjzMHPKb1JiSDF1w2agOXS/6KEmPR/K7HeLGJdvFZmTYnAmRHg/8sxhxFQf1npnsG89ltYbyFWMMfJh6DKPM4jEUgEEoFEIBFIBBKBRCARuGwRSMHish2abFgikAgkAolAInBWCHxHuW5XeoPI7y/rLNFi4Ugc+2xVZ4kVM+UY2bU5Ru/cFM0jR2JoWzcqNbtggoR1HAhIeZP8kO9YGSAgsAMdUaNIqEPm28WSLS0oB3dPLykRFPwLSk8ovV/pw0om/HkPwh+CjTqoCwIN8p8z7UAU4F0INp4jDiBcnMkygnKLMSr082R+Xxd3FRcFiqL1ha1IaIOFGp7bAgUcqIfkYynYd69XV5BtIhtU+tYU7TkJGI2Z6LUOxuILI3H048dj8qHJ6C0sCD2IRAKnPyyxgrLzuEgIFNxC7VWViGy4hGKuM3ctWOzSNWmn0iNKCBicCbpdjJkS7HxPK4uLNHjXaDWnsa7gu8y3/y1KWFj8lBLfyeLBnGZu85xvKqJxM91BXaMTKbudCCQCiUAikAgkAonAFYJAChZXyEBlMxOBRCARSAQSgZUQENl9UFYWWCUQOJjdtaMiwzfE7Hd7EizmY3RXJ9aLz5p/fibW3VWOsTdsjtqmiRjaCGGOEHCbEqQtJOxSQOglMh4SHrGCAysInhUJf1ss8NwCBtYVlEOw6lsHZ0j/P1R6uxLEGnkh0IjD8YZBXeThPqQa19SN+6hvDe5B6BPkGnLO9XG26MA177icousq5/e95a6hBkWeFDfIt2Qt8YPYGsSpQJgBD4s5YERflzDpCaNuuxvtEyOKI9KLxWf1TlUixkIv5p6ajskvHY/ZR5VnESzH1HL6/80UKwz/xT0PCNuGiGDWwcOD+cMcfetgTJ/XmQDqiBSMP2IaYgZzFwuiU0SLi9v6rC0R6IvIBNdmTjI3+R4xVxEtnlNCYONb9kUlhFG+pcc07+1aLyFMBBKBRCARSAQSgUQgEUgELlsEUrC4bIcmG5YIJAKJQCKQCJw1At9WTohzheTuE1iHRN1fH/N7ZqI9pX/ru7fG+vsa0do8Es0N90TzxcmYuG82quuxejishBCAqxBbWGBdgI9/XCKZ4IesL7pLWu5aicZCoHF/rxKuqh5SglizmxJbV2BhsXlQB4IJeRAkeBfiDXdSuKyiToQSfjuwLO6XuO+2Uq/bsrx9PMMiYikA9g/ab/GC5z6K92gPZSIucI2Qwhni2gd1uT5ZUfTmZM2CWDETjf21mH/2UMw8KguR9kKc+NyeaC5MqAVzajU7oMH8CxIrEJryuIQIQOBKtECA+N5gzP+Nzm9TQqzguE+JOflvlbAcYn0xp3inGMflEvYiq77GEOB7xveTucg85Pv9t5XuHuDA3MUS6JtKiHG4nTuaYsU1Nkuyu4lAIpAIJAKJQCKQCFzBCKRgcQUPXjY9EUgEEoFEIBEAARHfR2Rl8SVdIjr8LSV88y+IIJ+O1mQvph/eHtNf68b6t03Gtp+dj8qWksSKbTH6+g1Rqg5HuXxUwbgh6InRgFsnCFn+RiBB5CNssIsXocCuoYoEfzEoN+9jOcE9iDMCwHIN4W//6ZSDFQZnCDfqoXzECAQKWy+8bvAcNyavHbxj4cHumlw37XIcjmK8Cruu8s5i2gHRvNzSwu8gSrhMLFDcdiwruEbE4aCuuoSKstxAlaIlF1AzXzkUs9rkvLhnLI5/rqPYIaqlSz9b6iFnBAr6/DGNGbuhz+vo9XoarqUmcq3jlMDiepYBdc8NWcZ2vxJnxvVBpd9RulkJ12Wk9yn9e6XPK0EW2/LCweHPrcbMnQicOwIser6NfCMRgYkFhEj9i4N56xJf1MU/U+K7iRsovrHpdu7c8c43EoFEIBFIBBKBRCARSAQuEQIr7TC8RE3JahOBRCARSAQSgUTgQhCQaAGRhdulDylhxSBCvU/OD4lq70pqINDz+tj20xMi0m+MjR9ox9afOh7DN4/H0KjI+dKimHAEBqwAcBOFCADRj0UAu8sRQyB0HQC7KFSYJLflA9YJuNshGPhepRuUINuw3MBdCcGqyYOLHUQOxBKecSC4UD8HZ0h+CDoEjWJcCYSOovBAfvoLiQwWlE+cDt7BgsOufN48+E29uPbhHbuioo0WRWydYUGAvCb+qHdRtR+Nue924qWPzsXUF0rRoLsliRULHWFdVkL0oG7K/Bulryo9JMHivFyzFAQKcKbdxdgdS7E0dN+iRVHcAJw8VkZAVhbgiJjFeLFz/TeU/uEgN2O+VwnLo8eVPq1EvBjm2SHOGRMgZ9ZaIqD5abGCuck3irgrP6NEsHjm567B/KQZ/0LpY4O5ybenpfmZ1kBrOUBZdiKQCCQCiUAikAgkAonAqiKQFharCmcWlggkAolAIpAIXFIEsA54Ugmx4qeV5kWY46aJ+3VR5m8Rnb0YRx7AmuFozHxLroymb4mJtxyK9e+cjtoWW1cgHsC8IxxAeBHY+wEl/KD/shKiiINOW6gwuQ+xBrGPuGBLBv7ewK0TO36pA2KdeBckx66gPEQM8lInebjH7nbEDohkyoVYtjsmixfUbZGC9yDw+E2/EUEeUwIXykCQcSwKW31wn+vlbqP8HKsK9wsrEdp8MDpzJ2LP/9SM/f9qMZrTG5WjpkQbO2ol/ef4rhI79ek/vuQvVKwAH7vqoo9g5N/gQJ87EiosHJV03bNFxqBNeXolArawsQUNogRY36/0w0pY+HDsUmLeMg+fVkJQY84Vg9InvonAaiPAfEOE5fv1eiXirXx4WSW4f3pUibnLwVxGEE6Lq9UejSwvEUgEEoFEIBFIBBKBRGBNEUjBYk3hzcITgUQgEUgEEoGLh4B27YesLLAo+IIScRcQB4gFwa7cpYDWJRHzFV33RMY2jo3F9CO75VeoGcM3vCZK5WZUJ45HuQopz85xgrfaigKS/z8oQZixqxcyn2dOjvtAh9mJjqgAwYbYQBsgdh3MGnKXhCUHz4pBjXHNQ7sh4hE4cL+DkIDIwpmybVVhkthtsYUBRD4Hv3kGkYdw8HeVcFeFeybqJp/iTPTJZ9oHucd9iD4LMpSDpYhxoH1TMf2t52Lf/3pdHP/rsejMH1DLECpw0UK/LdCQ96ASAgz1f+0CLCtoI32nXVzTd3CwhQV9oV+0nfFbEk5+kJK0ZCRPf4APGGKFwzX4/YUS8wGBjnnk49d18fNK/1KJsX5SO+CZP920tDgzyPn09AhoDq30kO8Oa5zvN1ZmP6r0W0qI0sWD+frSYM7yzUF05rvlb2FCnwgkAolAIpAIJAKJQCKQCFwxCKRgccUMVTY0EUgEEoFEIBF4dQQQLXRA7v+pxAvILQQBSG7+zYdMRzQ4JPr9OqXhmH389dE81Ijyul5smG/FmMJO1LaL7CrvkHuom5UIRgxpdq8SggGBXCkPSwvIccqHGHcAaltaQPraZRNEO1YMJoIh10ykQa45wDZts4BAeexqh+xH0KAMRBN+Uy5tsVUExBwWDbxvKwPECgQPLBt+U2mnEowg5fMe+SjPlhx2CwU5CH7kRXDht9vwTHQWj8WxT+2OF/6HbTH3/Rv7rraWAjNz0C8Srqjor3fr4wbqrzU23D/nQwYS3l1tKxPKoG0WcBgPRAqek5c+uz/9QOGDMoh9ka5hzjwCS+tjiRBmbjgI965lr/GceYtIxdzDgueESOeFDG58zlP8mn/hNGIF3zm+UYi2iBWec8vFCvDDIo65imiBeMa3L61+rvmZlQAkAolAIpAIJAKJQCJwZSKQgsWVOW7Z6kQgEUgEEoFE4GwQQFzggOxybArIfXbfIkNskFgxEZ3p0Zh/bC5Grr8jeo1uNLfOxZA8MdW2tWRtsU75cKsE4X+jEmU+o4S1BSIGgbFx22TRwsGv+7EU+rUsnSHy+bsDQh0iHwGCZxDvdm0Euc5v7kPG845FCVtRWNCwNQVEPWQdZ/plF0mQzryP+xTawvu2qnC8AvI6CDckIBYK9hVvsYN3IQ2nYmHvd+OpXzwiqxRcPN2hnJuUeIaLIHCFvLYlCKIBYgzuqB6WWLHi9mk9O+MxcO3kuCG0z8HQwRkMITPBAtdfFmJcpt1j8Zs+4x7Klhm4iUrxYmX0wQhxCUsfcN2ntGuQFUED3JlzjMd/pkQAbsZhD3lFPmdci1eb2Pn8TAgU41XwTblV6S4lLH2YW8w9vsWei5TFHGWu8m3lu5NiRc6xRCARSAQSgUQgEUgEEoErFoEULK7YocuGJwKJQCKQCCQCZ0ZAJPm0rCy+MiC43quziXtcRCFEjEZXt9oLCzH9jZeisvm62P7hsajv2Rbl0amoT74Yo3eUolRjJzkuSSDnIcTYyf9RJQgzSHJ2mHPfBBpEuQNV00gTcHarVIx3YZdSjs2AiOBg0hDDdutE27lGEKBOXF9RHy58CArOGWKPPDwjDzE4LE7QPsqlfN7jjOUE9+ibg2/bQoPnlHNILp+ej8d+6UDMPDgR3cX3qjfEBgFD2k57HH+DuhB3IBlfVHpAY/A1nc/rKATYpu+IFhDkjo2BQEO9jIXxRmQBM/pKn0xacqatFpNoz6LKRyhCuEh3Ua8cIQSL55XYrQ5BzM71vzPAl9zg/p8OXpNZUjyk9GABY9yBpTue85r51/xLfLsQJBCCmVvvU3q3EkIph8VP1jrHnylhXUGsIb6DfN/ySAQSgUQgEUgEEoFEIBFIBK5YBFKwuGKHLhueCCQCiUAikAi8OgIizBclWnxfOdl1+3NKEGBYE2CNsCAaGyJ7LBb3bogT/7EVG95Sjsq6Rkw+OBIT9707yi93Y2jzk1EaVSDp2tAgiDcWFuz2XYrnsETSQ6Tb7RNkut0p0UhbWliw4B4kuWNa2GUVgoj/NnFex5LA+sL5EQn4za5iDupDIKAdkHo8h7R/zeAZeSCPKRsy0MnWHQ7QbcGFchAHTsTCc0/Gd3/tREx+9b2SPsbVf/oI8U8ZkNn2HU/9bxvce1znP1EiKPOFHLY0od0IELTTO/sRkcAVSw6ITTCwhQqYYfEBoYmwwn27qrKFC2XSfgJ09wNOI1xwmQG6Tw4Z84G5QLB0xAuEsd9WYlzs7ovMzDnEC/IjmrHeHpClxWTGtLiQ6X9Nvsvc4tvzTiVc4rG2LYwZEM891u3vKf2+ki3nUiS7JqdNdjoRSAQSgUQgEUgEEoGrC4EULK6u8czeJAKJQCKQCCQCr0BAogUEO7vv/1jixQ/p/DNKWB9gZQHpzfWxmH++FYf+eE+s/5FNMXH3cHQXDkTz+LpondgVwzfPR2V0Jsoj1ShVRKqV3q13KZN0QIly2PmLGOLA0A4ObSsKt82/7RaK35BvvIe1AAfkL/fIA9lul0/2z85zrA4QXmgDv2kD7+A2CtIPop6/dSiD5xB9ttQAE8okIZRARvPOl/vt6La/HzPfPhTf+7XxmH36HtWEUIHrJ/La/RXXiB62fKAsyvm0MCfI9oUeFiyom3rY9Q8xSR8gMjnssx7swMMWJBZ1cNtFexGZIDPBl7Jwj8U1GFFPcyBc9N1GXWuihYSFPpgrxBJg7jHnOP5IiblE8HYEQAQxH+xuxyUPAhLzAhdqbZXH/OylcFFAKi9XQsDfRL4lzB3mEGuZOcXcYh372KsL1v8fD+Yk34R+0PeENhFIBBKBRCARSAQSgUQgEbgaEEjB4moYxexDIpAIJAKJQCJwlgiISP+GRAvI6rcqQVZvVIJUfUwWBBNx4qFSNMR/tQ+Nx8T9YzF683RUt3SjfXxrtLqVKJVnY3jnO+QySsRsGcEDMhy/6hBskGgQ5Y5XQatsKWFCzqSa7zvWBWe7LYKYRxxAeMCCg79XIOUg2LnP89sG7aYO4mjwLhYfX1L6qcG7dpni2BkQ+tTvv38QGGgvdSC6cI34MR4v/8FcfO+3tqjUuwdiBTvscdMCXtRPXsrfrQRJ3bdWUPp9YUwZq3FYsKAs+k37ES84gxcCDInfiBD0C8GEdkB2IkR5fMnvuBe2hMFKBEwRmegPLrL67qEkWlj8uaYsLixcFAavj5uEB+Y0AhxCFLva2f1eFCwglElYHjEX/sEAb9bGgt5nrZ3W9dYK9RaakJdXEwIriGKsc9Yv31Asooid8g+VsKqyMFmE4Nv6gRUPc4s52dL8yZgVV9Mkyb4kAolAIpAIJAKJQCJwjSOQgsU1PgGy+4lAIpAIJALXHgIi1D8l0WKven63EjvFIfzfLnJ+REz1jph/RoR8e2/UbqjFuntr0Z6aiNZkR66hNsnCYlM0j1bkNuq6GNqkfGW5Qip19C5EOYQs5DcEOiIAZDmEWlEkKAoVkLg8Z+c/9xEA+NvEbpe4Jo/JOHYbQ+xB5EHg4xaJuogTgQsVhBiCi1M3hD1CAm1wfAq3C0LZBL5dS/XkFmsujn92Zxz55L6Y/Oz9atnYwAKFPOx85p0+AT1oL9eIEzz/G+H61zqvyjGIX0F7ORBWuEbAof92/wRmEJz0j34iQCC84JYILHhOX8EXrHjf7mQQJ+gH93i25BpsqS8IWA5qflK4WJWOXbmFgAlWKoz5HUoIVR8ajEexVxDMpJ9UspXLt3RNsHoskHIX/JU7B8675SuIFC6L7x/mPbiTQ0RmfbMm+SavdLA+/0oJAZXEt85WaefdvnwxEUgEEoFEIBFIBBKBRCARuJwQSMHichqNbEsikAgkAolAInCREBC5/qREC0QGyFVIsDcqyd2T7nW7jZjf3YoDv79BQabrMXanYleICy+Pj0vQaEZrqhdjd/SifawdzdlqVMbGY+SGab17RM83a0s+7pdIEGmID/57g7ODaBddOvk+pDyWFIgD5IOItxUARJ7dOSFGcM17kOxvVsL6ASEDUQMyHiLQ4ohjXyBgINBA4C/5eu+2JqM13YjF5+fi4B9ui6OfXojW4V3qx3a9DfnPu+x4RpigPRYNntU18Q0gsRErIA9X86D9JPrqINr0lTaBDXETwAuRh7oRKewKa/OgzcTVwJ0MhKhjgdBG3kfQgDxHYELs4KAsCxzgQ/l9F1GFjhHrYjX7eaWUxXxj/BEhGHfwI57F+5RwscbY+EDcQDj7W0pPDq7BmKDc4GtXad3cGX+lDP+FtbPgcow1xfjb2otvFnOIhOh6j9J/UGIO8R30gbj46cEcQvhiDtqa7cIal28nAolAIpAIJAKJQCKQCCQClxkCKVhcZgOSzUkEEoFEIBFIBC4WAiLZj0i0wFKB3eLvUnq/0nbRaTdErzMT9QPdePGfN2Pz+2di7HVvkFDRiZr0gPHXTsjKohyl6sZY3DMclRERZx0R/L29Ud2+Lyo1kbNlCLkDIv0RRCDCES7scggRApEEIh1SDuEE8pz7/G0CIw6RDjFn91Im+rAoYFcxpDzvkiCPedekseM0UI4DfkPu0VeIQMXn6A3F4jPzsbD71ph9/FAc/ctuLHx3Itp13Fw1lSifdyHracs+JUhDiH/KIiEGPKCEyLLah11lOUA4VhXUTZ9w9UQCQ+pGqID4tNUE4wl2e5V47y4lhBfyY03x+sH7BAWnPN53nBP6YZEJ7DnAnvf53Q/SfY2KFmABnrge48wYIGSB/Y8P7iEugdWuAXYQ0IhpTyhBSL+gxDgxPkME5h5gD/7pMmoA2tV00hjbtRvriG8J64hvH+sM13Z8a35pcKbrzB3mEN825hlz6iGljyt9TwnhlXXv9Xk1wZV9SQQSgUQgEUgEEoFEIBFIBE7ueEwoEoFEIBFIBBKBROAaRECiBeT+nISLzw3IsXfofINo7E2iT/dHp3lzHPns/hj9zmtiZOeJGBP3Xd2MWFGRqFGSayiRbt1uNI+M6J17JGDsV4DuI1HZMKQg3evkQmpRFhczegZBC/FmsQLyDgHgqBLEHNcQ6tznHhYVJIhcx26AoCMf+R2M2zuVObtMB6i2AII7Ho5tanNdQcS3R+NAJRaem4jF5+qx55+21M+NEmqqSrxL2Vhi0GYHUsYNEPeJYYBbIIjnTwk/yMO1OGxNAnHJgRhD/40F9yEzaRN4QIqCG23mTDBuBBfIUEhSzjcoQZJyRvzgDJ6IGMwDxgcSHisA+oWFBgIPmJD/pEuja1i0AFOwZ34gNiCwEaj9OSViWLxHCesU8CeeBQfY/67SXwzwtqUOeNqtmV2L2QXXacWLQZl5uowRGIgUrEmsKVg/rEF/yxhzrhFfEYl/YTBH3CPmDiIXB98uhFHmG3MMayrWfboWu4zHP5uWCCQCiUAikAgkAolAInBhCKSFxYXhl28nAolAIpAIJAJXBQIi3iHAvijhApdDLyv9hCjw40o7dX2LrC32ieSXXcEzG+Q2aXdseMdobPvJ66Iy3o3qpmq0ZbxQ3SAitrQ15r8zGjUZVtS2KUj3+HB0pk8o/sVBxbyAuJV7qTLWCRDvEHYkyFnEBYg4EgcEPW2CKOfvFcfBIJ/jMFCGd6ZztqsnCGF2sdtd0o3RqY9H4+iJaO4bjfpLnTj+mRNx/IF6NE701Mftag3vQixCMNJ/yqa9lIFAQTsfVcJK498IL4LertkxsGDoShhAUOBgRzaWEJCgCDt2DYUAgdiAixiek48DocUWKJTBOEKU4qIIixbil2A14ngf9B+cIePpLxjzvrEGU/A5GQ8E0UK/+8TpNWhxQb/BlXnAXMGKhVgqewZYL48rgDj0E0pfHWB+v84Q0BbyHJsETBGMEIoyfgiT6wo6BkIF3xDWDpY3rFfWEG7l+LaxPu9U4luCiMGcYG4UD+YOlhSIyMTF4ZvHb+aavwdXECrZ1EQgEUgEEoFEIBFIBBKBRODcEEjB4tzwytyJQCKQCCQCicBVjYCI+GclWuDyBkLtdiV8779eNP6zkhUUt2J6aRf+8U/W48SnZ2LdfRti4k3dqEwMyVXU9TFy86isL4aiM1uP+vyw4l5IsFgciebhHbLQmJZFxtHotWckXojKq+0WnfeW6HUJkLFkLbBkiYFIMK84EuvFhIO3yXSuIYcRPBAyIHS5RqyAuFfZnUp05majPVOTwCLXTrV7YkHxKWYfXx8NbVxuHh6K5svdWNx9k0SMivrF+5DD9BPCH0GCfrPLmTgVXFMP5OGfK+0RRhdz9zsCAdiAC2BwbZcyYOAYH+y8hiS1FQVYcQ1ejCf9JC9iBHjiFgrCFEsK+g8RinUF7rXYzQ1pCq4OhI6QAdnK3460BQxIlO8A3dR5rR3ghtUNmLxpgMlTOkNaLz8grX9aCZGI8SjOX+afrYd4jvCB6Dar+Afp+ucKmFUSK1hffIdIxJRhTFlbiK98W1grnIk/g8DFc+bE8gNBkTXIemOOfEOJ7xFCZR6JQCKQCCQCiUAikAgkAonAVY/ANRk18aof1exgIpAIJAKJQCKwCghIuIAQv0/pZ5UceBmC7U5R1biwKevupqhW6zG0tRLVkfUx9oZybHqv8pSHotdoRmV9KUqVhRh7zeZoT85F7cZSdOvTMXyD7g81lWdrlIYbfYuM6Ci2xEJLIoOECwkb0d0WlZII87IsHso7RNdD4GL18JKEiUZ021tUZk/nJRdRM984FOOvvzXmnxR5rBga88+0ozM/ElMPtmP2iTEJFHNqd03l1JWWXCxxvUS8QzjTJ8qHMOQ+4gW75iEPH+F8kcUKaTZ9bcRBehEPLJYwDpCfiAwIBrSRQM+Qovi3Jx8uiSBFIce9uxsynfcIVE65iDKIECQEDHzqQ5iTj75DolMX96ifd7EAgET//9u7tx7LrqsKwLuv6djGcexwEQKlcMgVB6xAQEASDJEAJcIgIRAPPCBEfgUSD0jwJ4J44gGRByBgcxOXBAMJOI65xBgnikuAk8iAHYc23V1dVc38Tq3Z2q50t7vTdbpP1RnLmtrn7LMva4+51nb1GGvOScQwLlx7q6IsbqWQU7e89a1I6SvdFI6EPCvnYQ4vItGvlBG8NN+NLX97i6bQfqNMlEXXRSEeIb3/oawFD4Q33/JDalzcepcv7ngVv3dv+NT7xEusC2UTGt5dZp6Yo+YNodAY+aVxIgGCT71nzF1N/ZlfHd+9h7x3jJFrpoHqlPBypgAAGvdJREFUot63CZ7cNggEgSAQBIJAEAgCQSAIHCgCESwOFM5cLAgEgSAQBILA0UOghAsknBQ2VgZbOWzbJNz/1BpgBO0TewW2j1fu9d3T0+l7T0ynv/GOKm59Zto9+8Xp5Nc/O9355m+rVFLfUHUwivjeLlHi9KXp1H070/nNi9OZN9a+YyVCnK+IjLMvVgTEy9M97/3mqoNRxN/Jz03HT99f4sPpEihK5Ni9uwSSM9PFF3emi/9VosPJ11RB8K3p/DMlkNx71/TljxWJvnt8OvuZS9PWFyoq5Cu7JXAopI0cRMzbeqYWKhDFyEHNs4lC+ETZp8seKZECQX9b2xAuiBGdIqujHUREIMsx6fyA8FTDgn+ksbLPMxEtHCMfvlQ1anIgWYkbriuFFHLVtZzn81+WIVP5HOGKYJV6ColOqPAbEnYRBVKCxf40SLV7PdpIBQQ7AlHPDULfzw/c3nYFJPjjowNHxHRHXIiucB1Yd7F1/uNXGH9VqqgQ1ssdZ1cQLLo+hfeJudOChDFgThL4et4QnwhZBKuHyzpt27zTT9cXQtZvlf1BGX97L7nO+fLvkRcDl+vBXD0IBIEgEASCQBAIAkHgMCEQweIweSt9DQJBIAgEgSBwGxEo4QKRjZh7Z9mPliFVkftW5X+p6H9phqzCR4CXsLD4T5qnF6bjx85VuMDF6a63vXa67+G7phN33F8iRdW6uO+l6exTr5nuevvxafvcuWmr+PNT9+5Mp+4pEeKF7emOt95dhbEvVWqpKvJ98Y7p0tZ2iQ+7JXIcKwGjKPTnjk0Xny8S15802yens09emC789/GxFv14rVNHFm7PxApEoD7a39EVSOBOtaQ2BBJZgeQXS6w4V8891fa2txIt9LkNMYq4RnIiTH32G394ljeWESas2H9LmfoV/1hmtTbyU7qo7y+TvkYBceKFz13TYqM+E2oIEn5zjs9ShRFFup4F0t39iBgX1rCWRT32XttXaJl/iHyEIb75UBl/sC6oTBDqwud8A//fH1gT1GBqYKs74hzjtAuqiwbq+i1TBIvLbljKh5lgwR/eb6KR1IUx94gW6t54L7YY2r77ydonMuy7yswj75cfHp10jjnGPlxm/krtZo51RMUi9Vr8uxS35qJBIAgEgSAQBIJAEAgCK4pAalisqGPSrSAQBIJAEAgCN4JAkdnFFS83JU+R9sjwaRTmLhp/en8ZQhYZfqaoVcQ3co5wgWrtdEJ3lVjx4kI0+N+nNypVU0VbPPjsdOL0mYqW+Lrp5BvOTS9XGYCTrzs1vfT42Tru9HTmW+6c7nzg9dP22Sr9/ej2dOp1xyqqYmva3Sox4uzJEisuTV/+1Pb0f8/u1vHSUVUUxfbZSg9FIDld1B9yvYtCI3oRyAje/UWkEZBWsuur/qtH0OmTtupZXWdVih/rRwsTnc++a0gQJrpOhWfhBwIT3/iuwDZiFMnaufRFXyDG/70MkaoQt30EHeQqktw1RWU8WdYpb1wPlsQrx3aNke0ahzvrKlqMVfCLMVcEN9xgJrXWRhkSWlookRa/UCbNk/n0fWUEIJEY/i63z5gkLFmRT3hqkQ05TgThq78uswK/a7gsip+nLQ2BTsvWadjeW3ciNhEmiEjmwXvKzDPzo8WLn67PXUTb3HuijO/NpT8rE1khHZQ5tjmO5dNEVCzNlblwEAgCQSAIBIEgEASCwKojEMFi1T2U/gWBIBAEgkAQuA4Eli1WzLswizqwGpyAoZAwkk29CwQr8g2hTcxA3lW9isV2u4SEl4qKu3v6ypMv1+eKfDhRYsHO3UXDv6FMbYmTC8Hh5Jmd6fnf3Zq2d3YW645PFa9+4p7TlV6q6lKUiLG7jXQnVaD2qpbGeYStcxF9nZpIn5pU1x/EOoIe2a/+AuIXsY9Ilmrpj8a5BAwk5Ll61q7dcR1eWO4hLQSUKOAZ9WsvemQvrVPn0fccfhcpgTyFgd88q1Q0iFZREVbtI027zoV9cCBSECvgaRU/fGydK9WN1FlIWse7B0zds1eer4q4U126fY14MUQLApmxb07wi0gKeMKLL2At6qL/JheJYeW9fbDnDz4yJvlSmqGOrJHqayFa1L2IbF0o/avI7qzQv/ZYuEqNih7TfMOPLVbAnxhIQPKeIPKZG3zlN5EyPzC+u7Hz+ZOv+dx1jQFjwVySWs0Y8U7qqK9rdzi/BoEgEASCQBAIAkEgCASBI4xABIsj7Nw8WhAIAkEgCBxtBEZdg6VHVlwJxXmKpPr8iLRJ1awmR16/vUwKFM3qYUQcUg/J9/xCvjhRKVUuTc9WeqdvrW+vL+r9/CgzXJEStVp55/yJRWHsPQniXEVabE0Xz+7UN8QhYWNPoCA+EDn2WhP5i/xQ47t7I3p9tx8xqKjxXtHwPSIf2ajvVq0TMxYk8CqkgRrP9YoNcWqIFp4XwUm8kKKp63PwgYbwJumInGiydS8aZi9NlPM8r8+iLxTZhlcLTYhzuBE2FAvuFf1qVrRIYWV5R37oz/Hq20K0WNdIi5mz4Gu8SfND6BExwX69DHEtrZpGeOgG164TA3+iENw7hZlIGlEavjfBzW/8byy4V6c3yyr9GbA38NF7As7miblga54QIXw25s0ZYgORwj5zRASFyAr7zLt5ax+bf39a5l3Db8QKZq5eTvF1A33NoUEgCASBIBAEgkAQCAJB4MghkBoWR86leaAgEASCQBBYFwSkgapnXSliuOs91NZqYuluEKnECgKG/vqMPO8c7epgIMURg/9W5jtST+Fix3T9BAQiQt4+BCHSnCESHdNRFfb1Kn/HiwRo0UKaHSuiP1KGCPbbCx1FUX0+XZ9FDByqVuMAOdr4ILy7ODecEKGI1sZIhAmBBhZWeL+v7K1lUmE9WvZQ2bvKkLHtDwQ5IvyZMpEWPtu6J7xEeIgA6ILQCx/cyqifVXbYqG1BYDAe+UH9A6vzv7NMRNIPlUknpMHSGEeKSx2EBFeE25g2ZtW9cJ6xa+zDf7NMKinjXMohq/n/o4xYov5BhIsB7rU2sxokfAR3Ip65wBfE1o0y88s7zfgXNaMehXcW/xKa4E684Avzz7tMe6zsY2WinpznPUQ03Ys8u0bauUTHDASzCQJBIAgEgSAQBIJAEFgbBCJYrI2r86BBIAgEgSBwlBC4ndEVN4pjCQHEB6QcIp2IgdiTtx8ZaMX5RpmoDCQf8g852ylUEHq+I//83dICBFIckYgEtjLZ9ZGGoimaXEfK/2sZkvBLq5Te6UYxvNbxQ7jqv+maFG9Rh2ABY0QrPyBe4Y8sVbPDym/7CBRqLsDU8UQKxDq8HSsShf8UWIe1Vf/2Ow/B3imLmkRf21oWV/LVSDnER/yC7Da+4WwLx18rU9odth0x9Pj4TOAT4aL9Thl/ESrMF/PA+OYPohMfEkDUJUGMEzkWYl6Ei4Hgvs0QKuyFu/cPQci8IDA8WCZCydwhLhHpzBHziUj0s+Ny3jUdySWFl9a+FH/2y2XmExFERIVtF6xPUe0ruyZ7g0AQCAJBIAgEgSAQBNYUgQgWa+r4PHYQCAJBIAgcTgRaqBi9X6noildDtKMv+rj6rmitFf8a4g9JjhhkViAjdIkRiHIrz6WXanECUY6olTaHQIEw3Cz74qqmcno1fG7m9zEu+hJIVYRqY9XpoBCm8Pb3H3IV6S3ipVPetKABU1EY0t6IskCG8xUyF9luFfnHYV3WK8mt4veZES0WaaKSFmrPJbMaCbBv4YKPpA9S8wDWiPJ3l4l6uVoz1kUjIcM3ywhJhAr+gvmny5DhxCiEOF8i1i+n7SrhIgW693xC4OQLW0YI4g9jnDBHTFKXx28EOcKFebBRRtxoX9THKzZzRPo5wpHoJOIhf5h3XatiEf2SKIqrQZj9QSAIBIEgEASCQBAIAuuIQGpYrKPX88xBIAgEgSBwmBFogu3QkcFzIWGIF1+obad/QrwiBYkTD5QhBv++zApx0RgECQIGsvy5uhYSPW0gMBcGSrzo+h3+ziNetICBqEZiEyi0LvSLSCUASYNjZbkV5EQHpLeV+vaLykDQEjD4hD9cj8iB2LWvUxl1bQ33CDn+ylEKGwZfeNkSkohLsH26jOgjhRCh6RfLuiizufLnZQQLvkV8i7xAsLvORpkogC4kT1DiJ8Q5n/PFc0XUO7brJTRhfqTTRs2iKFow8p6R2olA0fVBCEXwlNKJOEpIMvY3y95URtwTDdP/fuILuBJTpZHyfvrNMmKgFF+iYRS3h7v3lnNFxPQYqI9pQSAIBIEgEASCQBAIAkEgCOxHIIJFxkQQCAJBIAgEgUOCwFhF36uCD0mvr9rNYyVWIA+RpwoS/10Z8ptoYZU4Av3zJUwg1W+o7Y9CGSe30OPrgkQ/qjUWRlHurumBHEVs+05YgIPV+AQhhCxxAmHub0Kf/c4fvUIfwUrkQH5bqW/1PrLX+YSQLvZNsOAzJLuWAsIDiKtsmrTmm65n0Pj77T/LCBPEB2S3eiNEI2R4t4564U+pz/iT4GR8i1YiAkq1xrcdzaHYM18aD4QRPnu+CP3uzxXJ9FWPAJhFsMzhbnGit3ASYdSp5AgTip931MMH6jNMWb8vHA9XOLbI0ffgCxEUaoyo0WM+EPgIe64p8oVf4HzNOhXzTudzEAgCQSAIBIEgEASCQBBYdwSSEmrdR0CePwgEgSAQBA4FAoOER5j5fzdS8UjUCBiixaWOvhB54Rnr+w2v+IaRSINR02Ge7gWB20WPXR9JLELlSK/+n9c5GYW5ka/MSv2NMfCRsbAmUiC1pcD5mzIkKzECoW0FuXOkzOnV/gp1i3xBzLqm/Y5F2hIrRA8ciTE6cFrqZlaY24p9ZmW/SCN+EnnBRx8qIzqpA6PBH7lOUOI7wpPWNUaITfxI7LD6X/QFceSTZURBvidAETE0xxKebHcPa+qokerJfCdMSGNmqxEn4EcEMs7hqPi51HLGL9HBscYw8bQXdomM8M4QyUIEEm2hwRF+Hy7zXjYnNsv+pYzIZA4wWN7w+2zcI5sgEASCQBAIAkEgCASBILB2CESwWDuX54GDQBAIAkHgMCJQhHOn90FGXkxtgFd6cVZ4GjE4j6aYizw+w7FXPBM4kOtHvhU+TeASFxDiUtggYKW5gQFSVjSLFfrIb+Q2khbZLeoFMY7EFWUhjQ4i2OpygoXzkeNdC6ALQm8f1SiWgx4w+yIEjF9jlY/4h5+s5je2v7eMcCE6gIBEVJJGihAhCsDxGl8i3xHxrKOZCBdId8W5+ZR/CVT2d8RAi30iMdyTsNfzalx+4ev+rY/v6IwWVReFvokxr0bYD8Fmfo++RkdH7L/XXGycz3nHw6aPVxNE1A8MfrCMKOH5FdP2/PbD0PEwYN4PsNcIeaIkCBuiVkSEmQOwIVRIW+ee7kE4cjzsd17tmcf1swkCQSAIBIEgEASCQBAIAkFgHwJJCZUhEQSCQBAIAkFgxREYZLxVv4jBrFrf569ZRIVfmqhsQrNTIyGA/daRFosoFeeuA6kumqSeFRHb9RMQr53uyWer7ZG0xAmr0BG5SHBiBOLbuUhbx1iFb2W5/che57guMWSeUiiryr+2dwvcjFsEOBEBGd41KBDk0nWpsfCOMmmOpIpyLNHpJ8pEEGh8ZR6IvPBZ6iLX9vf/B4e/CE9IeiJV+5QQQnR6pIz/9UF/HNPF3M2nboQsfTRGEPkIe+cfLyHCvV5bW/uMN60XTPX48G7TP+OwUye5j33EB+NMH+Z1a/RLH9yHuY8+2OfZnE9YIPAYz4555zCRQISFfh8QLvQPVs7v4vHmxN+OPtknEsVYf6pMyi6RR/rknUIEeblEirUQQOtZ04JAEAgCQSAIBIEgEASCwNIQiGCxNGhz4SAQBIJAEAgCN4/ASOuD0EPyLVIZ3fxVj8YVBjb9ML0K/IoPJ5KijncMHOGJmBSpsjak+ky06PoFSFh/C8IAIY7kJVQsyNcy5Cuy129IWbghv6XQQdT67lxEceO/iADyPVFABzLP+KCLohuz/NI1RqQkIlYg3B0jVRGSvX0pSgaxjvC/v4y40SKUecBn0hiJyjAOCBYPlXXNEoQ8/xJCjAl+JW4QOXzXN/dw3Y2yZ8r0TwSOc/X3O8r0ybEEhP2EvmMIJLaeQd0Hx0hB5ruokbeUbZYRC4y9rqFCODNejUMYGJueS+onQofIFOPWGDYu9bvfAe7hOfXdMa5tPmju4V0rnRORQuotz+CZiT6OI650pNaiXksiKgZ62QSBIBAEgkAQCAJBIAgEgZtEIILFTQKY04NAEAgCQSAILBmBTo1yTUJ+yX1Y1ctfXql9PeT4ECcujIgMfwOdrM9rlbZoYLA9UkR1xAWhAjmMeGXIXaTtIqKnDBmM9EVoW4neK9C7ALTICgRur8TvVfKrOm5Wrl+vUtRaWqWOHOq6FPAW3aLIM1/xH+saFHz3U2XmCB+2qERwQOwTBogNfEvQQN7zo+MQ/XwsikMtDeLBRwdohA9EvigF5xFJjB+iB0L/R8oIDIQEwsn3lOmXY5xn+9i4FmHBfRxHICAKPD6O008CiPeea7uG33vsSc/kPNEm2sNlRBK1I5yr757FmOyaFB0JAS9CCmw8hzEt7RMhZLPs98Z9PZ/valK4t+Ph29FJl8XjVS9KPjDKJggEgSAQBIJAEAgCQSAIHAoEIlgcCjelk0EgCASBILCOCMwKbSPctKxanw2Em4iOQHoiL5GnyPu1SAs1n0Mj2qKFBWQx0hYpjLRGxCJmNSStvxet6kc4I8xbmHCeZovE7dXrGadzsA/+M5yNYbgTGtpPaoog/PkMmS89E0FBlIJ0XvxNeHJ+R21t1meiBUFEaqeub/K5+ixK4cfHOcYGEeJdZYQBhD9hg5hhXPidAGH8bJQh/4kBClv3+6s+LloXByduzJux5ZquQWQRPdKF3B2rb+8p88w+uzchgUDx/jKC2h+WeRbPa347zjU8O0Gli2qLPPEOcI7xrRYL0UI0xT+XeaZOb2Zsdzqqecqz2p0WBIJAEAgCQSAIBIEgEASCwEEjkKLbB41orhcEgkAQCAJB4AAQmKWCQrAhGNWu6JQlB3CH9b5E4YtQRWgiILcQ+OuKyIi26OLGXZcCYQwTBDdCl4ABMyRv1wywbQK3ozOM064bsq6Q3tbnrmgMPtK6DoQUTSIdRCWoC8Fn9iHipXsiSkiJhPi3T2QDAevby0RLOP6JMvUgjIXPjrEgQoMYYWwYJ2wZjajApHQiaoiQMN7eXGasqetBSDGG9Z3Y4jn1XRQKoUXqpz8uI5bYR6BwvOdUtJzQY1/X31AwfG3fCctwYq4ZBIJAEAgCQSAIBIEgEASuF4EIFteLVI4LAkEgCASBIHCLEBhihf9HI92QgFYvv7zOpPpBQz/SQiEukbuLXPQ3EbFx0N275dcbeLgvQppooSGFjUEYiapA4CLBpdpBFHdURdclQCYLV1mbuiC33FFfww2HgEFYQPh7n4hKQPYb93z6M2VSP/ErAYNfiRGiM4wF0TX2i9ToyAnHiGLga0S/FEwawt+YOYg2v5aICCKL96I6HOZuR2KIjCBESB3lmURJEDUcY7+xK1XUR8qMZc9EdPFeJYQQXC5GoDgIl+UaQSAIBIEgEASCQBAIAkHg5hFISqibxzBXCAJBIAgEgSBw0Ah0YWgko1XsVq1nte8BooxUHyQ98nKtim9fCcaBh58IEQSIrn3gO5La+OsxaGt/11VYCBYZowc4QA/wUoOIv1DChSgKZL8xL+oAob9R9k9lnygTQfFgmfRHnS7JlmChdV0TwgCxQpM6af7vCSLAQQkW82u5h3vps3sTTDbLjEXvSH3scarPRBkprp4sE4GhTwQ15zhXAfBFDZcUyx6ezCYIBIEgEASCQBAIAkEgCKwIAomwWBFHpBtBIAgEgSAQBCAwSwXVqVuQagj1CBYHPEQK645gkRPfam7RAQd8l6NxuZE2ChHMFinKyrogPLEiURWHyNUj6oIIIOJCrQoiBYJfrQifHyr77jJ1IswPJnKhi3s/UJ/Vp/irMpEPxA7nGROdWurj9fnHBiwErqstlJr/9id13PvKOpVT19YgOojk0K9PlnUhbMKESBC1L5j6Gp8a/fI8fzH65bOaHiIqthNNMbySTRAIAkEgCASBIBAEgkAQWEEE8q/yFXRKuhQEgkAQCALri8Aghq2AlnoHKWxVsXRF6wvKkp68sIYxclWz4nztIy2uBvUsTZlDFsLO2Lc4JeNzSYN0yZct4cKLxTwQnSAllOgJc8FWCiiFr6WDQvSrgyGtlBoRxAMFsB8pI14QN0QzOEY9id8u+0zZB8qkXHL+RpnIBudramR8U9lmGeHEtR8tU9D758rUzVBbQtQHEYJI8cGyx8qIJM53bcc4X/qnZ8ukiBJxYW7bSgnlXbqVaIoF7mlBIAgEgSAQBIJAEAgCQWClEQj7sdLuSeeCQBAIAkFgnRAYBDDyEHHn/9FWNZ/P6vXljILC24pvK8iRtVaHXwjWy8E6V11tBEq40EHvHHOCSUdHOLVPKiVplwgE95eJsjlbRiR4qkxUA2GD4OHd5R1GNCB0iHrw3fxyXZ+lpdLMPdcWYSECwj10hPBALPGdIEFwIEQ4/h1lxA/1K0T6fL6MAOK6+iwiYxGVNq67SF1WQsW4ZTZBIAgEgSAQBIJAEAgCQSAIrDoCqWGx6h5K/4JAEAgCQWAtEJitVkeed772rRDoS3U/whMZeqYM7ouogUQLLBXzXHx1EUD2I/qZOg/dCBTa02WEA78TB6RjMn+kUyNOEDiY64ho8Jti2c733f5OKeZ6IjnMQaKIiA2fu3aGItn2Ex8WtSbKRJu5j7RU3YcWJ7oAvOumBYEgEASCQBAIAkEgCASBIHCIEUiExSF2XroeBIJAEAgCRweBkQoKaY6YQwZqia5YsosLdwSrfPkd0bIbkWjJoOfyhw6BWQRG1yoxXy7XMJFqSXqpTrk0/3w9Dzuu34devu7sHv1vlv5t3o9EUFwPyDkmCASBIBAEgkAQCAJBIAgcEgQiWBwSR6WbQSAIBIEgcLQRKOK8U7BYKUy4SD2FW+DyUcdCvhjChRXf0tDsJMriFoCfWwSBIBAEgkAQCAJBIAgEgSAQBIJAENiHQId4B5ggEASCQBAIAkHgNiAgBVGZBQTSEskBz7LK/9b5Avb+HpITv9PZ3Lq7505BIAgEgSAQBIJAEAgCQSAIBIEgEASCwGUE/h+c8DHloh/riQAAAABJRU5ErkJggg==" }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOydZ5Qc1Zmwn0pdneN0T46a0YxyRAghRMZEG4NNcAIbbBZjL+B1WAcWe9cJr9PndcBejL3s2sbYGJtoY3IOQkgCoTzS5NTTOXdX1fejZxoJFEYgWRJTzzl15kzVrVu3urveuveNgizLdwqCcDomJiYme8EwjIcERVHixWLRfbgHY2JicuSiKEpSBITDPRATE5MjH/FwD8DExOTowBQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU8IUFiYmJlPCFBYmJiZTwhQWJiYmU0I+3AM4mhElCZfHT1UohNVqBUMnlYgxMjRILpc/3MMzMTmomMLiAKlvm8UpZ53HkmXL8XqcJKLjjI2OkMvlEQQRl9dPbX0Dol7khSce5M7f3sbYeOxwD9vE5O2jKEoCMMxt31vL7KXGTb/8o/H9m28xzjz7bMPv8+yzvdXhMc648HLjf+5+2FhxzILDPn5zM7e3symKkjCFxRS20y+5xvjl7X80ZnW2HfC5nppW47Z7/m54bMphv49DvwlG+6x5hkWWjoCxmNvB3BRFSZgKzv0we8W5vP+sY/j0ZZewcXP3AZ8fH97BC+v7mDOr+RCM7sji9A98mhtu+iGfvPpjh3soJocAU2exHz5y9af5/lc+RCZfest9DHRvYmw8fhBHdfixuYO865yzEYXXC9q97+NX8Phf7uDMc99P73jxTedsXvssG17b/I8cpslBxBQW+6ExaGNzz9jb6uOuX37nII3myEHXSiRiUSZlhcXbiJLspbu7G11+F/FY5E3n5POmhehoxhQW+yGWhfoqF/3h5OEeyhFFPh3lkQfurvzfuvg0Nq718Njjz3LpRafz8P137+Nsk6MRU2exH371s59y4w9upq666nAP5YjGW1VNbGyUmpZWhnbuONzDMTkESJIkfVHXdfVwD+RIZXD7qwxEilx/wzdZtmwJNqsVXStSLJUoFYsYh3uARwit848lKOeR/G1kBl/llde27rVt08z52MQiqUz2HzhCk7eDJEkFQVGURLFYdB3uwRzpCKJEW9d8lh63ks7ZcwhV12C32ygW8uSyGRKxCKNDg/T3bGfD2tVs27IN3ZiaKFEUC8ViYb/XlwQoadpbGTyyJFIqvXUlLQgoikSxuOc+VlzwceZ7M/gXv5s/fvtqtvS/WWcBoLpC3Pz7e+l94U/c+NVvv43xvBlZsVDaz+do8tZQFCVp+lm8zc2iWg2312fUNbUaC5Ydb5x38eXGjT/4pXHzbb816oK+cjtBNBatONlYdNwpxrd/fIvROaOxcv6CE8837n76FePYhTMNwGjuWmxcdtU1hstmqbQRZatx40//YPz05z8xBDBEWTXOvfRK44Tjl+82lqZZS42v//hXxqWXXLjLftH47Hd/bdz2u98YAhiIsnHGhZcZp5928m7nzli40jhuWdl5bPbSFYZD3dUvRDCu/uqPjd/ddZehyoKBIBonnXepcc45Z1baLD7jQ8bnPvcF45bf3V6+zsQWap5l3PjDW4yPf+IKQwSjedHJxt1Pvmz87YX1xvf/+3+N5XtwWGvsmG9c9sl/MS686CLDtss4nL4a46rPf9347s9vMy5473m7ndM85zjjD4+tNd5z9kkGYAQbO4zLrr7WCAV2d55T7W7jnIs/alxxzbVGe1vTYf/9HC2b6WdxECjkcyRiUQZ7d7Duhae55/e/5mvXX8Fv7nqMK//pCgDed/UNvPfcUzjroo+z5rknufraawEQFAfX/su13PHb/2Pm7DmEWubx79/+Jr7G2Zx71qmVa6x892UU+15ArmnDIgp89As3Mbs5yBWfuxFVmmgk2fjyN2/ijp99h5M/+GmCTgsAC055H1WlHpL2ahxSeSwrFrZxybU34FYmzZ4S//TZG0iMl60+H/zkv1LltVeu37HsXXQGivRnZTx2lbM+fD1nrlrEe676IiGnAsDoUB9nXHoFT913B0blTJHPfeMHPPTbn9K+8gLaG6voefkxvvWf/8Wz9/2O/739Xt797nN3+zyPO+dD3PgfNzK8czNqVSvHLJkPgGz38p+/uI2edY/xna99BdkdZPLWESSu+dcb+ONtv6Bz7nwc/nq+9aOforqr+dAHLq707fDV8L1f3UGt18L27l7OueD9b/l7n46YwuIQ0btjBy63B9kR5NxTFvH1G/6NzVs347GqeBtbEIDjz/4gI+sfIZaGbDrJ9V/9Jj/5t39m3YaNyMqEGkmQuOCiS7n3zjuRiznalp7BwiYL3/vOd8npQuULnLn0ZJzZPjbtHMUmlEjnNUDgI5+4iv+79RZUXSPQsYwzV3Twza9+jWROQ5qQFXVdx9DiSbNh+yAg4HY5SGcylXt534eu5M//92tUBJx1Xbz/3OP59698ifFUFnnCdppO5XBZSvzpj69bQYJtC+nylXju5U14nVbiyTRgcNLpZ/LwX+8DQSAcDlfah9oW8eUvfoovXvVh/nb/vSTDAzz97EsAvOfy69n06O389W8PITtDZMZ6mFyQ1XQsp5YRtvfFyKbifPwL/8HdN/8HTzzzPLLldXXcVV/+Li/+5Wfc8vOf0z84yiP33QWAI9DM1779zYP0zb9zMYXFAeCvCk2pnaw6+OjVV/H3++7F6vSQi4cpaAb3/M//o33lu6mrbeFfb/oJH7noFL7/3e/jDYVoX3wmpd5neWH9FrwuD+ls2VR7zBkXk+t9ko0DcYwSXHX99fzk2/+BJqhYpSJFDUTFxtXX/QuOQCPf/umt/P7HXydT1Fhw8oXofc/x6pYhZEHkqi/8Gzd/6wYKuoDTCpmigSAqfPLzNzDaV/ZOVd3VzGitQ1HKM4aW+atoccV56sVXUVULl137JW77/tfI5Et47QqpggaIXHX9dfQPJ5k7q638IQgSV3/+K6juAF/70a08fedPGYllaZm/ikZbjKdfWI8/UE0sMlJuLqtc/9Vv0f/qasbiGVR3HZ/6zKeRRAGbt5bLrriMdatfAODEcy5k5QknTFxH5qrPXM8tP/khnlAIb9182r057n3wid0+x7aFJ3H+eSfz1MOPAnDuB69i9sRYP3Ltl9nw7KNv78cxDTD9LKaMwJVf+j4tAZEnHvob69espr+vj1QyiW4YqDYH1XVNLD5uFWe/5708ducvePCx50FUyNrqOetdp7Kxe4hMOsmvf3Qba9a+ytbNm9A0nWBVkNNOWchHz1oJwNDQAGctXcFoMcCVV36Az11xMaqjgZa5S3jqjz9j044hQCJVsrN0+bGccsmneO3vvySy7CISG+7lgb8/ydzlp/OZa6/k8x97P4Lqp769k+hDt7P61e0AjMdKrFi5gnnv+gjp7udoPHYVC5ccwzkf+Wf6undw6eUf5fEXt3H1ddfz7esvpyQ6qWlqw4j8nSeeW1ce50iS4084gYZj3401vJZ//uT3uOk7PyT/jRs55qwPI4++xN3jrQRL3fzu93+hfcEKvvjVG/jWdR9GN2D7pnVc9JmP8vz6Ps7/6HWMbXicxpUnM2/BIs6/8nNY0TEM+Kcv38TA5vWsOPUs8t6ZnHH8PGSbk8VLlrD8vMvJb3+Cx59bxyXLLuKU897DZz9wBroBI8MDdJ13AUtXDXPNZ/6F559+gRWnnk5Lzs15Z5/CTx+/lfYlp7G0zcpVX/374fphHTWY1pADJNTQyvITTmHOgoXU1dfjcDoRgWwmxehgH+tXP8ujf7uPSOx1Jy5XoI5LP/YJqjwOHr//Dzz9zAu79bnirIupsab50133AiDKNj7y6c/hUzV+898/ZnQ8jmz1cM1nP8fvb/5PhsNl1/GOhSt5/8Xv4+Un7uOvD/wdqyfIJz//b8yZ1cnwzk3c/L2v0zswCqLKp750I/f+6gfsHCjrJRq7FvPBj3yEzasf5S93/YXOpSfz3gvezZrH7uWRJ17kQ1dfR8AhccevfkZP/zAICh//7Fd44k+3sHl7HwDVrbO5/MqP0/Pqc/zh9t+jGTBj3nIuvPgiBja/xO9/81sE1cWVn/kyS5csJDK4k1/+v2+xaevOyr2fcO6lrFq5jJceu4+//fUhFq46h3POPp0XHr6HD376y/zi57/m0nOWcN11X+TSq64j5JL4v1/8F866WVx0ycVsmhi/bsDsY09n2Zxa/ufW28p6E0Hiwo/9MzMa/Nxx608Jp+Gjn7wWLTVCwdlE8rUnOPOj1/HNT13M1p7hQ/abeSdgWkPM7QjeJOO3j79m/O7+h42Qz3nQ+7/kX24y7n1yrXHJBWcdAfd65G+mNcTkiMXi8OF2qfzgS59iNJo66P37AwHWP/4nfv+nBw563+9UTGFhcgQicO03/gt7coCX1m086L13LT+bS993Hs88/HeMg977OxdTWJgcccw54T3Ui8P0JzSE/Tc/IETFzvVf+Cz33XMPomj+/A8E89MyOcIQ+djVV/Oz732n/NY/yNJixTkfYMezf6Z7IIwgHGxR9M7GFBYmRxSN81aixjezuWcMYcJ0evAQueDii/n9//4vkiiivZU4m2mMKSxMjihOOvPdPHLvXSCqCOQOqrDwNs7BXRxg51AUp91GOpfZ/0kmFUxhYXJEsXDJQla/8CKKJ0gpNop+EPuevXgZG1Y/jQH4AzVEwqZvxYFgCguTIwgRv0NiNJqmub2Lvu6958R4K9Q0NtPf3Q0ItDYH6OkfP6j9v9MxhYXJEYRBoSTgsFk558KLeeqRBw9q7/lMBqfbTeuikykNbSCWfTv5PaYhpgenuR1J22kXf9L4zf1PGP/2tRsMSTi4fXuq24yb//Cgcesf/mJ0tNQd9ns9mjZFURJmbIiJicl+URQlaS5DTExMpoQpLExMTKaEKSxMTEymhCksTExMpoQpLExMTKaEKSxMTEymhCksTExMpoRoGMa0ERiiKNLU2o4oSftvPIGsKDS1zjiEozowbHbH4R7CW8IMBz+6MQxDFHVdn/qTc5RjUVW8fj/zFy+b8jkdXXOIjocJBKdWBuBQ0zKj45D2ryoQcEN9UKEhKFLjB48DpLf5SjEObqy5yT8YXdelaVUKwGq1MzTQR219Y2VfVaia8Ngoe4uFLhTKtTPHx0bf9vU9Pj/x6J5rgL4d3F4fiXhsr/ewP0QB3HZw2MBmVVHsIWRLeQZTyKXxCjp6MU0iESeRNsjkD+boTY4WJEEQvmIYxrQQGjPnzKO1fSY927fh9niZMXMWCAIOp4vOOfPp6JqNqloZD5cFg6JYCI8O0zVnAalUkmNXnkgsMs6chUtwe714vH5mzV9IJDzGsuNPRNd12jtnoWs6VpuNQDBEVaiGzjnzyGazHLvyJCLjYeYtPgZFUWhp78QwDOYuWspQfy8nnHomiViMto5OGltmkM2kWXLcCfT37gDDQJIkvL4ATreb2voGHE4XTS0z6Jo7n+j4GLnsgednsKtQVyXh8bpRHUEszlpEyQaIKIqKbLEhKXZkixuH04PdkkeRCuTyoJuThWmDIAilaaOvAMhlszzywD14/QHmLVlGNBJGUSzMnDWXfC7H0EA/Bq8/ATNnzwWgpJVomdHB8OAAzW3t5LIZ7A4XXXPnk0mlmD1/EfFohIamFrKZDNV19bjcXto6OmloaUXXdWw2O+tWP0/XnPnEImHaO2ezfs0LBKtrKeRzzF24FI/Ph2Kx0NDUglYq0dDcSi6bwdDLWR0CwWpi0QhdcxeQzWSw2uzIikzfju1Ex8N7vOd94bZDTUDC6m5AstZhsfmRZQuGYaDrOoZhoGkagiAgiCJFXcLiasLt8VMbAGVavGJMJpk2wsLhdOHx+WhqbSefz5GMRcllsxQnlhk2ux2LqtK3c0f5BEHA7fESqAqhKAqyrOD2eFGtNgb6ekglE8RjUXRdp1gsMjw4gNVmp1gokMtmaWxpo793J6VikWwmjdPtQpJlUqkEYyMjDA30oWsaVaFqqmvqaZvZSSaVQrVa2bppA6VSEZvdQaAqWFEOVlXXUCzkiYTHkCSJQFUISZKpa2w+4OSzbjtUByzI9jokxYnB60rIyb5yuRzJZBJN0xBFEYvFgiBIKPYabM4AdQFQpo3Gy0QQRTGr67r1cA/kUCNJEo0tbQz291HI53C63GQzaSRJRjcm8jEZUCoVK+coigWPz0d4dASrzUapVELXtMqDZUwsDSRRwsCgVCwiiCKGbiDLMgi8vs8wUGQFURIpFYvohoFWKrHkuJVkMxm2b3qNYrGIIApopRKyrDBr3gIkWWbti88BIMsyisWCLCvkczlOO/d8nn7kQQqFPNnM1JcgVgWa6pxgqUJW7FgsFjRNQ5Ik8vk8giCgqirFYrEys1DVcoFhwzAqWy7ZRyYZZSAM5orknY0oirlpIyyORNq75mCz2dny2ivk87ndjjU0teDxBxgZ7Cc8OvKmcxcsPZZSsciGdWsO+LpNIQmHr4lcAdxud2UmYRgGhUIBWZaRJIlSqVQ5JggCgiCg6zq5XA6bzYaua2SjWxmL5ogd/DpAJkcQoijmps0y5EhkoHcnyUTsTYICYGR4kEI+v0dBAdDfs2Ovx/aFyw4OlxtRtuHxeND117NcapqGoigYhkE+n6dUKlVMnvl8Hl3XEUURm80GgChKCIofv+vtm1ZNjnym5Vfs8nj3edzpcr9pn2Kx4N7PeQdKNpNm5/Y955ksFgps3fjqbvtq6hpobGkDyqbckaGBPZ7rCwT3ek2vQwDZg6JYKJVKJJOvF3CW5bLGUhAERFGszCYEQUBRFICK8lPX9fJ+mxcEBZdt6vdtcnQyLYVFW0fnXo9JskywuvZN+1vbO8nlsodyWPulKlRDapeHe280tbbtcb/LBk6HFUm2A+UH3+l07uYwVSwWEUURSZKQZZlSqVTRZ0wuSUqlUuV8SZKRrFX43ebs4p3OtPt6JUnepzdhVaiaSHgMYDehIcsyhQnlX80uTl2TWG12XG7Pfq8/a97CitUhEAxhdzjxeH1TGrsoikTHxwjV1O2zXalYVtK+0cXapoJssSKIUsUs+sbPYlKxOXm9siXodRvppLJTkiQEQUDTNHRBxWGTEd/g0S0IApIkoSgKiqIgHYCbvcmRx7RyyqpvamHpcSvp29lNTW098xcvw+5wYrGoJBNxAFpndNLf0w1AbUMjoZo6nC43oZpamtvay/00NjPQ1wOA2+Nl+aqTERAo5PMsWLocu9NJdW09/qoQ42NlvUJbRxftXbNJp5L4/FW0d85G1zUamlsxDIOaugZqGxqZvWARhlF2M5dkmUQsCoKA0+Umk0kTCIbonDOfWCTC8lUno+s6cxcdgyAIdM6dD4bBvEVLGR8dZulxJ+DxeEnEo2iaVp5ZON0YoqNiyVEUpfLQG4aBIAgVxebkUmRyP5T1GpOm1Ml9xUIBVcoxHi+i6aAoCna7Hbfbjc/no6qqikAggNPprJiaTffvo4tp55RVFaohEh6jkM/h9npxebwk4jEy6XSljTah1LNYVLSShsWi0tO9FbfHRywyjkVVWf3cU5X2HbPmMtTfhyRLBELVRCNhrFYb9Y3NDPX3Vtr5AlXUNTRhtdmpa2xmeKAfWVFIJ5P0dG+jvXM2Q/29SJJMJp3EZrczMjQIvL5sioRH8QWqGOrvJZmMI4rlpUGhkMPr87HmuaeormtgeKCPUE0N/kCAVDyK1WrFYrGAAAZa5YGfnDHsKgAm9RGT5lF4fYYyqa+YxDAMRFFEVmQmjaeCIOB0OvH7/Xi9XtxuNzabDYfDgcvlwuFwmDOMo5RpMaOYxGazUdfYTKGQxzBgqL8Hrz+AYRhEI2EEQaSlvYNCIY/L7aGvZwdtHZ34q4Js37IRRVGwqFaC1TWMDJaVi9lMmkwmTaimFk3T6NvZjdcfwJF07WblcLpcbN+yccLz0kY2myFYXQMC+PwBEvEokizz2vo1iKJEPBqlVCw7jKWTSVonBMbwYD9dcxaQTMZZ99Lz2B1OErEYdoeD5rYOSsUCFouCLxAkEY+RSiUpFAoTlg0wtAKSIlX0DgC6rpeFCWV9hNVqrZhJJ5Wdu/pXTC5BMpkMdrsdURAx9GK5/wlLis1mwzAMSqVSpX0+nyeZTO52bZOjh+nlZyEI+w+2EgREQUDXyyUTJqfhB36pvZ+3p2Nv3Len/2HP0Zu7LhUmj08uEyZnCQBVbgj6FQR7O6JYXoJomkYymcTtdlf0GJMKzmKxWLGETPpfTFpHoCxYZFkmkxpHKvSypR9KE7WGd509TF5/19mKydGFKIq5aTWzmFJUpmGg79Lurf6493Xeno69cd/+/t/TsV3b7LpcmCSeBo+ziCDEcbjL5lVRFLHb7RU9xeQMA96sIN1VUAAVa0kuNUoh/7qgAMwK5e9AppXOYrpT1CCZAS0/jq7rFaXm5EMvSVLl7T85a5jUa1gsZb+MfP71+PRSqUQqGUMmRzy9t6uavFMwhcU+mKpJcxJfoGqP+/dnUvX6Awd0HSgHximKgttzYGOMpkA08pQKqYqwKCt0LQiCULFUTAoQeH35IIoisixX3MLT6TRGYZxcATPHxTTAFBZ7QZKk3ZLkTIW9pd9rbtt3dqu3kravvqkFXdf36oC1N4oliKWBUhxjQp8xGTAG5fve1Yy66wxkV12GrusYpRSikWE8ccDDNzkKMYXFBI0tbdQ2NCFNJA9rbGljcKDvAHoQKuHuezi0V7w+P+HR4f32LooiXXMXVP6XJAmvP0A0Mr5fJ603Ek1COp1CEl9fhkx6Z05aPgRB2E2hOakwnRQcpUIasRQmmoJccT8XNHlHMK2csqpCNRyzYhWGUXYMamnvYO7CpahWG/lcDq/Pj8Wi0jazC6fLQyAYYnAXXwmAzjnzmT1vIbqu43C6UK1WFixZhqaVJs5zMzrhH1FT18CS5StJJxM4XW4WHXMcqtWK2+MhFhkHoLG1jYGeHtpmdrFw6XIEUaRzznxy2SxtHV20ts/EMHRaO7rQikX8wRC1DU0Yuo6qWhno3UldYzO+QID2ztk43R4amlr2GjcCZY+IdEbDrmooFgsGYkUhOumMNRmaPhlMNmnd0DSNfDaGnhsintKJ7N/73OQdwLRzyioU8gz09WC12uiYyI6lqiojg/3YbHZq6hoIhEKsffE5QrV19E14ck5SFarB5XLj8nhwuT0sXXECoZo6Xnr+adxeHz3bt+5mBaipbyAeizI6PIS/KoTb4yUejeyWe0KSZBzOssu3y+OlvrGF6HgYf1WQdCpBMpmga+5CnC43ikWltX0mo8OD5XgNWcZqs5PP5ZAlGQSBjq459O7Ytsf731VhWdKhZyBGIjoMWhr04m75KyYFhSzLlXwXuWyaVLQHLTNALKnttvyQZRmHw4HH48Hj8eD1evF4PNhstsoMxeToZtrMLARBYOUpZyBOxCt4vF5GhgYJj42W39ztnQwP9FEVqiabyeDx+pBkGa/fX0nWO3PWXEqlEol4jJr6BsKjIwiCiN3hQJZlBnp3Issy8VgUgIbmVjrnzCOViGOz2RkfGy3HW1gsRMbL8SeNLTMIVtei6zqR8BgCkM/lKBULNM/oIDI2hs8fQNd1tm58FbfXRyqRwOPxYVEtOJwucvkcdQ3NyJJMLpehf+eOSnzHJLIsV5ytJgWaYUAiXaCUT6JKWQQji65r6EhIklxZkmilAsV8HC07QCGXJRyHxBty7UiShNPpxOVy4fV6CQaD+Hw+gsEggUAAi8WCruuVBMgmRxeCIJSmlVNWeYotoWmligPTri7NwuS6vFSaWKdLdM6ex2uvvFxp83qchIAgChi6PpEdS3+TL4QoSsCki7SAIFBRGu7axjD03ZyqBEHA56/iuBNP4f677tjtmCTJaNqkmRPAQLXaOP7k03j+qcfJpFNob/CQlGUZVVUr7tr5fH4PYwWbZTLLt4SkWBBFC4IoUSgUiSfSJNI6heKes2IJgoDVasXlcmGz2bBardhstkpoO0A0GmXnzp2mB+dRiJkp6wjmmBWryOfzrH/p+f22nb9kGQIC69e88CYhYLFYsNlsiKJIqVQinU7v0WFrEkEQkCUQBQNRBE2HUmnqmbwnlaGKoqCqakV4KIpCPB5nbGzMnF0chZjC4gjG6w+Qz2bJTiG9v83uwKKqb6pJIggCLper4pWZSqXI5d6clWu3viYESyaTOWiu2ZIkVRSkZsTp0YmZVm8f+PeQbcrucOL1HbgDlSiK+Kv2nr1qV6w2O06Xm1hkHJd3apm5spk08WjkTSbUyfBzQRDIZrP7FRST57xx+QC7Z886UDRNo1AoUCgUTEFxFGMKiz0gyzIe35s9IxubW0kl4wfcX21DY8V/Y3/4Jrw5RVHEc4DemaGa3TN8lUolstks8XiczBSyf08Gje1JIAiCgM1mw+fz4XA4TOvGNGTaCYvJH7kgCKhWK6Haut32A9Q1NDM6PARQeVsLgoAoSZQ0DVGSKolwdsUXqKKxpa2SYWuyz2B1XSUJzm597uFN7fb68AWqWLRsBU1t7cxdtLTS165tBUHc7V4E4c1f5aT14UDe6JOzhzfOLCb1HKqq4na78Xq9psCYZrzjTaa7Mmv+ItxuD+PhUapr60nEypm1q4I12B0OVj/7JABur5fendsB8FcFqW1oJDI2RnVtPdV19ezYugWvz08PZX+GrrkLEEWRSHgMj8+PoqRYdMxytm7agC9QRW1DE2tffBYo1yLx+gPMXbS0ksLvyYf+SqGQp3POfJrb2nnmsYfI53J0b91MqKaWxceuwOevQrFY2Ll9Kz5/gKbWGYTHRnht/cvMmruQ0ZEhhgf63/ZnZBgGqqqSzb4532g6nUaWZbxeLw6HA1EUGR8ff9vXNDk6mFYzC6/Xx4vPPonN7iAWiVAsFti6aQO1DY1s2SWT9vF+xNwAAB5USURBVKRpz2qzUyjkKRYK9PV0IysK4ZFhFIuFV15+sdLeMHS8/gCtHZ2UikVi0QjpdIpUMsHo0OBuKfvrGpvo6d6G1+dnx7bNjI0Mkc/nkBUL3Vs20dO9jWQiTiAYqpQJaGhuI5VM0L11M6PDgwRratm+ZSMjgwO43F7CoyMUcjli0bf34O5aG2RvM5FEIkEsFkMQBGpra3E6nW/rmiZHD9PGKQvKyrvoeJiGphZy2SySJKFrOnaHg/DIcCUh76JlxyGJ5UCy8bERWts7iUUjpJIJEMo5dBTFUv6f8pKgWCzg8weIhMPkshni0SjFQpHZCxYRGx9nbGRyWVOLIAiMDA0giiLFYpHw6Ai6pmF3ONFKJdKpJG6Pt+xharWSSafKqf8Mg9GRoYqvRLFYIJVIoChK5QHPZt56rLgkSTgc5erp5f73HPRRKpWoqqqqBJ2lUmaFoXc6084py2TfTCbCURSFVCq1V2EBYLfb8Xg8pFKp3WqPmLwzMf0sTCooFgtVwWqcbjc2m510OgUGKKpKIZcjk04xPjZKsfi6Q9WuuTkPFS0zZrJz+5Y37bfZHVhtNmx2O4N9rwf7NTS3MtjX8ybHM4tFZfHy40nG4yQTMXp3bD9kY34nMv3S6pnshtVqo7F1BstWrGLJ8pWoNhs+r5dQTS1+r4dSsUAmnWLT1u3ouk42neLFZ59i9TNP0NfTTX4KfhtvB1lRsNnLBZEUxbKboGpoLgfcSZKMrCiVWiker4/+nh1v6qtQyJOIRXlt/cssWHosA7096Pqb66aY7B1TWLxF5ixYTLFYJJNO7fHHuS8amlsP+JyDhSiKtM3sYtWpZ3H8yaehyBLb17/II3/6Nc+v24DDH6KltZWL3nMeL6xZy+rVL9K9YweKJDFn7jxWnHASZ7/3/RTyeZ54+G889fDf2LFtC4axdxfyyaxb5bIBCoIgMnfhEja+shZZlslm0qjWcjZwp8vNyNAAgWAIp8szEawnUFPXwNjoMGVrrUB1bT0g0NO9leqaOqKRcaA8y7E7nGQz6XK+j/EwAKpqrVSUy+dyBIIhMpkUimJhxsxZbFi3hlw2g93hpJDPIyvlolL+qhD5XJZ8PoeiWMjncigWC5n09NPTmMLirSIIbHntlbd0qsfn301Y7PpmPJSEauq45KNXsfLk0xnavIaX/nwLvRtXYzHyeC0iMwMyL0fj9K7dwLJlx/I/f76vHMQmqmQMgWdeXs+zL76I125j+fIVnHDKGZx34aU8+uC9/P7Xv6hE576RjllzUa1WxoaHmDVvIePhcjtRFJm7aCnh0RG65s7nlZdXl53RfD4y6TTB6hpU1Trh1eqirqmZdCqJLMvYHS5sdnvZ1Gu1MXPWXHp2bKO9aw6+QBXh0RHcHi8vPvMEUE4XMNRfTmakWm0EgiGCYi2DE8WiNE1j0bIV1NY3MtC7E4uqEh4boVgo4K8K4nS5KeTzNLe1Exkf45nHHjrk39eRxrSyhkC5ZGAum8VfVYUgiNgcDuYvXkZ4dATVqmJRrThdbjSthK5pKIqFhccsL1ss9HJot0VVae+cRS6XJZ1KYnc6sahqJVOW1WbDolqRZRmb3Y4/ECQ3USfEMAz8gSqi42EsqhWLqhIIVpPLZrHZ7VitNmbOnsfocDmBzq4ZrGRFwWq1IUoibo+X3BTiRqBsEj35XefwpW/+gOG+Hbxw18/RNzxAU6mXjoBMjdeOy65iUVUSmkwGK8cuXsjTL61FECWQLQiSjKCoIKsYkkwqHiE8NEAmk2bp8pVccOnlOJwudF3HZrcjTzh1FYtF6ptaaG6bQSadYmxkGF3XyOfzqFYbUC4/sH3zRvp7dlDb0ISqWtm68VXaOroYHuynUMiDAf6qKuLRCCNDg1hUlXw2gyQr2OwORocHKBaKiJJIJp2muraeV15eTWGidktdQxNDA/00t7UTj0VRVSs93dsIBINoWglZknF7fYCBw+liPDxKeHSYmvoGBvt7ae+azcb1L+P1B0jG4/tMLvRORBCE0rQSFi0zOmhobsNmd9Dc1o7H5yMaHiNYXcPo8BBnvuf9jI4MMW/hUrx+P7lMhvauOUiSyPBgf0VpVtvQRF/PDtLJBAICZ51/Eds3b6ysqRcsXY7d4WD5qlPK1ca6ZiOKEg6ni2B1DVabjdr6Jqpr63C6XFitNuYuWkpDcyupZIJcNksiHgPKb2XD0Gnr6GL+4mVU19Zhd7iIRSPkp1CoWRRFPvTxa7j66ku4/9c3sPOJP7LAkWVOQEIUQEfEEEQkQ8MqaCQzOWJFmZbGRl566SWsFgsBn5fOmZ2ccfoZHLvsWOYvXIxqdzIyMsJLTz3KX26/jR3bNnPFpz5LeHSYZx9/mGwmU8my1dLWTm/3dtLpJKPDQ5RKpfKyYmQQt8dHIh5lqL+X5rZ2SsUCqrUsaBOxGCWt3Ec6mcDl8RIeHaZzzjx6d3bjdLuRJYlYNEJbRxe5XJad27agWCwUi0VKxQLpVBKLqjJn/mJsdns5GdHQAFXBUNkpbnyM+qaWCZN1ilgkQnhsBE3TcE8kWpblcp3WbDbLjon+o5HwIfqVHplMO9Np19wFuL0+ZFlm84b1iGK5UpbX5ycyPobb48Pr9xMeHcHhdNEyo4MnH/4b9U3NbN7w+pKjraOL7q2bgHLxZKfLxY5tZY293eFk6YoTePn5Z2hpn8kra15kzoLFyLLCupee57hVp7Bl4wbqGpsIVtfyyssvopVKHHfiqfTt7CaXze62vJm7aCnVtfVsWPsSnXPmEx4dZuf2rVTX1dO9ZdM+71cQBN576WV85MPv5pW7r0PK9eIuglXz49YsZPNFYlmd8ZxBUNWYUV/NDksLT4zbqZsxm2eef4FMQUOULSgWhS1btpDMFzAEEYoFKBUgkyj/BWbMnMWN3/0Jt//q59x/1x3sOfOFydGIKIq5aTWzaGhuo66hiYG+Hgxdp76hibHRYRqaWkjEYwwP9CGIIjZ7OVCqWCgw2LeTlvbOcgasiRDwxtY2gtU1BKvr0HWN/t6dGBVTnUFVsJpMOs3wYD8erw+n24OmlXC43ETHw4iiyNBAH/6qIMV8gXwuW15PGwa6pmNRVdKpsu9CIBiiUCgwNjrMyOAAuq4Tqq0nNj6+XyXbiaefzYWXfpD7//sqqm2DuOwgqyDrOaLpLIMjWXLpLNlMDhcFQl4XFqePLTv6GU2M47drvLJ+M7XV1VSHQvRsfIVcfBzyWSjmoZCrCAqA6HiYZx9/mE9+7iuMj43Qt7N7H6MzOZqYVjMLi0VlzsLF5LJZNr6y9nAP55Dj8fn5+e/u5n+//ykWBtcypxkUGdI5yBcgmQJHCga3g6RDwApzjllJ1WlX8vXPXUNKcaEqIn9ZM4hu7Lt84htZsnwln7nhG3zikvNIJ806Ae8EplU+C68/gNcXYOf2rQelv13L/B1MrNaDI7c/eMUn2b75VeqU9bTXgUUp1wxRFXDZIeCDhANq68FjBasEw7oTb+s83vWhTzK/IYRLteNQy4rKA3G+evnFZ+ndsZ1LLvvEQbkXkyODaTOzgH0XKz5QRFHcZ3q6t8rBGKPT7eF/7vo7P7zhCt7V+Qp+N4xGwa6W41pkqZwuz2mD1zZCp+Jm0Xuuo6/k5KGHHmFb7yDWXIRNQ2Ul60giS6ZwYLVL5y1ayldu+hGXn3/abtnMTY5OptXMAvY+hRYliZo3VB9rbuvYZ74GXdepb2rB7fHidLkP+RgPhJNOP5vI+CiJkQ1YFMCAXAHS+XIuzXgaWmqgusrNinM+zDFX/4j1D/+J3930eX5z998JD/czp87HkpYqCiWdQunAheJr69eSzaRZcdJpb/t+TI4MpoVic3/4A1WUisVKlm4Ap9u93wfXHwhitzvo6d5znY7DgSCKnH7u+dx75++o8RvYVfC5IJ4BpxXa6yGWsTLz2MsJNCzjrw/cz/svvxJLvsRoDjJFDV3T2R5Os64vxmjGoDTVbL27oGkl7rvzdk4753weeeAe0636HcC0EhayomCxqJSKRVo7ZiLLSiXT9M7tW6itbyQWGUfTShi6XrbX75KJ2ulyUyiU/QDyuSzFCZ8AcSIZ7T8ap9NZLv6Ty1UeRo/XR9vMWXz1O9/BFlzJsfmXcRRSZHJgVSDUcjyLFl7Dq8/dwX1/+gR3PlGip1zCBLvTz4zmZlqbGugzqljWplKbkomO9hIL9xIe2UYhN3U358cevI8Pf+LTOJyuSji/ydHLtDKdzlt8DMHqWlxuTzl7di5HKpnA7fWSiEVxulw0tpQ9DRcfezxer5+R4QEUiwXVaqO9aw41dfW0zOjA6XIz2N/L7AWLCQRDUzIT+l2wsB1WzIbj50IqV14SvIUXN4sXL+b666+npqaGnTt3VjJbnXLmefgaZ3DvlkEKNbPIpArkh/poqPVx8nu/hM3TyhN/+ld+decr/Plpne5hsNoDdCxYzruumkftzEZSxgLsnhBFaxCbO4DV6cWq2nG5a8ll4hTyUxMY+VyOk844h1hknB3bNh/4TZocMQiCUJoWQmISi0Vl9bNPMm/RMWRSKXRdZ6C3B4/XRyBYjcPpZNumDdjsdja+shZFseDzV5XdsG12DENH0wyG+npBEIhHI4wODexzim2R4Z/fC+87UaatbQaSWkVBkxkbHeDCVduJpwxWb4ZH18GarWXF4/6YP38+N910E3PnzsVisfDHP/4RmKi6duqZ/P3Fl6FjKSVfNWv6VDqrZ1J92mnc9+oDqDv+xKPPZXn4ZcgXBQLVM+hcfBb+hmrcNWsoFrtJRLwUM/UUi3lkRcfi6qdlRpTEoAOLeiKvrbmffG7/OSw0rcRjf7uXE08/m4cfuAfTSevoZlrNLAQgEY9RFaommYhPJL0Fn78KXdNIJRM0trRRLBYqbsND/b3EohHsDiedcxYw1N+LKEnkc1lEUSQQrCYSDlMqFssxDLswvxW+8mE4ZdUSaLyOHv3dxGznIdRegtr0IeLKSSQKfoIejVPnRljWpdE3BmP7SCAeCAT4+Mc/jtvtJhwOc/PNN7N5c/mt7XS5ufpfv8Z/r95Grnk+XTNaufLEhWwdSfPDe59nICMwnLLx7ON9ZPJQVdvJ3OMuwOr2UCxA/2tWxnbUoshN6Fo5taAjMIq7SqRUzDPzhFFiIzlkvYVouGefkaaT5HI5Lr/6Wv58+23/kGA5k0PDtJtZDExEGG5Yt2a3/btGS05GIQK7RYZabXaG+nvYumnDbudGwmNvuo4gwPnHw+XvEik4T0Ge9VU0Q6be6aSxsZH8RPq+lSedTWrpKtatW8fY4CaaPHfxjdrHuO1BjXuehdIbrJWiKLJq1Sqqq6tZv349t956K319fZXjS445llS+gG518k8L68hJVr73yIvkS0GMqma2lAw29yTRchKKxcKsZasIdWjUdq0l3CcQ2bmQUkGkWMiBYSAIItHhDJnUMIGmMfJZhdmnQqmgUSisoHvjE+xvttDTvZVcNsuMmV28uvalfbY1ObKZVsLi7RAIhhibKA+wPy49GT5yTjVVi/6DtoXvQ1XVSjJcwzCIx+MkEglsNhtOp5NZs2YRCASAFQxseoBL9W8R8qb45QO7CwyHw0FLSwt9fX3cd9999Pb27nZdb7CG9oYQFxy/iLv7MgxGhjEsDigmECxWjGQEPTYGhoavqon248bwNmynVFDwVbdgd0YY2NBYFhSiiOqMEAmvxsBOOipSzFQTHy1h8+/E7W/BaveQy8T2+VkUCwVSqQT1Ta2msDjKMYXFFHn28Yen1O74OfChM33MOP02Qs3LkWWZVCqF3W5HlmU0TSMYDBIKhSq6jkAggMPhYGRkhJlL3s+Ap45TuYZoMsMdj7/et9PppL+/n76+Pl566c0Pnmq18vi2EbyqTDhTwCgWQNMQVFs5+KuQwxgqz5aqalpx+NNYrCLhHTVE+2YiynrZt0QQ0Up5xgcjlIqdCMUZpMZ20DBbxF9noNj9JAbjeAONDO9HWCAICAhYbbapfdAmRyymsDiIBD1wxdkK3rlfpLbteJLJJG63m1wuRz6fJxgM0t/fj6qqiKJIKBQCYHBwEJ/PR1NTE8ViEZ/vXF6I7eAy63d56tUMgxMZ/tPpNM8//zyRSGSPSlVd14knEty+ZiuulgUUchYMrViOHlMsoJUgl8Rm9+LwqYwPGBRyVUT75mDoAlpBAyTK5dkLeGsEajrTZGP9xAariQ5voq4rw9YXI0RHLTjd+y/JaOg6qVRyl0A7k6OVaeXBeah53yponX8BgbbzyGaz9PX1YRgGsixXygJ6PB5kWaZYLKJpGoIgkEwmKRQK5PN5FEXB6XSy6KSr8M79Ny4/x8ekI2kikaC3t3evqfdlScatKvTF04wnkhjZFGglRKsN0eVFKmUhl8aiOlBUDVmpRy9pGKSxB3pBjAEGCAKipYfmxZuoaspSN6sPb9PzhHts5JIiVvkMQg2nTakimSAIOBzOSmFkk6MXc2ZxkAi44dRlAZqXXovN48VmszF79mxEUcTn81X0FV6vt1LjY3R0lHw+T0dHB1Cu1WEYBtlsFo/HS6j9TC543yD3P/0j1k4hGXUul0XUyhYHAwEkGWQFPREFq6s8YdB18tkk2YQNQciTCjdgsaWIDthQbVXouoEoGBhaE6Pd3WAYOP0yrQucaIUUO1d3YbU7USxixWKyP3RdJzuFRD0mRzbmzOIgsWAGzFn+IQqCrzJjkGWZdDrNwMDrvhiTMw1BEKipqaGxsXG38O9IJEJ3dzf5fB5/sJFQ22mctXzPcX6CICBJEpIkIYoi0fEwqghCYhzBMKBYwOjZgDG4HSObRJ9w4shlE2RTSYY3zSaT0Ji5ai3uukfIpiIICBiGjmA4ifacRt+62cRHCpSKOoGGAgg6VoeXfDpGLrt/r0xRFLGoaiVxrsnRizmzOEg0VVtwNZ5LVirXAgUoFApkMhk8Hg/ZbBZFUXbLdG0YBvl8HlEUsdlsFItFnE4nM2bMQFEURkZGcPs6mN+qI1A2UsqyjN1up6Ghgfr6+oqlJRwO07djGzXVNTgcdtJ6CWQZIxVDcPkREBGCjeXZhp5nbGgrVY2zyOcT5FIatR0y1W0vs+3ZWhR5LgCiYUErBEjHDSRLnsEtYHc2oGslsvFxYpH911YN1tQSqAqxdeOG/bY1ObIxhcVBQAAWzGnCkL3U1dZRLBYrBYOrqqrIZrNkMhlEUSQYDCJJErlcjqGhoYriU5Zl4vE4VqsVq9XK8PAwLpeLbHocr0vBYdOobWijo6ODqqoq3G439fX15PN5stksa9asobe3j/G+bmZ47KyPjSHUtiHUd5QVm4oFweEBqwOKeRLRQXKJCH7vTIa2DLLsfBkEgaFNObLRAloxj6LawbDi8vsx9HGcPjvx/ijJMY1YuI9Mcv+1VRctW0Hvju1vuw6ryeHHXIYcBBQZ2htU+ofKafc2b97Mq6+WCy3n83k0TcPhcGCfKJij6zqyLNPc3ExjYyMul4tkMkljYzlMvmwR8WG320nGx8nkNFSrlbq6OgKBAMFgEFVV2b59O1u2bKG/v5+dO3cyNDTIUw/dz3FtdRhjfVDIITh9kCvXScUdQPCULRjFQoahnvWkIyPIUhO5dImX7smQicxCki1Iiko+myQZzdH/yiyKeQvFTBBJ2kl8pIeBnWv268EpCALHrTqFxx68D107sHwYJkce5sziYCCAVBojGKotF/FpayOXy+HxeCgWi8TjcSwWC3a7vVKlfHR0lPr6eiRJqhzL5XJEo1E0TSMUCpHNZtFS29jcmyORlNiyZQvd3d1omkY2my0f18pVtSb/PvbA3dz0gSu49b4HKTbNAkVF8IYwinlIJ8Dpqwx7uO8V3N4aVLeOYEnQt24JLn/ZH0KSLYiSgmHopCNJ4kMqO56XiA7F2bnl+SkFk9kdThYuXc5PvvPvh+yjN/nHYQqLg0CxBPG8G6fDRjKZJBaLVd7+drudSKQ84/B4PAwNDZFOpykWiySTSbLZLA0NDaiqyuDgIC6XC7fbTSaTIZFIkE8NsqUfiiWNoaH9e5CODA+iJ2PM8lhYn4qBOwCiiCCqGHYXQnULxqbnKdfrKLLttcco5I8h3F2LO6SQiY6hlQoU8xkc3iClQp5UeJC+9TrhkWcZH9k+pZgQgIXHLGdsZIjwXooPmRxdmMLiIGAYsGbDCEtG1iC4F5cL7dhsDA8Po2ka9fX1GIbB1q1baW1tpaamhlKpRDqdxm63V3QV9fX1QFkxWiqVGB0Zxq287pQ1FYqFAo8/eC/vO3EFa+95CqHzWIzoMILLhxEeLCs4JRkmTKzFQobtGx/HojqwO/2oNjeSpEykDdTIZZNk01FymfiUhQSUlyAXfvCjPPLXe9BKUzOxmhzZmDqLg8T9zyTZ8dx/okp5QqEQ1dXVQFn/kEqlKJVKdHR0oKoqhUKBXC6H1+vF6/ViGAYDAwNs3ryZsbExVq9eTSaTweuyEI8MsPYAE3Hdf9cdzOrswjO0CaIjCLIFEhGMHa+gv/pkWeH5Bgr5NLHxPkb6NzDYs5b+HWsY7FlHZLSbbDp6QIICyvVUZsycxd/uvvPABm9yxDKtQtQPBbIso+s64Tj41EHcwnbqZ72XUknD7XYTCASw2+1YLJaKuVQQBOLxchz68PBwJfFvQ0MDmqbh8Xiw2awYqS3ccfut/PWZA7MkpJJJ5i8+htraOl7uGSzHhkSG0J/9M0RH+EfklfjYNZ8hFo3w17/84ZBfy+TQIwhCyZxZHCQM4LePQGn8KQa7n6avr4/BwUGKxSKCIFRqlhaLRURRpLq6GqvVSjabJZ/PVwQFQDKZJBPrpX/rw/zyzi0HPhZD59Yff48zTz4Z/8CraOsfQ3v8DkhG+EcIivrGZk561zn8+mc/MHNvvoMwZxZvk13LAWTykMoWWdg4iuSejzdQh9PpRBRFhoeHWb16NV6vl0gkgsvlQlEUQqEQfr8foOKPYZULZPv/zBdu/BmvbM/v7dL7JBoJ4/J4OGHJYp6/45doqehBud/9oVqtXPeVr/PcE4/yxEN//Ydc0+TQM+0KI/8j2D4IUn4HjeoLFIQAYzGBXD5PVVUVqVQKSZJIp9NIkoTNZmNgYIBEIoHFYsEwDAY338voC5/lx7fcxV+eLAsKi8WCxWKpzDymyoZ1a1h5yhksPGY5Lz331CH3dVBVK9d++d8p5PLc8qP/RJti7IjJkY8pLA4BhgHruiEajTAv8CKeqna29yWpClbT1taGy+Uqe2Zms6xbtw6Xy4Xf76d76wbW3HMNhR0/5pa7w9z+aHnBoCgKHR0dBIPBSrWyYrE4pem9Viqx7qUXOP+SD3PS6Wfz3JOPUsi/tZnK/vD6/HzjR/+N1Wrju//+JbKZ9CG5jsnhwRQWhwjDgK0D8MJraULi/2/v/n2aCOMwgD/v3ZWm0uMaWmkYFFATIYIWlB8SJYIaXR2Ngw5ObA7GTWdNjHExjhonjQuTg42QAlWUQApRokHTVkAjEOz1SgstqQPQaIL2ChWoPp9/4N4b7snd5X2/jx91VUByMY5kSiAWTyK1Mv7KVaphKf4Z02MPEAlcw1R4DLeeAN0/VbFaLBY4nU7YbDaUl5ejpqYGqqrCMIxMjcGfLCTi8Hmfoa6hCZc6r+Dr5ATmY0ZmGvhGCCHg3OlGfVMrbty+h/dvR3Hz+tWshc1UeP6rYuStIgng4B6g3QO01NpQuc+DUocKTS2CtBDEoj6O4JcEuvzAnafA4hpv7quBUV1djYqKCmiahlAohN7e3syGr6zrkGW0nTyLC5c7MTc7g9f9Pgz0dWMyHMy5hlGSZeyqqEJLWwcaW9uglmh4eP8uXvle/JVKR9p6kiQlGBabSJGBSvdycERiQPgbMD4lMBcFlrKUhwgh4HA44PF44Ha7kUgkEAgEEA6Hc/qXYVdLcO78RbSeOAXNUYrBlz74e7x4NzIMXY+sTMla+/olmgMHDjXgWMcZNDS3YnZmGv3dz9H1+BFiRvZqACpcDIs8Wz1+nitZlk0/8DabDWVlZXC5XAgGg78dsZdNkdWKqn370Xy8HfWNR2FXVYwMvcFSKoUdxcWwqxoggKgewbxhoMhqRa3nCKL6dwwN+DHQ14Pgxw+/NLbRv4thkUeKomQOdOVKkiTIsoxkDr0a+WyElxUFuyv3orb+MIrtKko0Ryb0FMUCPTIHQ9cxOjyIidCndd0jFTZJkhJCUZRoKpWyb/ViCt3yWYr1f6/n8nZBtNkURTEkIQS32OXBRn/sMShoOxNCpLndm4hMYVgQkSkMCyIyhWFBRKYwLIjIFIYFEZnCsCAiUxgWRGQKw4KITGFYEJEpDAsiMoVhQUSmSNiM2fBEVPCUdDrttVgsp7d6IUS0faXTae8PYCyFZC+IDU8AAAAASUVORK5CYII="}
,{"background-color":"linear-gradient(180deg, #000000 0%, #000000 100%)","background-pattern":"","items":[{"x":-626,"y":96,"w":2749,"h":510,"type":"text","text":"","text-data":"Qm9udXNmcmFnZQ==","font":"sacramento","color":"rgb(202, 222, 236)","font-size":42,"font-style":"regular","justification":1,"align":1},{"x":-656,"y":602,"w":2803,"h":770,"type":"color","background_color":"linear-gradient(to bottom, rgba(0,0,0,0.423645) 0%, rgba(0,0,0,0.423645) 100%)","border-radius":0},{"x":-611,"y":599,"w":2740,"h":776,"type":"image","image":"png","image-data":"iVBORw0KGgoAAAANSUhEUgAABiwAAAHCCAYAAAB8COEEAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4XuydBXgUyRLHT7AD7nGHu0uQKBLc3fVwDnfncHfncHeH4O4ECAnEPUECwd3d7l7/Q5obJrPZ3WRDsuG/3zcv7ExL9a97eu9VdVX98AM/JEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJGCGBFL89nvK1GnTZ/hJfMxQfIpMAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRgzgRKlq9cffdpr4teN57/i+vcpXuv/16xaZdN0eKlzHlclJ0ESIAESIAESIAESIAESIAESIAESIAEvncCP37vADh+EiABEiAB8yGQJl2GjPucfa9cDPT3cTyyf3fixImT5MpXoFDpClVqJEqcJMn2DauWTh05sNeHD+/fm8+oKCkJkAAJkAAJkAAJkAAJkAAJkAAJkAAJkAAJkAAJkAAJkIBZEWjbre8gz+vP/kmZOk1apeAIDzVhzrJ18LhYsmnPsUSJEic2q4FRWBIgARIgARIgARIgARIgARIgARIgARIgARIgARIgARIgAfMhMGravGVzVm3dq0viP7v2GQijxYyl67ebz6goKQmQAAmQAAmQAAmQAAmQAAmQAAmQAAmQAAmQAAmQAAmQgFkRSJAgYcIfxScyoXsOGjURRotWnXr0M6vBUVgSIAESIAESIAESIAESIAESIAESIAESIAESIAESIAESIIH4QwAGjRXbD51GMu70mTJnjT8j40hIgARIgARIgARIgARIgARIgARIgARIgARIgARIgARIgATMikDOPBYFPK49/YS8FmYlOIUlARIgARIgARIgARIgARIgARIgARIgARIgARIgARIgARKIXwSQx8L96uMP9LKIX/PK0ZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZCAWRGwLVqiNHJZ9Bg0coJZCR7Dwqb47feU+vKAxLAI30XzSZMlS56voJWNsYNNlChx4i79ho7+JWnSZMbW/Z7KZ86WI9f3NF6O9T8CiZP88stvKVOlNgWTHLnz5U+UOEkSU7QVl9tI8XvKVHFZPspGAiRAAiRAAiRAAiRAAiRAAiRAAiRAAnGKQO8hYyaPmjZvmaFC9R0+flq1uo2b6Su/96xvyD5nvyv6yn0vz5G0/EzgzacDRk2eZW5jrtWoWev1+xxdzUXuweOmz9150j3IWHmxrmFoy5Yzd15j634v5S1ti9iDUd4Cltbfy5hNPc7sufNaHHAJCE2fMXMWU7cd0+0t3bLvxIptB09Ft588FgUtXa88fFesVLmK0W0rLtcvaG1XFO9LuSo168ZlOSkbCZAACZAACZAACZAACUgCPxEFCZAACZAACcQ2gRr1/2hh6ClXKHL/7NpnYLO2nXvqk/v4gd3bM2URR7Hz5i+or+z38Dx7rjz5kv/6vxQf3r97Z27jrVC1Vj1zCu+V26KA5ePHDx8YyzlXPouC/3z69OnOrZvXja37vZQvXLx0OYz15fNnz76XMZt6nMVLl6+cIXOWbEnMzJMH+xfmv5AwWiVMmChRdLj0GTZuKtp48/rVq+i0E9frwsAHGc1x34/rbCkfCZAACZAACZAACZBAzBCgwSJmuLJVEiABEiABIwj8+NOPPz1+9OC+IVXy5C9khXJpM2TMpK/8+TMnj6FM0VJl4/UJWn0c5PM8+QuGsfP39jAbTwUpu02xEqWvXrpgtMeCoWxMXS5jlmzZH9y9fcvYdgtaFy56IdDP+/27t2+Nrfu9lIeyWtiC7t++eT30exmzqceJ9+nDh/fvb4ZeDTF12zHZnnUR+5I/iQ9Cp1lYWttFtS+bosVLlapQpQbqv3zx4nlU2zGHevI3M8DH080c5KWMJEACJEACJEACJEACJJCACEiABEiABEggtgkIvdm7H3/48UdD5JCxy3/++We9v2FB/j6eaDNvuJHDkPbjcxkZQifQz8vDnMYJL5lUqdOmO7jTYaM5yP1zggQJ0mfIlOXo7VsOxsj7k1jU1oWLlXBYt2KxMfW+t7KFbAoX8/NyPx/T44ZSHIrtLNlz5hb/TPL44cP7rmcdjz95ZLznTEzLamz71nb2JUIuBAV8/Pjhg7F1Y7M8chPJ/q3sihb383Q7FxV5eg4aNVHWe/3q5YuotGEudbDv37px7eqzp08em4vMlJMESIAESIAESIAESOD7JqBX2fN94+HoSYAESIAEvgUBYa9492uKFL8Z0lcioUVEuZcvnusNB/P08aOHz548fpQ2vX5vDEP6NvcyFoWsbXEy/a6ZhRsqZFs0LKRJoK+nuznMQVphrYDx4c7NG9eMkTdXHosCyUTMG56E1k0ttYCbLkOmzNvWrYxRo07dJi3bImRQytRp0iqlCfb38Wpeo0yUT/Ybsx5iqmyqNOnSI7ya86ljh2Oqj5hq19a+ZJmH9+/e+V+K3363sitWYsMPC2cb21eJshWryrBi4b8l8dbDAvuQ2FYsTx09uNdYTixPAiRAAiRAAiRAAiRAArFFgAaL2CLPfkmABEiABL4QEB4W71Om+loxqA+PoUp3nCpN8ssvSfW19z08tyhoZWuO4aAKWtsWwfyYiyIfCnXIe+tG6FVj1lXO8FwrVy4GBxpT73sqi1P1GK+fd8x5WCBHTt/h46fBk2LZ3GkTQoKD/BMkSpjot99TproQ4Odt7rzN7X2SvOHxAu8apxNHDqRJlyGjMFiErQVjP90GDB+LPDEhl4IDc+crUCg+e1jkzJ0vf2LxAxjo62UWxl5j55LlSYAESIAESIAESIAE4icBGizi57xyVCRAAiRgVgTgLaE+yaxrAFA04dkVoWwyZJBIqPr2zZvXhpSNz2VwohrhtMzFS0E5FwWsbIs8F5anG6FXLpvDHKUTsCHnrevXjDJYZM2RK88/4nPzmnnlFfiWc4L8Ff+KT4C3R4zE47crVrIMPCtg2OvZplFNeGh9y/F9i77wPqEfczNeFrS2KwqjBQyXaYSnTbN2XXrBcPHg3p3bhnJD3gpLYfQ6sHPrBuE8k/5NltevsJ4MrW9u5WSeDxoszG3mKC8JkAAJkAAJkAAJfN8EmHT7+55/jp4ESIAE4gQBnGQWET5SGiLMRxF0HeWC/LzD8lPo+yT5JWlSGC30lYvvzwtY2hbGGM1NcfWj+OQraGUDJaW5KBYzZM6SDbIibrwx6yqbMFjcu33rBkKkGVPveyqLHB+hly8GGxISzlguSOY8dNKshdiPerdtUjs+GivAxKKQjR2MuJcvBPobyyg2y9sVL1UW/fuL/CX+3u6u+Dc8LoyRqUu/oaPxbq6cP3MyfhtevXweb8NBgQv2fYxX7PtmlbfImDllWRIgARIgARIgARIggfhHgAaL+DenHBEJkAAJmB2BJyKxAmL3GyL4TyIoN8oF+/t6GVI+abJkyWNCuWlI33GpTH4rmzCDhb+3Z4ycTI+psWbKmj2nWBop/L3cYjzJsqnGAIPFvTu3br5/9/atMW1irDdCQ8zCi8SYcZmqLOLxF7CyKxJT4aAq1qjbECGCZk0Y/ld8SKyti7tFISvbQD8vD+mtZqr5iel24P0CD6QAHw833/Bk2/C6MLTf0hWr1rQUHjonDu7ZEXIxKEDYK5K9ehm/E27nt7QpfO3K5Ysir3i8NswYugZYjgRIgARIgARIgARIwDwI0GBhHvNEKUmABEggXhOAcjDZr4YZLOzsS5QBjH+Etk0flJ8TJEiABLO3VcmPU4hY9JWEchLGDH1txOZzU8pZ0LpwUSjRHz24dzc2x2Rs30gUjjrmFL4mU5bsOa5fDblk7FgzZ8ue8+b10CuR1UOyYBnSx9j2zb183vyFrJCPxt/LI+x0vak/TVp36Abl7sFdDhtN3XZcaQ9h4ZBjRYTUihGGMTVOGKusixQvFSK8QmBkQHg4eMAY42EhvSuWzpk2HnL+In4A3rx+HW+978AM+6e55P6JqbXDdkmABEiABEiABEiABMyPAA0W5jdnlJgESIAE4h0BoUO/jdjk+pJjI2SLfekKlQEA5fWBSJc+Y2bUuX3zWqgsCyPGhv2n3GYsXb+9TuOWf+prI7aem1rOAuKkbVSV/pgX5FeIDRbWhe1Lot8AH/NJGpstZ+68xhossPhTi7j8kRks6jdr02G5wwHHBet2HIyNuYjtPpG/AjL4e5ve2wZK/KIly1bYvmHVUkM8Dxq3at9l71nfkBJlK1ZVcsF+07X/0DFzVzvsM2SP+tZMzfF9AiPh+GKdLHnyX308XF0kM+xnBaztiiBsnD6O8K6AcQPeFRcD/XxQHvvamzfxN1wgEm6HGfjCw2fpY8TnJEACJEACJEACJEACJBBXCNBgEVdmgnKQAAmQwHdM4M6tG9cx/JSp0qSNDAPCW+CEMMr8KBSD+pDlLWBpjTLKJMYJEiRM+D+RMANxvUOvXLqgr43Yem5KOTNlyZYD3hpRPWk7eNz0uaNnLFgRGyxsihYvdf/u7Vvm4hmCecuYOWv26+KkvjG8UAflb0XiYSET018NuRhsTNvxpSwUzgizJaL5+Jp6TOWr1qqHNpGM2ZC2+42YOENMWc6WHXv0VZZv2LJdZ5zkL1OpWq3/GZiXx5D+TFUG7xPaCvT1dDdVm9+iHTv7z/krfDzOO8v+YLwQ0eJ+M8SYijlBOKnFsyaPkfWRw+JtPPawkOGyorrvf4t5ZR8kQAIkQAIkQAIkQAIkoEUgAbGQAAmQAAmQQGwTuHvrZpjBIk36DBlviyPmuuQpXbFaTfnMkFO1SNaM09IXAny9Zb13Ittsg3KFLYReOSFCJMX22HX1b0o5C9oUDovzHhXFFU6JV6ndoMleh41rvjUrnA5GvH1nx+OHv3XfUe0vS/acuRGKxVhjWKas2XKgT2Fc0xkSatWCWVNOHTmwx1jvjaiOJa7VgwIWuWs+ffz40dSylSxfuTr2CUMNY69fvXiRJEmSXxzWLV+klEUs2WT4fvLwvl0P79+9Y2o5o9uebdESpZHPQGnEjW6b36K+rchfgX683c6dlf35ebqew7+xLhDKS5ccpSpUqQFj1+G927coE42HeVi8jr8eFgVt7IriXbkQ4Pfl9+9bzBX7IAESIAESIAESIAESIIHoEqDBIroEWZ8ESIAESCDaBO7cun4NjaRNnzFTZI1B8QTPCEOMFWjHzr5k2ZBLwYHCRvFa2e6jh/fvRVvob9CAqeSEQg/cAn2MP1WNMDxIiO7p6nzmGwz5qy4sbYvaw2PhYtDnEC7m8CkQntw8NCSi9w7yqYglngXrPE26DBnhLYQT4r+mSPEbkj1jfMMm/b0QJ8GFPQ22osT4E3YlTpT4xx9+/LFH64bVP3x4/94cWJhSRiRIRoibzauXzjdlu2gL4deKlChTfvvGVUsNbXv0gO7tRTShl15uLk7KOuuXzZ/l5+V2LjAOhjDDgsov1idkw35g6FjjQjkk3MZ+qDS0+Hm5n8e7UsimSLHIPGPCvCuE4XrxzEmj5VgQugt7S3zOYYG8RfBGgldSXJhDykACJEACJEACJEACJEAChhKgwcJQUixHAiRAAiQQYwTEIdeXz589fZI+Q6YsujpJlTptOpySDfLz9kDSYX1Gi0SJkySxKWJfcv+OLeuVbeYQSs+nIss3En3rGxAUWh8/fvigr5yxzxGiKWWatOmuCaU2xq1V35RywuiAvsTB6mfGyioV6bERB91GnAaHvJeDg/z1yQ2lM5SSuhSxUHgLvd0bKDj1tRWd5xaFbOxwqlnYeFI0bt2hq6Vgnytv/oLZc+XJB8OPsm3IgtPuYlqeovz79+/eie8vhD3iHYwS4us7/Bv/+CA+P/zw778hF4ICdMmHPAwx4TUE5S6MLQ/u3bkdHTb66kY2hxYFrW3huSKMAef1tWPsc+wnIv9y8mA/b09D6zo7HjukVRbrT+kFoCzzrdagrjFg/4TRQulloKusvvfJUE6mKIe98PdUqdMcF/knlO3h3bkiDNKRJd6GkRvv4B6HDauVRkTx8/AL2norLBaGyBiTPGC4RFgrhL6T3oaGyITfOF3GCMxzXpH3Y9emtdEO5RdTv4OGjJFlSIAESIAESIAESIAESIAESIAESIAESCDWCGw+5OQ1cMzU2boEqN+0dXuvG8//7dhr4HD8lfG5dZUvV6VGHZSrXKt+Y1kGRg6noFvPZi3fuDOygVasXqfB1qMuvqi//YRrQPpMmbOaAgxOyiPZN9rF5Xrl4bvOfYeMUrdtSjmh5HW+cPfluFmLV8t+IMcfbTp1x71mbTv3VBt/wHrB+p2HZq/csmeno0ew5/Vn/8xYsm4brmmL1mwdMmHGfCh4TcFEtlGyXKVqaH/L4bPeizbuPmJRyNoWMoATFP66+oJBZeGGXYfdrz7+4Oh37ZE6CbKshwTJvYeOnSK/I2cB+tl44LQ71lR0x4LwMrUbN29z8FzgNTm/HteefgI/rLfeQ8ZMrvdHq3aQD+NBHhUldyRpRjJ4XXK07tSzP9pFmDOtMsjXgv4s7YoWl89hIOk/atLMQ65BN455XrqDuZbPYIRo2KJtp23Hz/uDW90mLdvq6rtZuy69zl++/0YpL0JfYS2c8r/+eNcpzwsINSTrw/jSc9Coieh3n7PflfyW1naR8TVkDlt16tEP48+cLUeu6M4V3uf+IyfOgPxYc1gDaHvZ1v0n5TrH3wmzl65FAnXl/jH+7yVrIlOQoyySQ2vJGNNrUNlnzjwWBUZOnbt0/T5HV1zV6jRq2q5H/yEYZ9M/O/eIzvsEwxg4KHNHQKHfrnu/wWCK8FrRnSNl/UYiLwjkxhpQt4sxYm2if60+1+45cc7t6qP3MkeMLAMjAdrEOoju2owOD8wJ9i65Z+D3AXuJLpkwTuxXeJ9RZ9PBM54yr5OyDow0eK58r2H0R0L40dPnL0eOFX1zZMjvYLFS5SqOmDJniTLBPORB3iP1GtHXH5+TAAmQAAmQAAmQAAmQAAmQAAmQAAmQQJwi8PeKTbtmLtvw1QlapYBQnu938b8KZRgUMUrFrNZAoCzxCH3yESF3lM+hQIYxQtfg23brOwjtr9l1zBlKl/MhD96aKuG0VDpjnN0GDBt73CvkHvqyKlyshFoeU8mZx6KgJfpo0rpjN/SBk/JQcuEeDBH4qzaajJo2b9mSzXuPT1+81sEp6PZzR9/Qh1B6wpgAdvPXbj9gKoMFFHDoTzKfOHf5+tMBN55A2Q3jEowtMLpozRfC+LhcvPfqgEtAKBSPqAOlsLqssA2kRPvSYAHjAb6D/0mfqw/QD04RR+WFgLJ98PgZ884E3nwqlY5TF67eUrxMhSpqj4rI2j94PvD6pHkrdCZ8rla3cTO0X6lG3YZa7cD4gOcw9OA5EnTDGIF76/aePI95hEED8oIHlPNQ9E5ZsHIT+j536d5rXQwgFxjJfrFe8R0Gt5U7Dp/BOjrsFnwThjD0D6PNUY+LtyfMWbYOfSzeuPuorrEbOoeT56/ciHUYlTlS14ERE2sZBqJVO444gQ3GsueM9yWsIYwFf9fuPu6iNJZJJXBkBguMWcvwFJNrUD0+KPgxnr1OPpdhlMTfMOPZSfegyPZOQ+eiQ6+/hqGdlh27hyUchyELa16ufxgIEPLMFHOFNsBUl5EaRkA80zKKQSmPZ8MmzVqolgVGBjzr/tfwcdFdm1HlAZnx7mw8cMajU5/BI+W+3L7ngKFaMsEoAONsmAFZGDZgrAnb18R+pi4PIyOewTsFz5BsHXud3PexHjDf0f0dhNFXaUjFOpfrDPdh8DfVOmA7JEACJEACJEACJEACJEACJEACJEACJPBNCQwaO20OFDZanSKUChSqKFO0ZNkKUIQoT3Sr60DxCqX3iu2HTqufQeE+ZeGqzVr94NQ92oaxAyfQUQaKoa1HnE2SQwHt4DS6PKmePXdeC3gRqE//ol9TySlPJ0M5hpPfDsfO+eFEPZR5+A7FLBT3WjxgTIDCWd8p5OgsFCjDoYCr36xNB9kOFOJS+bnc4YCjVvtghtP9YAolGcpIJR28F5R1KlSrXR/twbtBGo1weh7rCsYQdXlDxoOY+pAN7ULRjdPl8FpRGg0MaQdl0D/qQWmpqw4MFSiDNaNVBu8GniM/Btbu0i37TsBgV71e4+YoD2ON7AOGDCjspbdCvxETpuOZ5BjhnRGMMUbch8HrmNflu7hgDMM9nGJHfZzmhvIfxgVp0ILyXpeB0Jg5RP8L1u04aChTY8pBob9i28FT+upAMQ2jidwb1OWRnB4cYIBTP4uJNaglr3zfYWSVXgcw2mK+IBsMsMrT8LINY+Zi9srNuz8bCWwKo770fsHpfbnOGjT/s6M+noY+h0EShkstLwqEWoMs0iAr28QeizWO343UadNnUPcF7xDUw5xGd3+JKg/5zkrjDvYjGH7KVq5eW0umsbMWrcJeKd9plMEehD0a4aGUdfAOwogKDnhPzwbfeQEvRnjewBsLY0dfWv0Y+juIttEHfmvl3ODgAfqq1bBpK+khB28sQ+ea5UiABEiABEiABEiABEiABEiABEiABEggzhBo3bnXACigtQRCOBMoWOzsS5WVp5xxgl2X8AhloaXEQqgNhN9AX+q6UOpBcQ+lDk6Ky+dQkuIErClAQZm7ZNOeY/raMqWcY2YuXAmlHRRKMA7AI0EqGiHHvDXb9oOVWuGFZ1KxhdP9+mSOynMYKXSdEJandBFaSKttnDSGYgz5QORzGA3QnjokD0JYQakHrxzM//BJfy+Kiryog3UCgxb6gSIehgSpwEY/UGjry6+i7hvrGu2Vq1Kzri65wAFeDbrahkcMxggDjDScKEPoIDQU+sDJe4RAQtgm2RcUl7iv1XeY0UoouaWXBEL+4AQ93kNZHu+HbBunvpUy4p3CKezozCGYo/3ITsNHdT5h3IRhB14y+trAmoN3kVY5cIdXFOTU8sAw5RrUJSeU0ZgreL2ovZKw5iHb6p1Hz0ZnLlAXRk545eDfCK8FY4LklyFzlmzoRyvUnT6+Ws+lJ4QuLx2sNRhg8U4q60OpDzn6Dh8/TavdPPkLWeG51m8Byhuzv0SVB7wGsR8ZwkUaLNXeFDDuao0Bodjw3uG3ZPdpr4vYT5WGWfwOwNCo7tuY30EYPMEQHjBop1LNeo3wHX/xvU6TFn/K321DxsgyJEACJEACJEACJEACJCAJhJ0e5YcESIAESIAEYpvA3ds3r0OhohVGp0qdBn8gmbCXq/OZVy9fvoCsopxmnHg8a9KmYzckyz6yb8dW5bgKWNoWhgJWJO6NoKj5s2ufgQijM3Fo365IeIx6KJvbooDlpWB/nSGkjOH2/OmTx+kzZdGbD8OUckKxHCgSlZepWK1WjfpNWkwe3r8HEpdLuRMK68znBM9v36rHIhWvfp6uEXgZM26tspjrvsPGTX14/+6dpXOmjleXeRGeINzz/NkIXjIwVsFbYpmod+vGtauybr5CVrZiGYXKNSLvFy5eupy3+3lnnGj283I/P2XUwF5RkR/hgcKMFEIhN2lY/+7Nqpe2RSJgmcjbvlT5Sm7Op0/qSvytq0+Z2PxSkO51BmOLv5e7q6620YbIP+wnUov82mPQyAmuZ0+d2LB84ZecMNlz5smH/l8+f/6sb/tm9ZQJ2HPmtShw61roFS35sooj7DiRHxzg6wXDCrwIls2ZPgEcUR7Gmqw5Pp+gxr1Jw/t3lzKm+D1lKrxTN0OvRAjTZcwcFrC2K4L2A3w8deb4iMp8ok7mbNlzQrkfGXs5TisxB0H+2om5awgFOU77Xwz08/H39nBVy2OqNRjZOGEUgbF1+uhBfZCAXlnWVO8Tkl/DiHD25NEwbxe8w48fPbg/e+LIQfge1dBqusZlE54bxeO8c4R9AHWw1vw83c4pQwRi3+42YPhYJOVetWDWl7w1yj4SJ04c5pEg8tlH2PeMWZvR4YHfA8iqL3wW3r+/xkyZjd9A9V7p6+Hqsm7pvJnKseGdgyEXCep7Dho9UUTnyjygc6tGz589fSLLYd9X7gHyvjG/gzL8nNOJwwew7gaMnDTz8J5tm48f2L09JtZCVN9x1iMBEiABEiABEiABEjA/AjRYmN+cUWISIAESiJcEoIzBwERokmzKAcKAUaZi1ZpH9u7YAuUUlFB4nlRHYluEn7AvXb6y04kjB549efxI2RZOo8KQEej7n8IezxOLY6h//Nmp+5njh/dLRSzuI8QNQuzs27ZprSmgn3c6eQyhSJTJarXaNZWcOEWPGOYX/H29Bo6dOvvU0YN79zhsWK3sM1O2HDmvXw0JC/ej/kBBDYMCjACmGL+yjaZtu/SEQnvxrMlj3r5581rdvojikunTx48fvd3PRTgR3qZrn7+ePn70cNOqJV9OxSNUUuUa9Rrt27bxq7lCaCIYGsA8X0FLm7EDe3RAu8aOB6eJcXJd6GbvNq1W0sZh3fJFSqUw1glkcD17+oSxbYuD8ZbCPvNUF2co1AvZFCnm6+nqotU2ktxCSRns7+PVpmvvvzDmScP6dZOGAyhFEcMedWFQuH/39i3ZDhSu4OMtNMJabefK9znhOdruNXj0JKwVpRJYJAG3xTuKORzRp1NrJVuEb0NdrbaNmcMCVrbhBgsvd2PZ6isvk2qHXAyKNNY+vBcwzgJFoK0AACAASURBVEtBARGMl+ArPQoO7nLYqO7TVGswsrEgRBl4H96zfXOQn0+E0HpYn6jvfs4pQugrY+YCXldox835zEkYyarUbvjHjDFD+r0TCwD3M4QbZNV7r7550PVcrlsYq3WVgdIe84j9BGUat2zfBe/72iXzZgodvabXnvQoE/aKCAaLb8UDvweQV18CbHiipc+YOcuC6eNHaO2Vai7S++m1MO43a9u554Jp40dcEdZMWQ5tYc1ev3r5q33f2N9B7KdyLSAEGPahmeOGf/FeFHatMOO8qdZCVNcQ65EACZAACZAACZAACZgfARoszG/OKDEJkAAJxEsCUomaMUvW7MoBVhEJcqFcOrhra5giUNggwhLv6so7AO8KhAlxWLs8QtgfGAKgzFN7E1SoVqs+QmFsXrX4iwIcyb1xYnmvw8Y1ODVvCug7N69dgXYat2rfJbL2TCVnQZvCRcECngcpU6VJO2XkgJ7KfqFIxUnci4H+mjk6oAT1cnVxMsXYlW1AWQZFGoxP+7ZvDgsnovxA8YVT3EH+Pp6vX716qXwGxSsMUjs3rVkulaQYA0J3Xbt6+eLqRbO/CgGTW8RvBwMo6XZsXL0sNOTShaiM56/RU/6+feNaaPtG1cveCL1yWd1GsdLlKuGe61nH48a2DyXwhQBfb131oBjGXMFLRKuM9NCA0r2ZMAQ5rF2x6NqVyxdlWcwj1je8VY7t37VN2QY8VcBHy5MF5YS9qxD+igPUiaA8njNp1GDpgYT75at+DmO1dsmcGXdu3rimbLtkuUrV8N3r/NfKZmPnsKC1XdEH9+7chvHMWLb6ysODBGVCL18MjqysNJoIg4WfuhwSP0sjJIye6uemWoORydciPAH25tVL5muVsxB7AIxJPioDoLFzka/AZyW1r+d5l469/xoOQ4Ljkf27ZZ/Zwj15boSGRHhH9M2F1nObIvalsN6UhmR1OZ9wY5u12N9hpEUuDSjJNyyf/7euPv/zsPjaYPEtecA7C4ZKfb8H2CsxnsO7t2vmXlKPsZDwqoOxEiHmsCdsWLlojrJMnvwFrfBdve8b+zuYr4CVDYysT588etiuR78h2APwnirXAuQQTnARPKyishZYhwRIgARIgARIgARI4PshQIPF9zPXHCkJkAAJxGkCD+/duwPlRnphsVAKWrdpq3aXLwT6y1PDMDZA0Y3kv+oBwYjRsHnbTlA+upw+ESFuPkK6+GgofUuUq1T10cP79845OR6DYhfx/pHbwU2clh83qFcnU4HDSWBPoeBr2KJd58gSPZtKTkuh7YPs1nbFSqycP3Py3Vs3w+LOy49UpCKMjXqMUNwhHj3kNdX4ZTvWhe1LwiPgqFCeS6ODsg+ZUN1D4zS4fZnylRGGaP+OLeth+ECS4S1HnMOU/d1bNqj25vXrV8q2ZGJoKGtXL5w9NapjEUo+S3cXJ0et0Flos3jpCpXhJaQ0FBjSF7wncFL5QoCfToMFDFh4N7B+tNrMW6BQ2Kn3nMK6gJA8K+bNmKQsJ5P0rtQIj4PwVghpBY8k7bYtrTGuKrUaNAn09XI/cWjvTmU55DfBqe+NKxfPVd7HuJC891JwgJ/ac8TYOUSINPRtCE9jy2QVJ/MfP3xwX9dJfNkePE2gOL8uLF7KPsC7Y6+Bw3EPymflSXZZzlRrUNfYYNAtVb5K9ZtCMay1vyGZOjxEENZLHS7N2LkQHjU2Qj/9ALJUrlm/8dwpY4Yq5cqVzyLMI+fK5QtBxs6FujySUOcVuSYCfbzctfYJWd7f290Vaxjho5BEGwbPVQv/nqoeq7L9/zwsvg4J9S154L2BgQk5hezLVKisxQveEjny5MsPzzgRt08zz4y6HvZ97BfWRexLTh05sJc6PBjyd6COet839ncQ+1aAt4db1doN/hCpMpKqQ1PhncG7r2vPjO76YH0SIAESIAESIAESIIH4S4AGi/g7txwZCZAACZgVAYRqQoxtxNuWgkPJBuX19g2rlioH80BEKUojYgapB9isXddeSLgM5ak61r8INZUdRg6tEEMIfeTv5eHaqfegESKZ7LXm7br0WvL3lLG92/1RB3KZEuTimZNGQ8amf3buodWuKeXESVv0cV+cel2rinOO+1AGaimucE/GhFefyDYFC3ny/ujer3OMyLaLl/2cUF3LuwNzBeMSTowjmeyIKXOWODseO9y8emk7GVZMKaP0PsApcJEn5UZU5e/fsUUD5MzQVR8eFjBwGdt+jlx5LRCKJTjAx0tXXSvbosVxUlor5jzqwMAFJXLpitVqblmzdAH4yLbQdtU6DcNywAhOh5R9wGujlPAkwgl1qYRWy4C2Hz98eL+0CMu2aObE0crnMKQgFM/Jw/t2qcO+FClRpjzCTSlP38u6xswhlO0wnGmFOTKWtVZ5yB96Rb/XDcJm3Qy9GqIOJ1b3j5ZtU6ZOnRbeH8hdoZVjxFRrUNd4hT2yDJIrH92300GrTLHS5SvBi8YU7xNO518QSXGai7323JmTR9VGNOzZMNyojaNRmSuEQYPhS5f3j2wTXlh4P5CYukWHbn0wF5tXL9X0NPnvvUgSlsPig8oIYMzaRP3o8lgnwlbBAN++e78hWowqVK/TAPdFSMSv8jHp4ol5hmcdjLrwptIyOIulbAUDDw4CKNsx5ncQ7yWM2lgLIul3f3i2KQ1EMCbD60jLGB6VtcA6JEACJEACJEACJEACJEACJEACJEACJBArBKCAnjBn2ZcQQcMmzVp47tK91/B6UAqE8D8rth/6KgkrTuM6+oY+POZ56Q6UtOoBIOG0143n/6o9M/Ad93G5X338Af0L20bOmASwdvdxl2Nel+9qJag1pZzHvULuYVzIxaE1HvDVYoKy/UZMmO584e5LKAxNzWLuaod9HqFPPsJwo247TNEm2EAunJRWP9/p6BEs5wtrAMmMI5Nv2db9J1G+bOXqtU09Dtkeclegj9qNm7cxto9aDZu2Ql15Cl+rPt6L4ZNnL9bV9gGXgFDwxLuSKnXadMpyNRv80RLtI6SVuj48L/CsZXg4IfVzGM/wHG1vPHDmS6J2WW7UtHnL8ByeFOq6MCThGU7kR2cOi5UqVxHtlKtSo46xbA0pf9gt+Obo6fOX6yu786R70OyVm7+EPkJ5JBoGe7B1vfLwXbcBw8ZqtRPTa7BNl95/gVGpClVqaPU/bdGarXgOb5rozAXG63b10XusxdMBN54oE13LdrHnLHc44KiPpyHP2/ccMDSycSnbkOsN5RFCSV/7eFdRVhpPZXlj9hdT8eg9ZMzksD0g3ICslH3D/lNuYI19Ud+Y8Bw5i+RvGfI5adXZccItEONUPjP2dxD5UtBP76Fjp+B3F7+/yvakHAjPZYjcLEMCJEACJEACJEACJEACSgIG/ccvkZEACZAACZDAtyCAU9pp0qYL85yAshqK9kMiiSxO7Cr7R9gdhL9R3mvcqkNXJF1F2But8CFWhe1LiOgUVx49uHdXWU96dOwXuRRql7bKhcTBKBeT4123bP4sKJa1kq2aSk6cSkfYJYSJ2bcjYp4IjC+PcFPAaWQ1EzyDMjLIz8tDHU7EFFxyCAW/ONzroxWyBXHXwSYsNnp4vpKv5ytT5gAfT7fWdSrYdxD5JLTCRinLIz8E1o+z4/HDppBdq43iZT57hLg6nTI6fwUU+gj1oiuEDt4DnFTW8gxCn1A0Yq5hWNq1Zd1KpXcFniO/Av4eP7B7u1r2anUbNQ17JmLpa43L0q5YcdxH2ysXzJysLIMT/fDcwOl251Nfs8Xpapx2x3uklZsD+UkMnUOZMyGykFlRnVeMIY3YAAzJa5JGnCYXTipfhVRr1KpdF+w5Z04c3g/lta+n2zktWWJ6DeJ9gmeHVjgovEvlwvOMBPp6RgirZcxcwDAHIytyRQT5eXv6qcYrk7+byhsG3j3wBNAal5qzv5f7edyDF9WOjWuW6VsTiRIlTowyIlLcVx50scEDHoHYZ+s3bd1eKTdYI9ybp8gBAw76xoTnhWwLF8Pf/Tu3rNfKtYNxw6soWOQHUrZn7O9gbosClqhfWhjJNqxYNEcdig/hoPDcVGvBkLGzDAmQAAmQAAmQAAmQQPwhQINF/JlLjoQESIAEzJ4AEmqnFBYLDKRJ647dEGccITPUA0OceCjHpLcETuq379F/CBJ+blu/aokWCCjZfNzOnVU/E5EtUuHewd0Om0wRxsSQSXA8vH83wvtonfo3lZyWtkXDwkEh0bQuowPyMuhSKOHEf6Cvd4RT9YaMT18ZzN2t61c1jUI4LY76WqFEoGzDSV4kQUf4HX39wEMAuUKQCNnUob2UfQuDRWWsSZk4Xp9cyufZRUgoGJXUoYZkGSht8W+ttYv7WC/4C4Xm+mULvvKiQMiWIuIkNORSGzwQDgqny5EbQte6l23fEllzT6iMGvCqSCYyHJ8+dnCvOkY9wkFhjtV1IKexcyiV/dEJ56VrPrLmyJ0HIXS08k4o68BjC3vMo/v/GTsx9s59Bo/cuHLhnPQZMmVBeS0F8bdYg2ANY69WyLBm7bv0AnM8UydFN3YuRLSnMCU1PAFWixwRaq4Im4V7wf7eXynDjXkflGUL2RQuhn1AVyg0ZVkvNxcnfF80Y+IoQ3I9wMCE8sJg8VG2E1s8YDRGeC3174FI55QdRovb4v0zlCFyXqDstnUrND2ykGMEBkgYnJRtGvs7KD3CMmfLmWuLRqL3/9bC14YRQ8fBciRAAiRAAiRAAiRAAt83ARosvu/55+hJgARIIE4RePPm1SucCIahAmE9oGhGbHK1kOJ0aFi8f9tiJUrjL5TcUNotnT11nFaCT5ykFvkarL1FrH51W/8TmhrcE/l0DUpoagpgSN4b6OPpjqTXyvZMKSeUfWgb+QW0ZIYiFUrXS0H+vurnUHSLRyn0KXKjykLYHJKLPMdfebqgrSq1GzSxKVq8FP6NRLu658qw5LMWhaxt0cbZk0cORlVWffWg/IOC/tzpk0f1ldV6jrAtkSXqRoJyeE3o8vqRYXnczp46AcOHsg8YFRBK5sTBvTvUuRVKlK1UFe/ZqaMH9+qSW7a9a9PaFeoT3hXDY+sjTr66fnnhJYN7Wm3/974ZNoc581oUuHIxODAqbPXVQdgalLl6KfIE0TDuoNzr1y9fyjY79x088p9///lHJHKfBhlxX9hLb6r7/BZrULxOvz5UeY5BDnjetOrYs9/n9ymid4WxcyH3K+Q+cDl94oh6rFJJLfJtf5UbQd88aD2HpwMM0sK74KvQf7rawjvUoHxhCySnNqS/nxP8nADlPglLoSwfmzy8hTE9c7YcuZThDJEDBrKJrfKOIWNCGeT9kPlUtOrAqw731fu+sb+Dci3scVi/GrmnIq4Fi4IwNGnlFTJ0LCxHAiRAAiRAAiRAAiTw/RKgweL7nXuOnARIgATiHIGP7z+8x4n4z4ls06TVOsULoYP9fb3evnnzGqF4UK5Vp179cRJ3x6Y1mrHoC1jZFUGYGnWCWLT1WmQ8xV+hu42Q98JUgKDIQ5JSZXs/CkWyyOf9VTgSU8opEq8Ww8l5XeFuZLx0deJVyIiTvfirDBUFAweUiKZg8l4Yh2CcUbYFA8nAMVNmY15xXytE0utXL8LnKmKOEi258hW0DMuf4OZ85qQp5NZqo6C1XVEYfs6dOWG0wQKn+zNlzZZD62S+7AtGA611K58XFknI8e9Du7dtUssn8z4c1TAqlK5UrRbKOzse/SoRt2wDnizCxmcX1vaebZuVbePUd8nylathrpxOHo1gDELbSCSMZN5qmYydw3QZM2W5dvXyxZiYv5x58uaH8RDhxyJrP7HYHPD83du3b/AXRoiWHbr3nT9l7DCMM1OWbDmEzvaxVii6b7EGRUSxt0nEhKnHMHTCrAXyntDnB0V3LmTycIe1KxZp8cLpfRi2xHR9lR8hKnOH9wr1tJJG62rPkNBesu7P4gcB/1buwcauzajygCEGYZmU48DvAdgpveGwP6DML6q9Evey58qTT52PCR4iSAJ+/ozjMa3k76j3377/tVHJmN9ByCWNU1vXLF+ovRbyF4wpQ2NU1hPrkAAJkAAJkAAJkAAJmBcBGizMa74oLQmQAAnEawJQHsKw0KHngGGuTo7HZZgP9aAR3sdVnCivLJLIdus/bCxOQE8fM6SvrtBHdsVKlkGMbS3l/PWrIZfQvtrbAUrIQWOnzdGVyNaYiUBy6JnLNuyQCigkLIWi2c3l9FeKdFPJiVP1+QvZ2EWW3wGhdjAG9al83JPKvF+SJg87WY7wH5sOOXk2b9+1tzHj1lUWXjMwNsk48pjzCXOWrkU+Acwr6t29deOrfAG4h3wJOD2sniuE62knQoK17dZ3kLJPKOdgdEGoMFPIrdVG8dIVKmM96suloVUXhg6Epnks3E20nuMZQnv5hcfnV5eBUaGAlW0RhMBR56HAWrMuUrwU8oBo5b+wEZ4beN9g/NPq27ZoidKYF4TeUq8RxNWH7M6njh1WK+mhREXSeoSc0QpzZewciqn935NHDx/ExPwhHBfCJOnLD/BGCC37h+Fx6sLVWy4G+fvs3rp+Fe4LW9tv90WCCy0Zv8UaxPsE5lKJDDn+7NpnIHLknBf7qKneJ+QlwHwf2Lllg9ZY0f9zYbjR8nIzdv7yW9kURh0vV+czxtY1pLzci0XqiC8eFsauzajyGDZp1sLVO4+ehbEdsqZOmz5DwxZ/doKBD++klP9G6GePKbtwo6S8j++bDzl51Wv6OT+N/OC9hDHR3eWMoy4GKIM5VO+JxvwOps+UOSt+c2FI1fLCgwzIuxOVEHmGzB3LkAAJkAAJkAAJkAAJxH8CYaeL+CEBEiABEiCBuEBAKmvSZ8ycZXD3tmEJgXV9juzbsRUxvxu37tAVYWkiU9Lktshf6NnTx4+h0Ea4mjb1KoXF/ccHp3KRx+FPEVYKSnKcGkeS2poN/mgJBRYSGUeXzamjB/YggfiSzXuPI8mrfalylXCqe/3S+bOUbZtKTihiocwOiiSWvIxHr06WCnmgvMIJ3ZYdu/fFSWCE5xLODc/XLJ4zPbosUH/fto1rB4+fMW/u6q37xOl/hxr1m7QoXLx0uYO7HDYG+Xp5YF6FziuhVl8HhScBTrfDQIGEzggL1rhl+y7wzBk7sGdHZR0YZbzdI57yN8UYZBv2ZcpXRrJlrBVj203+v/+lQB2t5OK4D+8LeKJAIb7xwBmPxbMmjj597NA+2Q/Cv8Co4Hhg/251YnqEmoIhZ/+O/bu1DHlIIn3rWugVXbk9rIvYl0Q/+7dvWqcelwxzhJBt6mdp06fPGPZeRXLK3pg5FPrvRwg/derIgT058uTLjzW5f8eW9Svnf50E3Fj2KI9T6rpCbSnbQ8gbeFD80aZjd4Sfg2Gtf8cWDeQpdpyOfyk8LbRk+BZrcP/2zetgoJi9cvPutSLnTwFr2yJI4AzPnTWLZk+Dp0103yesQ5GqI9tusR/qyikBg4WutWzs/OQrYGWDvVmXMc/Y9nSVFwaLT8pnhq7N6PBwPLJ/N9b08q0HHEOvXLqAkHIwTg7s2qaJUhYYW5HQHrlmhkyYMf+0CN+W38q2cKfeA0dgve3ZumG1sjw89PBd2NJ05hCB8Vl6sSnrGvM7KEOpbV27TNO7Ar8ZMFqYai2Yaq7ZDgmQAAmQAAmQAAmQAAmQAAmQAAmQAAkYTaDX4NGTvG48/3fElDmaibOVDSL+/mG34JuHXINuIO9FZJ31Hjp2Cto95X/9cfV6jZury+LEqvOFuy9RBpdT0O3nUKirQ24YPaDwClA4r9h28BTaPhN48+n4v5esUYeIQlFTyVmpRt2G6EtrrHIMM5as2+Zx7ekn5KvQGlf/kRNnSB5QliO+elTHr64Hz4qVOw6fke17Xn/2z5iZC1cifjs8BnAfBh6t/nAqea+Tz2VZ1yP0yce/V2zald/yc/gi+YGyHu1GxiC644HS0vXKw3edRPLlqLSVPXdeC4xD5u1Qt4EwWedDHrxFmQXrdx7COlKW6dR70AiMP7/l59Poyg+8eFBP5ppQP9/n7Hdl0rwVmiflUXbJpj3H8H6pQ3fhWbcBw8a6XX30Xp4QV7aNvAnot2GLtp10MTF0DlG/frM2HTBGOd+7T3tdlAaTqDCXdXDC3uXivVdQBBvSjnw38f5CgaysM3Hu8vXuVx9/yFfQKiwE2bdcg7KvfiMmTJeM8BfvF95ZKI5PB9x4Mm7W4tVa4zR0LrDHHjwfeB2h4bTagcId+0lka8oQzrLM3rO+IdiDjaljTNkmrTt2g7xS+S7rfgseWHuDx02fi/0J7xHeNZnEWj0GKP/xHirndu3u4y7wYFCXlW3CoKbFAv2e9Ln6YKejh2bILkN/B/H7gvUFY6lWP/ZlKlTWtwcYM1csSwIkQAIkQAIkQAIkQAIkQAIkQAIkQAKxRgDKmUYt23XWpQhRCwaFnD5jBepA6YoQRPA60DW4FL+nTCXi8ldHWKbIykUHDpKoRjY2U8kJ+S1ti9gjNJQueeGRkFO4WUQ2HijMkcw8OmPWVReyQVGPeVEbTXCKXiac1aoP5ShOJZcoW7GqltIcdaCohdJchn6JiTFAQQ1FtTIUjzH9IGE31lxkdRBSSMbKV5fD6f1ipctX0qqPtuG1omv8YXlVxJrX1XfpilVrwgNB6znWhcwxoPUc84r+IxuXIXMo60MBixBV6rj/xrBWl8XYoFRt1q5LL0PawXrFfCMUlro8ZJu1fONO9V70LdagUhbMKcJAwRCmvF9JhM7TMmrJMsbMRWSsECoI+4ohPPWVgfJci7W+eoY+xxrGHhLV/cWQfvTxgFFVJnSPrD3s5+Wr1qpXq1Gz1mrDrLIe9lF9ezpCHeoyaKAtU/wOYs/BGsS6MoQTy5AACZAACZAACZAACZAACZAACZAACZAACZAACZiIQGRKfxN1wWZigEC1uo2bwWABo1cMNM8mSYAESIAESIAESIAESIAESIAEokiASbejCI7VSIAESIAESIAESOCZyLFACuZHQJ5UvxQc6Gd+0lNiEiABEiABEiABEiABEiABEoi/BGiwiL9zy5GRAAmQAAmQAAmQAAloEChWqnylJ48ePnh4/+4dAiIBEiABEiABEiABEiABEiABEog7BGiwiDtzQUlIgARIgARIgARIgARimADyo1gUsrL1cnNxiuGu2DwJkAAJkAAJkAAJkAAJkAAJkICRBGiwMBIYi5MACZAACZAACZAACZgvgTIVq9VCYmBXp1PHzXcUlJwESIAESIAESIAESIAESIAESIAESIAESIAESIAESIAESMCsCWw8cMbD49rTT2nTZ8xk1gOh8CRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAiRAAuZJwM6+VFmvG8//nb92+wHzHAGlJgESIAESIAESIAESIAESIAESIAESIAESIAESIAESIAESMGsCP4nP6p1Hz8JgUaREmfJmPRgKTwIkQAIkQAIkQAIkQAIkQAIkQAIkQAIkQAIkQAIkQAIkYJ4Eug0YNhbGitkrN+82zxFQahIgARIgARIgARIgARIgARIgARIgARIgARIgARIgARIggThHoFyVmnW3HnXxLVu5eu3IhEOC7c59h4yCseKI+4VbqdOmzxDnBkOBSIAESIAESIAESIAESIAESIAESIAESIAESIAESIAESIAEzJNAzjwWBU76XH0AQ8T0xWsdrAoXK5EgQcKEcjTJkif/tXKt+o3X73N0RZnjXiH38uQvZGWeo6XUJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACJEACcZZAmnQZMk6YvXStR+iTjzBKuF199P6E95X7pwNuPMF3XJ7Xn/0zY8m6bfSsiLPTSMFIgARIgARIgARIgARIgARI4AuBH8mCBEiABEiABEiABEiABMyZQPqMmbOUr1arfgFL28IpU6dJ+1F8njx++OCCv4/XmeOH99+6ce2qOY+PspMACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAACZAAvMfQuwAAIABJREFUCZAACZAACZAACZAACZDA90Lg5+9loBwnCZAACZAACZBA3CGQOMkvv/z6vxS/vX3z5nV0pcqRO1/+169evfz06ePH6LbF+iRAArFP4EfxSZchU+ZXL188j640qdKkS580WfLkb16/ehndtlg/egRS/PZ7SrtiJcsUti9VNm+BQtbJxY/Aw/v37vzzz6dP0WuZtUmABEiABEiABEiABEiABEiABEiABEiABGKcQK1GzVqv3+foGuMdxUIHS7fsO7Fi28FT0e06j0VBS9crD98VK1WuYnTb+lb1s+fOa3HAJSA0fcbMWUzVJ5Syjn7XHpUsX7m6qdpkO3GbwM8JEiTYfMjJq1LNeo3itqTGS9e575BR5y7de/1L0qTJjK/9Xw0YRvc5+13p/tfwcdFph3WjR8C6iH3J+Wu3H/AIffLR68bzf5XXUY+Lt+s0afFn9HpgbRIgARIgARIgARIggfhEIEF8GgzHQgIkQAIkQALxiUCFqrXqpc+UOWt8GhPGglO1hYuXLvfx44cPCRMmSvThw/v3UR1jn2HjpqINcXr6VVTb+Nb1ipcuXzlD5izZkkRTGauU27pwsRI4vfxJuJl86/Gwv9ghkCNXXot8Ba1sfk+VOk3sSBBzvZavWrMujA0FrOyKeJxzirJhs3m7Lr0yZcmW483r12azP8Qc1W/fcqLESZL8NXrSrCatO3a7ffN66OpFs6f5erq63L1968a/4pOvoKVN5z6DR46duWjVTz/+9NPuretXfXsp2SMJkAAJkAAJkAAJkAAJkAAJkAAJkAAJkIBBBI55Xb67bOv+kwYVNqNCpSpUqSFP2FraFS0eVdFtihYvJdtBWKiotvOt601ZuGozvEISJEiY0FR9dxswbCxYpE6bPoOp2mQ7cZtA49YdumLOYfyL25IaJ13SZMmSy5P47Xr0H2Jc7f9KJxOWUXgdgREU5lFth/WiRgBhvWYsWbfN/erjD6079xoAjyCtloRdKik8hTBXmLOo9cZaJEACJEACJEACJEAC8YkAPSzi02xyLCRAAiRAAjFGIFGixImhIM+SPWdu8c8kjx8+vO961vH4k0cPH8REpzgVnCp12nQHdzpsjIn2Y7NN26IlSsv+rYTBws/T7VxU5Ok5aNREWU+Ep38RlTZio461nX2JkAtBAfAwMVX/OGn//NnTJw/v371jqjbZjuEEoJzFHOQrYGmT7Ndf//fqxYvnPh7nnUNDLl0wvBXjSlrbFSuBU+oXAny9jasZt0tbiXH99PPPYXn2sD9EVdo2XXoNgNcR6r8WExLVdlgvagTKVKpWC+HKxg/u3XnHxtXLdLWCPEZzJo0avHDDrsM1GzRt6bBu+aKo9chaJEACJEACJEACJEAC8YUADRbxZSY5DhIgARIggRgjULdJy7YIPZQydZq0yk6C/X28mtcoYxcTHReyLWqPdgN9Pd1jov3YbNPWvmQZKNZFzu3foZzc8MPC2cbKU6JsxarKk+UiN2+0k/MaK0NUyiPXBMJ8OZ86djgq9XXVyVfAyuZycICfKdtkW4YRgJfQyKlzlyKfirLGP+JT3jJbqhfCkmRYS8aVKmRbxP5G6JXLYu0/M65m3C5tJ/YHSHjrxrWrUfXASvF7ylQtO/bsJ0f6UhiQ4vao4590lWvWb3zn5o1rOzetWa5vdK7Op0/AcIG5p8FCHy0+JwESIAESIAESIIH4T4AGi/g/xxwhCZAACZBANAj82bXPwL7Dx0+DJ8WyudMmhAQH+SdIlDCROLib6kKAX4ydbC5obVsEYgf4eLpFQ/w4VxWeKoVsChdzOnHkQJp0GTIKg0WUTlB3GzB87D8iYUPIpeDA3PkKFDIXD4uYmNffUqZKDSPIqWMH9sa5CY/nAtnZlyq7aMPOwyL8/k84Re7l5uIkHGc+pPgtZcrXr1/ClhAjxgqEzsmWM3feQ7u3bYpviMEU3kJH9+10aNut7yB4m8F4Ycw4sW8nS578VxiVLQpZ2woHLBosjAFogrLpMmbKcvlCoD+8gPQ19+njx493bl6/lipN2vT6yvI5CZAACZAACZAACZBA/CdAg0X8n2OOkARIgARIIIoE7IqVLAPPCn9vD9eebRrVfPbk8aMoNmV0tQJWtkWgtMMJaqMrx+EKBa3tisJoAUOM0E1laCaS4sJw8eDenduGio0cGDh5fWDn1g3C6SX9myyvXxmiFDO0/Zgsh3lF+1hTpupHRCEqjLYuBvr7mKpNtqOfAMINTVu8ZusrYZfo0bpB9SA/H0/9tUxTIr+ljR3CUPl7u5tsHZlGsui1kjBhokQwaIq8zGf8vdzPozUrkVDeGIMFDHjN2nbpidP9p44e2BNusGBIqOhNjdG13wgrcsbMWbMbWvH9+3fvdOW5MLQNcy23ol2YU9GP4vop/K/8/+ifxPePHVad0Wv0MdexU24SIAESIAESIAES0CKA/yjihwRIgARIgARIQEVAHJj+aeikWQvhWdG7bZPa39JYIePhQ6lvLop4QxeQXfFSZVEWykipbIWC0tD6KNel39DR4LJy/szJSX5JmvTVS/MIBwXZLQrZ2CH0CU4eGzPmyMrmt7INM1jgNLmp2mQ7+gl0HzhifEpxJHxw97ZNv6WxApLlL2QdForOlIYv/SOO+RIFhGdZYpGF2d/LTewPn416hWyKGLU/wLtCbAvJVi+aPQ0GELRBD4uYnzt1D65nT53ILcKkwYBkSO+p06XPgNwvhpSNL2VgqBAXjBM5xVVLXNbiqigueE5tE9dcceURZRKLCwYNfkiABEiABEiABEjguyBAD4vvYpo5SBIgARIgAWMJVKxRtyFCDY3o27lNTCXW1iVTpqzZc4qILymgtDNW7rheHl4riO0f4OPhllIkFYe88Lo4eXjfLkNkL12xak1LEbv/+IHd20MuBgVAMYkT7obUjQtlLApZ2Qb6eXkgnJWp5AE/hFS5HBzIHBamgqqnHXgFNWj+Z8fdW9evcnM+ffIbdfulm3wizBGStgf7+8YrIxX2BwzS19Pt3L07t27ev3v7Fta3oXx/T5U6TdM/O/dAvV2b165AOD/UNac9wtCxxvVym1cvnf/44YP779+9fatP1szZcuRKJX4PQkMuBusrG8+eJxbjgZGinrjqi+ujuKxUY6wsvu8Q1zxx3Yxn4+dwSIAESIAESIAESECTAD0suDBIgARIgARIQINAk9Ydul27cvniwV0OG781IIQwQZ/x7fT0Tz///LN1keKlQoR3ARSICHcFzxVjPCykd8XSOdPGg9EvSZMle/P69atvPUdR6Q8njdNlyJQ5wIThoCCHCA9U+JJIuI2QKlGRy5R1EPIKikdTthkX26rfrE2Hn0TiiuVzpk2IDflg+LoUFOBriDI4NuSLap/IXwHvKT9hsEAbfsITC2M1NFSQ9K5YtfDvqXgfYNBEO2/fvDKLPSKq3OJiPRhlkWPl9atXL/XJV0kcEEAZZ8djh/WVjQ/Pwz0r4DGRVFw9xNVcXAXEBWPFP6ox5hbfB4lruqiXPD6Mn2MgARIgARIgARIgAX0EaLDQR4jPSYAESIAEvjsCUCoXLVm2wvYNq5aa8iS8oSCtC9uXRNkAHy93Q+uYQznhsGKNRLg+Hq4uUl4YZQpY2xVBGCx9Y4B3BYwbJw7u2XEx0C8sX4OIHpP0jZkoI2NiXnGiPH3GzFniQnJ2KIfX7D7mvPesbwhyk+ibT3N+Xqdx8zZnHY8dMia3gqnGK5yvfsuRO19+Mefxan9AGD7rIvYlYSgW6XsegxdCxyFEFLzd9PHDu/BHm07d4V2xY8PqpZ/3h6RQCP9gLkZNfWOMj88TJEiYsHn7rr3v3rp53ePc2VPxcYzKMSnyVaQR95eJq424coSXeSP+LhdXH3ENFRdCQt0Pf4bfyLDwf/yQAAmQAAmQAAmQQHwnQINFfJ9hjo8ESIAESMBoAuWr1kJ4hh+Q1NnoyiaoYFO0eCko3R49uHfXBM3FmSZwehrC+Hicd5ZCwXgBBWzWHLny6BMU3hUIJ7V41uQxsiwUkm/NxMMC8wq5A31Np2iWuQzigsECSuF+HZrXf/ni2bPB46bPRY4HfXNqjs9z5c1fMEv2nLkP7NiyPjbkRxJqKPcDfeOXQTNP/kJW2AuU+4NvuHHTEC8s6V2xYt7MSdLbCAZNeKFg34iNuWKf+gk0atmuMw4JzJs6ZtiHD+/f668RL0ogFNQkcTUKH81R8XeBuLqIa5a44Nk5VVz9xAUjBTy5EC4rf3jOi3gBgYMgARIgARIgARIgAV0EaLDg2iABEiABEiABFYGS5StXvxDg6x0bBgMo2BACJb7Fpgdi2/D49N5u585K5H6ermGhX/TFqS9VoUoNKC2P7t/poExYHeZhIWKOmMMiti1aojSS/968djXEVPIilwHawkl0U7UZnXacThw50KhisYKY4w49/xqGE/PRaS8u1sX+AM8rl9PHj8SGfFhH6De+JVm3LVYiLH+Fcn8IEEYZ5GfRtz8g3Bq8K3BKf+emNTihHvaBQZPeFbGxSg3rE+HjegwaOeHovp0OsXVAwDBJTV7qN9GiNFag8QBxzRfXIXFlFheMFAnFBa8KeF/kD/+OexmE0SKTuH5nIm6TzwsbJAESIAESIAESiCMEaLCIIxNBMUiABEiABOIGAcRKL1KiTHk3lzPfPJEuCFjaFrVHiIyLQZ9DHsWnDxLqPnp4/55SYY8Y9Tj9XMimSLHIxhrmXSGUxItnThoty+GUOViZg0IyUaLEifNbiVwTQQF+iNFvqnm1KGhlixjxSEBuqjaj286L58+eDu3ZvjmSQrfs0L1vdNuLa/WLl6lQWaRh8RHDfBIbsgnFfmm8CyEXgvxjo/+Y6rNI8dLl0La3+38GzXdv37y5GOTvo8/DQnpXLJ0zdbzylL547ZKYw/4QU0zjertDJ81aiPBf4wb16hTXZTWxfPgNUCYjDxLfEQ4ql7hSigvGu27ighcGPLlg3LAX1zVxZQwv9z/xl/9f3sQTw+ZIgARIgARIgATiBgH+R07cmAdKQQIkQAIkEEcIIGmwyOOcPNjP2zM2RLIJPz19OVi/MhLGlchyP8D7IMVvv0P5EesfxNxHjHnl6WkIBY+DK5eCAyNTSMK7wtK2iP2+HZvXhYZcuiAHkzhJkl/w77dCIxnrA9QjAMYHo4XSO8QUMiNBO0JMxbWQN3dv37xx8tDenWUrV69tSH4SU7D4Fm3gncM7GuwfO/tDwoSJEsHb4LpIWK8vyTq4R5asGga/NOkyQPkZJz42whDz7MnjR9cU7zgEQ9g4hOHCfqYlKLwrmv7ZuccNwWSPw4bVyjJii/glJveHZMl/hdLYoA94I+wVfmOwFxhUyQwKZcqSLYelXdHiIprX78aIi8T12B8GdW3zh/gZeGZM3XhQFp4S6RXjWCL+jbBQME5sFddwcc0WF5JtZxUXvAhh0PggLnhnIMcL7jHUWTxYDBwCCZAACZAACZBARAIJCIUESIAESIAEzIUAEq/iJG2GzFmybV69dP6x/bu2acneqlOPfm/fvn2zbd2KxbrGhuTPr16+fJE+U+asLdp36y0SF2eFQiljlmzZUadB8z87Vqxep4GsLw76vl42d9oEJIQ1Fa+S5SpVa9iibSfEw38sXA/mTBo1WOY5uBwc4KerH3DoP2rSzGIly1YUQ3g+tEe75i6nT0QITzNhzrJ1vwjrS49WDarLtsTp8Cqd+g4ema+ApXWQMMoM69Wx5YN7d27jOeSAJwOUSJeC/H2Rj8BUp8jt7EuGh3txcVKPC3Hqazdq1hrKVYR/UT+HTDitv2TW5LHKZ0jGi+9iaiINCYV2MZ9VatZrnCptuvQXxen4vyeMGCjHrWwTsdR7Dho1EXN9/WrIJTxD/Tadew3Ib2lTeNeWdSudRbLlyNZAzjwWBVp27N43X0ErG5Rbt2TezIxZs4UlVb0cHKhzXo1dVzCsYc5OCMMA6kIR2rZb30EwDEFxu9dh4xplm32GjZtaWOQREa/GG4H5w7+wcoR//hVfxKH9T/if806Ox7atX7kEiefLValZd8bYIYijHuFTvV7j5mUqVa81vHfHVlrPvd3PO1er27gZFMpPHj18YOz4jC0Pb5smbTp0Qw6aB3fv3Jo8YkBPGMTU7WBcVes0bDpxaN+uuvoAW5zMTygUy5j7XPnyF0worAV4n/AMeSRmLFn3Zf8Bu73bNq5BSCxj5dZVHtxaiGTEhYXHF3I7OB7ZvxtrD+s+sv0BRkrMNdgnSJgg4bLZ08Yvnzd9orqfP/4UG+Xw8dOK50mXVHr9YD31Gjx6kr3wIsGcjf2rRwcvt8/vrNDNp8D6qi0SjmP9DOzSqrFwBDOJYTdbztx5ER7o1NEDe9QeSL4e512ate3cM38hGzspi3Is0rti8axJY9T7B4ya+vYHZVt4d9AeDKTuLmccFyk8utT8wGHUtHnLKljlSIN1Bu5d+w8bI/bw0mJLvYn9/OrlCzg5/wN+Z+av3X4Ahhd8fyo2/FH9u7Y9c/zwflOtF3U7ho7FmPdBOTcwnk1esHJTpRp1G6JveLYsnztj4tLZU8bpGxOMHAPHTJ0NvuJ3yENf+Xj4HAYaeMWFrYfwj648Tk/Fc+wryGtxWVyPxPWsw6ozn+IhFw6JBEiABEiABEiABMII0MOCC4EESIAESMAsCDRu3aHrxoOnPaAkKixChwydMBMJKiN8oLTs2n/4WGGP0HnyFcrrM4G3nkHxiFBE9qXLV86UNXuOVGnSpc+aI3deKF6guC4klFY4OYq/SAqNtk0BCwpwKLoWrN95CCechU7LH6emZ6/cvMdaKEKhKL0achEJNiN8EK5q3d6T57PnzJNv48pFc3B6eNjk2Yu0yloJ2T+8f/dOPoPSb+GGXYdzCYW6CMt0BW0NGjt1Dp7Xati01dYjLj5Cn2blcc7pFBJkIya8KcaLNmT+Ci9XbYNFIqFZRN/q/spUqlYLykPEpb9983qo8rmI9pIE3yM7QQ2l7+qdR88On/T3IhijoIStWrvBH3+v2LRL6+Q/1hcu9Iu2UWbS3OUbeg8dO6VK7QZN5qzasieyU+lIILv5sJNXsVLlKl65GBwIJeak+Ss21m3c4k+0F+jnZTLlXF5hdIJ8/t4erpVr1W+8Zvcx5xLlKlUFr3GzFq+WY5DMYPRBiJzkv6ZIAcXjC5Ec+5PQ8OLkOtY+1gPa+T1l6jSoA8U/DC9QJmutgzqNW7SpUb9JC12n+BEaCvWMOYUe1fWWOm36DCt3HD4zaOy0OWBfSxjAajVspmlIgdI9Q6YsOLWs+YHXyhH3i7dKV6xaM33GTFkq1qjTAAzQhzBcFEIlGA0KWhcuiv0BFwwaSYUVNKryq+uhTYejLr7N2nXthbwMb0TYr069B40YMWUOTmKLdaSt5E0rBMb+UL1ek+b7tm9ce8Hf16vbX8PHwcir7sPKrljxD2Kzk0poGGE2HTzjUb5arXoIMYY9b8rCVZuhmAYTh6PnfOs1bdXO3cXJMU3adBn6DB2HpMAm+ejbH9CJlheWWKpp4V0Bz6VDu7dtUguDPUIYLAzywIKxGMxhsMD+17nvkFEwPuoaYEEruyI/i8UPUx8MPZsPn/VuKvZY5M2A0bdclRp1ZN0h42fOxxravGrJvE0rF8+FAWrKgtVhbE0CUNWIMWMx5n1QdoPfExgrYDCFkUJsJ0+7DRg2FutI35hGTZ+/HEbxNYtmT9NXNp4+h5Ed4Z7Uhlx4UGC9Ivk4LnhSnBYX/nvnuDBSXBLXYxor4umq4LBIgARIgARIgARIgARIgARIgATMh0C7Hv2HeN14/u/es74hUCKK09F/4PvEucvXq8OEIMkvniH0htYIobg7d+ne6z1nvMNOz6s/e518Lq/YdvBUTNKZNG/FBs/rz/5BSAzZD5Q8kBvXcocDjlr9CyeQ7Kf8rz/eesTZR4Z6atauSy/UUYfjwHfch2EEbRUrXb6Sx7Wnn1btOOKEZ1C44vlJn6sPGrdq38X96uMPbbr0/gsKcKFvS4Zng8dNn2sqDgdcAkKdL9x9qaXczp4rTz7016R1R8Ts/vKBLFuEEhDzBWWxWhYoVFGvQ6+/hmnJib7W7j7ugrGhbWmgaC1OzKMePBLU9YTRaDeewZsCz+Ctg+9d+w8dA6MF/g2Dl1Z/MFbg+egZC1bIcUIxeczr8l3cPx/y4K0pQ8FgTGi3RNmKVc9fvv8GRhjMHYxfuA/jlKHzB5ZOQbeezVm1da/kVKdJiz/RDt43dTswMLlcvPcKz2Hc0+oHimQ8h1LZUDmiUg79430OW7PjZ8wT3lJZhOLdc8cJt0B4GSjbhNER67C58FzQ6gteVluF0hrvCtpRlxktFK1uVx+9jylFM/qDcQAybjxw2h2n5HEPc7Jg3Y6Dco+AcUktG8YGY4VT0O3naAPP81gUtEQdpbeYrId9RO6DMFhhneJCHZRZu+fEOdSt26RlW7Q5ef7KjTDy4tmG/afcwCkq86VVBwY29AVDjdbzY56X7kxduHqL+hn2KNSrUK12fa16R9wv3Fq0cbfe5OgwcmE9nw2+8wKKeLHV5sS+gb1Y128J9qY1u445Yy/G/oa9FO1AjhS/p0wl3yM8h4wjp85dKmWEon/G0vXbTcVP2Y4xY4nO+4D1s+uU5wU5zuy581rACI/fqcjGhbGHzbUwrMbE+ON6myJR9g/h1//E39HichfXU3G9FtcDcT0W10FxOYhrhLiKikszHFpcHyvlIwESIAESIAESIAESIAESIAESIIF4SQBhZ6DcgPJMKukRrgT3oPTHCXrlwNv3HDAUSicoHrWAQIGPujhVqn4O5Y1H6JOPUHrGFEwYKdB/7yFjJqv72HnSPQjPEJJIq38ooDE2hNOQz9t17zcYdRDiSlkHCa5xv2OvgcNh1Nnv4n8VSjVp2EB5PMd4oZiDh4Wsj3wTkRkCjGUDhTLaW7xxN2J0R/hA4eXod+3R+L+XfBXCSM59XxG2RqseFIloFwYIrecIbSMVrsrnMEbgPsJxqesdcg26cfB84HXcRxgXKI7leoCxC/Vw8lpdDyexYZDAKf+ffv75Z+VzeHegHjw9jGUXWfkhE2bMhyIXfcIwI5Xo4AnlK5SJhvSH9eFw7JzfYbfgm8r3CUpvyI2QXOp24L0hlee68o/A2wHGJl3voiGy6SsD2WGcgIEBnjGyPAxzYQYMldFNGgZ1yVyzwR8tUQ/he7T6XrH90Gmw0idXVJ/DELT7tNdFvA9qT55qdRo1hWx4X7XyOWDvw3N4Asn+oRTGPeVpfzyDQQ3rVb6T0xat2QpDjFKJvPHAGQ/Udb3y8B2U7UqPpONeIfcMMQQYygHGaKxZXV5sM5dt2HHwXCASDn/54H2EbDDS6OoHBl4Y4SKTA4p2GOtgcJBh3DAP2BsxfhnySNkGDEn4/cG7MX3xWgfMlwz3pO4rv6W1HdqBh4yhPKJaztixROd9gBFryaY9x4yVFesKxlVj68XH8sIQkUBcucVVQ1z7xXVXXHfEtVBc+cUFowYjIsTHyeeYSIAESIAESIAEIiXAHBZcICRAAiRAAnGWABTLY8RpdYT7QB4GGWKmTqPPislAXy93xAJXDsC6sH3Ji4F+PlpJiKHox6lxhMZRJ2dFG5mzZc8JZTNCVcQEFBgL+orY8g/v372zdM7U8eo+XoQnHvU8fxYhIL76IPcETtIjLvqtG9euyof5ClnZIlQS8nEoK+QSeS7wPTjAx6tNlz5/iRA42Tr9UauCzEmRTYSUwnOMd+X8mZP379iCZJ9hn5x5P4dBuRl6NcQUHGQicY/zzhHGhfYRksbP0+2c8nQ1FKrdBgwfi9jwqxbMmqIlR2IR7wX3RdSrt+rnMCC0FcacI3t3bFXP9WvRKMqrE5JDCQnjyvYNq8JOQmOuHj96cH/2xJFhxq3IQoLBeACDwfTRg/ogD4RSnsjmNTp8YVj6nzi9bVHQ2rZxpWKFEMpM8nz16sULQxPZjpgyd0lO0VbnZnUqKd+na1cuheVryZE7j4Vazko16zWS93SFyMJ8Ikl6TCYEHztz0SoYVsYN6tVp37ZNayETvEVkWJqzjke/yjeC/QHzIyIeRXjH8S506jN4JNqQa0A97myibdezp09EZ94iqwtDKuSfOW5of3WOFYTwQl3se8ipo2wHa7l9D2GsPXn04NF9Ox3ks3zhnhaXgr7OiZNVuDXB2yc4wNcL4Y9g5EA+AT8v9zDlP4xMWXPkzI1/496k4f27y9BR8B6A18zN0Csm2R/g3QGPBtezp05gb9bigzw38BKBpxX2T5RBvgi8c/OnjUOCYs0P9oj3795G2B9kYXhAzV6xeTd8WLq2qFflQoCvN57VFKHOsB6QE0PkdDmubhzMYMBB+wij1rNNo5oIo6UlxLMnTxDWJ8wAGlPrBu1GZSzReR+eP33yOH0kodW0xop9GQacBdPHxbjxJiZZq9sONyogvBfCRiIMo/wNQFLsf0UIJ01xxH3kbLos6sNInklcCN32r7jw3zVXxfMIa1eURT8IeflS6/m3HDf7IgESIAESIAESIIGYIkCDRUyRZbskQAIkQALRIgDlPk5hvn///l3vtk1qS2MFFFs4eY/GXTUUScjbcHT/fwo7pRCd+w0ZBaUzlHqPHz64rxZQxurXpXiK1oBE5aZtu/SEsm/CkD5d1ApHtC10cZmgIPN2PxfhJH6brn3+gjJ5k4iBLuXAadrKNeo1WjF/BmJhf/XJlc8iLJkn4t9PWbBqE5S5yE0hCyEPCP4N48yCGRPClLTyU7RkmQr4t4+wMER3zKgvE4l7uTpra21EGSgkEe4LfJ49efyoccv2XaC4hRL1mVCMacmBU9C4L+wVEZQ6UPwitvzsSZ+NDcqPDGujroecECjn5nzmJBKbV6nd8I8BnVo2fCcmC/dl3gPIp2wP3ixIXIsY+lpJiJFXAOXdFfxNwVXYnPJDYQtNuD26AAAgAElEQVRG6vweyOGii5uyb4QDg3fNwukTRirXB8ogl8qjB/fuZs2R56scFugTymORByUks9Dgayli4amBkFtbVi+db4qxarWBEGYIV7V+2YK/keNEloGnARTueJfUY0KOmGtXLl/UUmKDA8KTwdCjlQwZXklQrsfU/oD2W3fu2R9zuWX1sgg5eiJbR43EPKL+whkTvnj/IOwbEobDAKpeH8i5AV7B/j5e8ERCgnmlYVB4Gtgi9wj2qRF9OrVWJrPGWkdd72+8P6BPzN/xg3t2wLuqtjBcuzmfPnn+zEmdp/yRNP2dhkFTrhWEFcS+369D8/rSWAFDBdYQysA4pGX4gycKDF/w6sHeit8UXesc7PGulKpQpQaMHOqk4qZ6P6Iylui8D+edTh6DxyD2aawfQ8aBPR77qavTqQhGIEPqx+Ey8IJIJq5c4kocfiGcG0KouQkjA5Jlw8gIA8aXj8KQASMF8lmgzO/iuiGuMAM0PqL+j+FtYi/GgQL0dV/cPyLaCMtTFW40wf+3h9EERg0YTZAr45Mug4lSFv6bBEiABEiABEiABOISAbqYxqXZoCwkQAIkQAJfCPQcPGoiTruPH9y7852bN76EAunUd/BImR/AV5zKVyJD7GwoSi8FBUYI2QJFZO2GzVqjvJYyEvdx6hh/Qy9rJ7yOzvRAZsRGh8fAvu2b16nbgtwYb5C/j+drkWBX+RyKSiQGh1JWKs/hLYKY9teuXr64WiNxKRTu4IaT8KLrhOpTyOWr1qyLPqaPGdJX7RFQslzlalCy3b19E0qTaH9sitiXwul/eXpbq0FpHIECTehJUyBnBAwDG5bP/1uXAP95WHxtsACvGg2atDi8Z8cW5dqR7UjFr9rwkK+ApQ3K+Hqed+nY+6/hMLA4HtkvTl9//kivlBuhIVA+ffm0EImp8WXz6iWaynkL4QUDha+PhiEqqnDBCKfNYZTYvGrxVyHMEC4Iyupb169eiax9nHQeKJKuu5w+cUTL6IW6N4SXjTxpL9uC0hGnuRdMHx9m6MqQOWuEhM5VajVoAqOB04nDmqGVojpuWQ/veneRTBoK97mTRw+R92FAke85PLNgdFH2VUAkSr4U/LW3AZ7DkIkT+/j3udMnjmqd9IdiFs9jYn9Au3VErgjM646Nq5dJbxml7FhH+K42wuAe8kzASwkKdnzHGpixZN02GFimjPirp5q3cKgJ88AStqdEMCjCc0vZp9wf1i6ZM0P9DpUsV6ka6nqd122ANGZ+bYoUL4Xynjo8sPBMOIK4Y06Qowjf+4+cOAPrS6xBnSf1YVhDGV0eFjB2IbTZ1rXLFirfcxiukEQb/ah/Y+S4YNyEYQOeLZF5eMjyOzevXYH9Hf0Zw8bQslEdS3TeB4wJ8sHoaaicWGtgqrW+DW0jLpYL95TA7zaM6zAYwAuotLiaigvGR+Qrwe9EWXEVFRfy4ySHkSHcGIEcFdhf8P/NYYCHNxWMFDBEwPiQX1z475de4e3CQ7K8uIqL578hdJT4N4wZOcPbxt/fxMXDiXFxwVAmEiABEiABEiABvQRosNCLiAVIgARIgAS+NQGEgmokTtjj5KoyvAmU8FBGSu8Eoaz0VMomTw2HCEWlWmbEGpe5BXR5DmQVJ23heWHIyXRjmSD0BsKoHN2/a5s0OijbsC1aAsoNTWWkfZnylaF4Q9gmGD6Q3HnLEeew0CXdWzaoplbK4hRvbpE4N9DX0x1Gkq1rly+8f/f2LdkfFGcI0+Tv7eGKE8pKOXByGcq600cPRhr33dDxIwl0XtFmoI+Xu9a4ZTv+3u6uCB0EuZBEGwacVQv/nqoOdaXs9z8Pi69DQlWr26gZFNAO65Yv0pITbHD/yqXgQOVzxK9/8ughTrn+ULlm/cZzp4wJO2UtP9Jr5crlC0HyHmQoVb5KdZyg9nGP6JEChSbCoCD0TmRjMZSnLAcDHP59ZO/2Ler5F4aVMI8IrbBHsj4U49MWr3OA187w3h1b6QrbhPBjOGkvkz+jPhS6WDtQ8uK0eEZhPVPLj8Tkjx7ev3fOydHoGPeGsBg0btocvM9De3VooVR+wlsA9XEPxj9lW/CsgTeImL4I+0O9pq3ayWTBOveHcE+TK5f+m39DZDW0DLxWwHP/js1fwrMp62KPgHHR283FSXkfuRzgJSDDuiHp8pbDzt7wlBrQqUVDLQMNFO737ty6CcMSjBwnDu3dqWwTycqxz25cuXiu8j6Yl69aqx7aVHttGDpOdTkYKWGM8PV0/coArSwHo8OFAD9v7A/wVECIPKcTRw5ovXP/vZufQ8ZpeVhgLQwYNWkWQpbNHDf8Sw4cvM/d+g8fK39jgvy9v1pDsm3xSoftIXvFbxQ46hv7tnUrFsNY3a57/y/GNX11DH0e1bFE932AV5ynMOo2bNGus8yNpE/mgtZ2RaVRTV9Zc3sOTwdxwZgNz8Tb4oIBA8aLzOKCkQK/J8hdhXCQ8IRqKy4YIgqHP0fCeRguEB4KoaKSCUMEjOgdxQUjoZ24UogLHhjpxIUQY/A2xVrEHoznaA+eHfjAW+Or8ITh9/mHBEiABEiABEiABOI8ARos4vwUUUASIAES+L4IQNk+bNLfC5GXYI7i5DQoDBg9eRYUkefOnDiKMB1qDwCZ9DRUaBSV1BA6SZxAbQqlMhRRF3XkqIDST13XVPTlqeSjIqeCVpvFy1aogvterl8rI3EP8dKh/MUJayTkHTFlzhJnx2OHm1cvbfd/9u4EXre5+h/4uffiKlPJVFInQ+Yx0YAokqgoCoWkImme+5eGnzShQZMiNJJIiCShDJmVTBm6hmSeMrvDf72PZ932fTxnuGe495x71n691ms/z97f/R0+e5/vfs7n811rdSLLjANRbuX7gqEYIP6bbW79ph13IYA0w+jk+S222bYnYe8ZDc+CoWCwxjrrb4Dk7JSXo1kvrxKhdiS43XmP93xAnPqj+gknFNxiDyH5RDwszbp4AIj/j1DriHWQnQjQ666elbheadXV17rmyssv22n3vd7317+ccVr79YQHocmE2cp619vgpRtbzd4U1pptbrDRpq/yTHe6r0PB1TPt+vM7hFYh+Dknl0tvbXzhoO8f/uxg6D+59+47pkjTqewtNz6ZpyBXnCMmN978Ndv89lc/O9zf0u23/vvmZSNMW/Naq6h5b/zqyEO/1+69M5Qx57Xu7yu2eO3rhU1qejto10rzP558/K+trr+uzZPC/XMvIjfHLPMDcUsIIPODNnpbVe/vyniy3HCMJevwDK27QYiIkS+i+Xzl+WctsdTSxERzV7vwZX5Q7pH4I5IU/JCjTjydOPjWrTd9see4Uz+FzrvnrrvugOX3D/zSLEnV5f8w1jNOPen4di+k9V+68abEq6ZHwlBwkEdjlXhWrvr7ZRd3CpPXrJsHiefqo/t++SDCTl/eFa7rbX5w7t0f/OS+PK3kp2l6YAjJRQA667TfnaDcdVc/1VvP3Mq7yfmBhjyTO+jnh373m57RFKeHglvz2sGOZah/D/rwgwhHJxTZW3Z793v7G49nGOYZequ/8mP1vLwSYfdG/78edniYcGG8FeVn4TnB+0JYtbeH/SiMePGeMF49BAtChLBP7wh7fxghgvcFYWKJMF5jt4UJa8n7QnioF4QJK3V7mPBcl0cf7uL5UeGgAo3aCoFCoBAoBAqBQmDMIVCCxZi7ZdXhQqAQKATmbQSEzFhjnRdt8LMIBZTJVY14sy232daq2p/+6DsHIYv+1WGVszBJVrG256fY60Of/JxVnQQOXge9kahIupsivv1IIGxFs3Y7rd4mHmQS407nhUxB9uz3rR/9lEDxzh1eu+nH37PbmzOBdnt/1woW3bFVIg79MT877AfthPQb3vy23YUoEgu+/dpXR94GJGWnsDODwSUTaV/cIZF4e30EAmF3kJiHHXzA/n15ZLg2ivUIFrE4e2aiXlgSSS467+wzO8WK5y0grIwwSM2V+QjuF4QIEGT0DeKyH/LNr3yxvX8EsXYRIPNe9Da+LbZ+UgDqlJdkMHjmNRmeqNPfgRwDkfrlMSvSO7Xxtne990NW8x/81S98+tK21frt5SMyWE9YqRQsXvOGHXryx5z6218fZc9LZbnuFXrC5+S2xz4f/TQB6uheQmQNZdyu3fujn/kiwfLQg7/+payLKPbxL3ztWz35J2LlvePt2Cy7XDdSr6s93v62O+7yjmcECy9Bt2fi6stn9czINswPvApGIpwN8phw0ttzZH4gtlx20flPyW+TIZWIUAjhz334PbvvuNXG6/WWa4MniVBR4bC29tX/+PulPBWa92Tbt+yCKA3vnaeKq6/eZrs3O3f6yScIcTPkjVjhb28g80PMjefBiFj3p5i7hAPrqwOd5gflCS48zzz7Z512co8wYVvmOc9dTuJyx2Oavcn8wQOjvY300Lrq8ssu7uS90luffnHY97/FG+ptIYoMGbhWBUMZy1D/HnSBhx4h6S27v3sf96avca3cCmk25frhD7k4XHgOZz0Eg6iPt9RBYceECVX5QBjRgReEeZOnnHxS64cRwRZv2VaxXytM/qRJYQQMuTEIEjys1EX84MkhZKa/BV5SvJSIGY+Hd8ZwDqfqKgQKgUKgECgECoFCYI4iUILFHIW7GisECoFCoBDoD4FdIkmslbY/+cG3D8iywgP9v6988wfI0yO//62vC8chVE17XUsGWfeff988c/W781Ylv/p1b3rL9yMZrZA/va2etsJ5yaWf/ZxOBFV/fR7IeWR4RKr6W6ewQFaLEySQoUL0tNcnhNMVf7vkwl1et9mGe7zpNZv0JyakSDAtFJKfHnLwgc36rO5FdqvjKTkcAp+eldXhXdFMsjuQ8fVWxkpu4Yb6Ct2S11pd7jNh6bhfHGnlaZ8bYUOB0F5mChZLhduAUCe9kZmRqHcXBKnQXM3KkaAIN+Fpgoi8BAnXPO8ZFNKrPam2+4rY7DQ+9/QVrVwhhLL+xjM755/z3Od3K98U9XxH3PPm0Z9Ogo/V8x/49Be/+uc//v6knxzyv7+x3tpOb4LQAiWTjTwLO+925qm/+y1PE9+vD8Eik1H7Tmy0av/Yn//4kJEIrSZZPA+SXx35o+81n989gmh2/Ntf/vynEM/60j5HSGrveHOOEALoXR/4+GflAXEdkYfY0wkPfzcjOT9osz3cU/bjjTvv9i6fOz1H5gfzxkff/bY3vWHjdVY64ZifH9GXZ8ua620g9EzPs/Lj7x4oRM3MzTzIS4XgdO5Zp5/aPCccHQ8o8/BwrZI3P2hDvpj+nv+cH8wnEs33V/5/88P/BE3XvHnXd+0tx8uPvvlVoXl6NmLQ5w/47o/nX2D+Bb762Y+9b5U11l5XwvlOf0Mrr/5krptTTzj26P760Dzv7+HEX//8yE3CQ6kZYm126mgvO5SxDPXvIftiEYG5rr/8HJEjaG3XSHo/lDGPpWtbHg7G6+9s+7C9wzx3QuVdGHZ8GI8LmzwUvCWEffJZnhlCxbPCzgz7ZRjBkjghlKPcGLwnr4l2bm55dkznUZE2lrCqvhYChUAhUAgUAoVAIdBEoASLeh4KgUKgECgERg0CQnEgJP9w0nG/SkJU54RAEobjU+/dfafgRZZBNt16841T2jv+rCWXWvruO263unDm9qHP7Pd15K1V1RIF3zzlhlkSJmfB571gxZWQVu15DYYLHIR3b0mQd93z/R/VTqcQPkg3eSCsZJU3YCD9Qbord+pvjz1KaKTmNcJB+f6Hk37zlNBUm2/9BoRKl9XLA2lnIGUQ2MZl5Xt/5XO1//cP+NK+vZHGzToID76HYCHed8+2ZCtUSzuRn+ff9Na3vxvRfdpJx1vxOnPLmPQEriPaQmgplOHGrm6Lae++qq/T+HZ8x57vc/+c65T8uz88+jr/zGgXKd3uZbPxK7fcWp863cPF4qKvfu+Io++6/fb/7PuhPXdreqAYt3A/7W2mN4K/D6KO+4kQz3I3XHPVFT5nTo0P/r//+xovJ8LiUMbX27UEE+eO/fnhP8wyhIp3f+gT+wpTJG+Je2ls7ZgvHvMDIa4pdPA2Ca+bRX7yw4MPXHm1tdbpbX7QFjFvJOcHbdxy45MeLc1tw40325zY6tg/Q/RsPx9T47OICDymestF0rwm5weCTvtzIj8FL6Q///GUE9uTVXs+enu2BnuvPU/6PJCQacZoPvvdsUf9tDfvkWY//jc/TJs5Pzi/zfY77WrszXBZO+6+5/vgLPk4McYzdOvNN03pNK5VVl+7J/l5e96PgWAgLxNhNEMEDuSavsoMZSxD/XvIfhEwzXGEmL76GusQHpZnhRg21HGPwevlkvhvmKTchIqdw3gy/TiMZ4SQUYRSz6rQTjwtlgmTgPvMMPPdD1r7f4Qg8e+W/Tf208cgHtXlQqAQKAQKgUKgECgE+kRgvsKnECgECoFCoBAYLQhstNmWryUanPH7k6w67Nne9YFPfNaqXrHGEfZJikQOaf/gz7JZWd8k6K34FEZqt203f9kLVlpZMsqu3hKkvmDFJ893CrEzHPiE5rBw5POeRUxR7xbbbLeDuOY+S0zd3taiwUY61p6nobc+wWCFiPXi/LG/+B+p6ztsN91y6zcgujuRbTw9rCjulBdhMBhY+S30zKknHDeglchW3m636YtWGegq9knzTer5HTMtWOjsHzHL5/ZE1I4Jq4OYF26qnYzNMC/XhRuMcFHt403Boj1hc9zWRe6Kldjt5Ylvb3vnPh968r4Or3eFOsMx4GmPBAPY3u5OQbwSe049cVbM3fsvRUgxgs47tn/NJu3eD4Q9+Thes+Fqz2t6+QivRhQhSLx++5138/fVxCdD4qwYzxxRkeD49c9/4oNyrgzmmenvGt4bCOVM+Oz5+sZhvzw+mrvt8x/ZuyeUEXFFGLR20cvfRkTkmUmWCi0nBNCh3/7afp4HCblvP6FzAmXtEDxHbH5YaJFF9L39WeLV8JHPfqnHS0ofr28JRE2czBGzg3d6YB3/y58c1i5wCBWm7j+2eSA5tmnMD/ZnnXbKif3dp4GeX33tF71YrpGmQN3XtW/fdouXx73OFel9NgM7BZrzg3k+ImIt//NDv/fNFOyEUPvIZ/c/8C+nn/o7xz0n7vfFfz3nz50akEuIsNWXuNVbx3jKCSmW881AcepUbqhjGcrfQ7M/xmOO629MRx1+yMFdXYcMZchj9tq2PBIECeKE3zA3R+gm4Z2EfZK7wmJCZj4g8nu3med5Xtwd9Tw+ZkGojhcChUAhUAgUAoVAITAbCJSHxWyAVUULgUKgECgERhaB1dZeVxznrstboYG22naHnd/zkU9/wcrhDF+zdDDByjz43/ufsmJfeJfg9MR87hKm5pP7Hfidk2NFp/A+8ls4fsd/br2l0yiWX+mFqyJekggd7pE+HuypcCvNemMh82If+/xXvpnJZm8INry93Ycf+q9VmUFQP0nE97eJZy+Pg8S97WGKrGYWukO8+Pa8FsLhrLTK6mvK/dBO5vfXZm/nV197vRc7d8kAwr1kHQMVK5SfFIykfTOHxd13PkmUC9/U7Bf8kJKI+iN/8NTV/wh35Y/5yWHf7zSeFVZeZXXk7r+umzX+uuTwEpu3X/Op/Q4SrqNnCx3mKfd1sJjmdVY0R87xWZ4JxKtV4ice84sj2+/vO9//8c+8fLMttvrO1774/zolI/9DhLeBUaeEwDf88+orl19p5dV45xx/9E9/3Aw3ZKU7XNzrj37uK98gYBx95I9mjn2o42xe7xn1/Ob8wBPgW4cffQJvk4/vtesOKcKEULZcJ4+XJ+eHR3rmB9sn9zvgO/cE+42kznj+vQmaMf4eQXOkwtnk31xMEbM8S2/dY+8PIoL1OxwMrovoZzPDn+U4QoP5bzwKA5ofeGutusbakvh2/f6EJ/OQ5Naz8n/Tzbc0H519xmkSBc+ybRQCMO+ZTnl2BnOfJXB/boQau+SC8/oNB5X1m58H4n2lfES8esr80P6OIUR+/ZCf/jrChN342Q++e1fX/e8d81SvsJ5cN/Es8HgbyJiFYBN6K8tOjC8+d7qPA6mvWWaoYxns3wPMiJPNvkyId05zHp7dsYzX8iFW+Lv1ntwkTE4mXoP+P+eJwfPC4g2/AZYOe0aUr8WG4/VhqXEXAoVAIVAIFALjDIESLMbZDa/hFgKFQCEwmhFAPOrffcG2CnWx3zd/+JPIRXDJZz7wrl1yNewCkxfoyVuApGsfyyMRa8IxhP3nvv7dw54ZrPW3vvy5Tzq2yKLPeIZ9b4Rk9wovXEUImYGEVBkMhohd3h4ZV93q3/2+9cOfyJtxwTln/Umdt7Xl33hynA89KLxR++pVgszu7/3wJ9/+ng9+vNmfDOuDjGxPOr3uBi/rycJ5xqn/82DJa9d+0YYv8znJ4MGMsf2aVdda50WODSQ+/WDa4zXgunAYmelh8e9gdZHVvEWadf6//b/xfV4PX/nMR/bptJp7hZVXXR0pfPJvjv55p74g6R4IsaNdzHFfrdhODwzX7rbXBz7Gu+f8s888vbf7OpjxNq9BnHuGhGlyXKiefb/+nUPlSDnkG1/5QrPsBhtt+qq9Pvypz/OM6CTWKJuYPBquKe19swKemLFErDo/7hdHzJJbBLkNc3+v8BX/v5n/xN8ibDI8z1DGbYyuNz8guw856sQ/rrbWuuvv++G9d28+txGFa3KnXDGPhntFti/pMs+tA7/46Y8QKnlPONeboGl+cD6TkA9lHJ2uzRBHm2y+1evyPPFon0/s+6XzIpcEMYEI2elaz0Imq8/zcN/6jW952+cO+O5hzWvU6bnhrZb5SfL8CyMJNxHo3LP+eGp77gYeB55z+V2GK7/Nqmut2zM/XBIC6nDjqb7/zQ//88BqvmOE2Tr0mJPPVO59b99hmxS8PD+uj6n3Ke8YYoV7IeF2f33mzXXk8X88d88PfmLfLGvO9rdw4bl/GZDg0VcbQx3LYP8eDjv2938+8Ec/Py7xJZS+aMOXb3Lheb2LOP52JYU/+Mhf/y7/1vrDb14/3xIrnhnj5NVkbhPaybuMqPqLsG+E/STst2HyVtwlJ8a8jkuNrxAoBAqBQqAQKAQKAQjUKo16DgqBQqAQKARGDQJ33vZkvoVjT7/gCgSckBvv23X7rdMDwblMmv2hz3zpgOtj5XeTdFOeKBBE5umI+899+D27Z4goK0AR+J1IKPUKeTNSZKT6T/r1L37yif874OBvH/GrkyLh8zG8R4TPOeX4Y35x1d8vvVioq+DB5u90M0757a9/aaU1sks4nHU3eOlG27/1HXsibb/wsX3e2bxm7fWfFB7EeW+vSyJZx4Q+aT+XCVintHkQDOXhkBOAx4SwQkOpp79rQ7AQH7xns/r6d8cd9bO37Pbu93543/0PPP8vZ/xx27fs8o7Nt952e2T97wPL9vp4vsSi/Of/NrwHesu1gXTvlBAdzgSKb/74qN/+JBKcW/WsPc/ikd//5tdescVWr+vtvvY3rr7Oe27kPtn3awf/6A8nHvernXbf630I5c9GbopmWDSC2JcPPuwXCOwNXrbJK3920pkXnPmHk0+48Nyz/uTvbaFFFl10zXXX35An0x0RZ63TavcrW+TsmaedfEIn0lwYo+W6l1/x9JN/e2x7QviDDv3l8TCQx2TnrV+x/lDIbmGf/A1LNPzGnd7+Ll40B4XgcGqbp4A5wjyw54c+9blDvvHlmeLNTVOuv04YqAN++LNjhT7iiXJWjAnO5gf70Hse6IS7+YFY1VtulKHcS9f+9c9nnCbJs9BcER1q0eDMF9x1zw981HiFwzv8N6ed09tz9PvfHvPL17xh+508CwS350dfd3jbHnsh13nEdJ4ffjmb88Myz1HP8M4PTyavvuT8/hNuDwXf5vxw52239bxjPve17xy6+BJLLDVjRteMvd+67ZbNcd14w7X/FAZtux133eOi8KSQoD7bJ+r43O691ql/RCjzwB77fPTTwvTFHPM8AptwfBe0xMyhjGuoYxns34O/mdfv8Na3e89GSpgnNnz5K17F8+VnP/zOQb2N5zNf/uYPhORzfpnAYaAhwIaCz2i9NoQKQjvPCp5O6V2R7/774hgvwavDJNImUDzFq2q0jq36VQgUAoVAIVAIFAKFQCFQCBQChUAhUAjMcwhIanvsny644uyrbn3g6z/4yTFW9XYa5D4f3/dLF/7r7sfbV9ELeXPJTfdPv/jG+6a9Y5+PfKp57XY77fbOS29+YIaV1e11Wil63j9vf0iImJEClWfFj4879S/6wPTz8wd+78dWriOxHEMCdWofMXvi2X+7Lq+9eMq9U8XtX3XNJ0O75KaNc6+57cGDDv2FUBJP2Q779Sln/eoP5z4laa+CVsjrUyZPHg4cTjzn79cTaYajrk517LDLO9/jXmf+kSwjubRxJl6ep53esdf7e+uHMEOnnH/lTc8Jxr9TGSuitbP/wYd19L5AMmdb9u6zUDdWYv/5ipvv/eJBPzhiJDD49P4HfS/b9fxuv8see7W38/5PfeErZ1/17/v3/thn/k++lA9/9ksH/PGSa//T7K/Pvznz4qszsXN7HXIeXPSve54gbHQax7ePOOakP112wx1yQDTP+7s6//o7H1U//NrDdA0Gk/d94nP7u58n/OWyaz2zneogdjr/y1P+cknzPPHmzMtvvFt/rBBvhlkjuDh+QIQH6lTnd3963Cm/Pv38fwymzwO9hohywQ13PZb35uTzrpjy0k1e+WrXw9j3TnXBmWDWvKeEqSSIm9cc8ssT/njqhVff0h6eThmilXm1033iPaP+N+789ncNdDz9leP9ccwf/yp+/4hs5gV93v5t79gzGxAGyb3098L7obdnWvJxfzcf2ffLs5Dw/tb9raR3QX8dJxK7b/phjnn3Bz+5bzNEVH/X93V+qGMZ7N8DDwnvEmP6y5W33Pd/3zjkyPYQUe39Pvy4P5ytvL/L4TJ8EUYAACAASURBVBr/ULCbm9eGYDE57FU/3n3jA2J/StilYX8P+03YEWFHh50Q1j03+1ltFwKFQCFQCBQChUAhUAgUAoVAIVAIFAKFwGwikAlV2y9DPEr23H5cSIpvHf6rEzPBdfM8kr5HzIiExbPZjdkqbpW79q3+XmqZ5yzbvPit79z7g8981hJL9lYh0pzXCAKzN+JX/a/bYefdegu5IY8HIr1TG+rPZLyzNag+Cq8XYUKEmBmu+trrkQMkQ2C1n0OKCX8Dr+EIQYKM59HS21h4YAgDlSGashzSeNU1nwyNNRIbQjTyDrwmwyW1tyF0GJyax2HjXr92uze/laeP/BP9EbB93UfEZ2/P5HoRhownCA+ikRh/X3V2miPg1Azf1byeh0KT3G6eI/LwzBjpMfAA8Rx5ZjJ8nDZfuNqaa7/6dW98c1/tu8a15sDeykla3pso6TnJvDOdrjd3DSfZnEmjRxJTeAy2z65r/7sw32S+m4H2Wx1E0YGWH4lyncaincH+PbjW+6q393D7GIiIBLHe3j8jMea5Wedj7+ya0LCJrc8Tf7b7Sxf98e4bvSvs54fvvtH3D9/95X89YveXXxT2tTi3WhzfJ4SKv8b+/LC9TnrHWgs265qbY6q2C4FCoBAoBAqBQqAQmJMI9MR+rq0QKAQKgUKgEBjPCGz5+u13/Mp3f/xLoUHE+R/PWNTYC4FCYFYEeHoRLH78nQO/fPBXv/DpwqcQKATGFwJEgxjxjNaom58d8r3n2ORDu2ZEWYnVmdDLQs0J6TTjounLL3b9jGV2i8+bT+ia8bQZXROuCZsWn29aYsIDR2048bp7/jb9+YvcPONZH4vKnju9a8Kz5+uadshrJl32m0W6HhUaik2LNqa1+jOzTZ2IY9mXWfoZ5WsrBAqBQqAQKAQKgUJgzCFQOSzG3C2rDhcChUAhUAgMNwIZWunaq68csfAkw93nqq8QKATmDAL/mx+uqPlhzkBerRQCcwWBlhDQbJsI0UWIaIkCRAIiRIoWhAn5JxybHtdLnO3/a8cWdPyeGQv/N0SIJW7vWuy9k7qmvzrsaRO7pj86vWvifYtOeHj/F0y486bnTbhrWogTz3jJxGunzjd9+qG3z1jsy491zbdICBrbXzN92RvXn3j9P6OuR8OeiDYIF9rLNgki8jhln6a3+pt91vVZFinmeOYKyNVoIVAIFAKFQCFQCBQCA0CgBIsBgFRFCoFCoBAoBOZtBDZ4+aavuvfuu+4cqYS68zZ6NbpCYN5GYIONNn2VEf7zyn90zP8yb4++RlcIzHsIpDDRJkSkGEF0SIKfx0QKFHmMSNEjRrSQeUbsJ4cREmzEikda35d4vGu+JR/sWvA94SXxhskTpirzwMJdj96++IQHL15hwu0LhYDxwji2kAvj830bTLxu4lUzlr361hnPfP5jXfM/679dC773nzOe/ZUXTvjPvVFEsu5Mwu3/+MfCJOq26TdRgweGjWDBZhmPfreElR6PEAUbQk16Z7Sq7BFraisECoFCoBAoBAqBQmCOI1CCxRyHvBosBAqBQqAQGE0IiMO9yhprrXvGqScdP5r6VX0pBAqB0YHAy17xqi3vv/eeu/913TVXjY4eVS8KgUJgdhFo857oERviGILeZyKEPbHh8TDH03NCUecWaZ0jGDw7jIBxT5g8Tc8KuztsmTDiw3WtY8+L/VqLTXh4i8dmzD95oa7H7glR4m/PmXDPP5eY8N8rJnbNyLaeHuUIHwtGiKjFVplw643zd027+8EZk5cPT4zF752x0EemTph0QHhhLB9lHgq7rdEmcWTxVp//0+r3ArH/bxixwmav3/rsnM88QnhmNAWNLO+ap4gXrbpqVwgUAoVAIVAIFAKFwIgjUILFiENcDRQChUAhUAiMZgQ2fuWWW0uKesHZZ50+mvtZfSsECoE5j4BE9ZJ0//F3x/96RmxzvgfVYiFQCMwuAm3iRHpGpEeEv2MeEbwkEPf+H2bKEQ14LPBkQN4/GIbUXzKMGGFzbIkwwgGBQD2ECQLHM8N4URAtXjqta+K08LB4elR8fwgR8y884dGJy0y4b8qiXY/whOBZsWqrXW3ol/YXiZBRty074e7Tbut6xuohWMhnscaUGUuuvcKE2x6OurRhI5roAy8Look2iRELt84TNW4PI8YsFmb8xI0co/YyN4a+65O6Eq8e8aIl6vRU2R5KiidHeWC00K5dIVAIFAKFQCFQCAwrAiVYDCucVVkhUAgUAoXAWENgx933et/02MrDYqzduepvITDyCLxl9z330crpp5xw3Mi3Vi0UAoXAUBBoJKNu5pjIz8h8QoXvCHqf7ZH2PB0Q9rwoEPlECN4TCH4CAQ8I/zc/t3VeGdcg+FcLWzOMl4ONULAim9o18ZHwqHjGol0PPzh9wsSpS0544Oandz1G7NAuEYQ4oj8EhztbbfUIKk/venzGcyfcc+19M56++NSuScs92jX/hjO6Jv51Qtd01z+n1RfX6seyYca3dKu+W1p9JmJkKCmihXaN8a4wY3TeuAg36XmhfeNSb2LXkyOjJV7MDCUVx2orBAqBQqAQKAQKgUJgRBAowWJEYK1KC4FCoBAoBMYCAutt+PJNJNQ954zTTrnjtlv/PRb6XH0sBAqBOYPAQgsvvMgbd9rtnfffd+89f/r9Sb+ZM61WK4VAITC7CLR5VPj/lleBjaeE7wh35DzhgUAhXBKBojuMJ8HDYUQD3xH1/2od93mlMGS/MsouF+b3gjZco27CBiFAe0QD7Sy+QKSTCIHimeFlcf8iEx695Gldj+kLYYCpi4BAIFBH9pUHhz5OXqBr6uKLTXhkvodmTI4Lpq4Sxx6Lwo+HiqAv2nSdPmRIK8LFzWGEBv107srW3vjXarWtrzDQJs+Lq8NsxBl9VD/vDfXqi7Zs2pP4e2aOj9bx2hUChUAhUAgUAoVAITCsCJRgMaxwVmWFQCFQCBQCYwWBibG9/5Of/7L+HvH9b35trPS7+lkIFAJzBoE99vnopxdaeJFFD/nGl7/w+GOPIjdrKwQKgVGEQIs4z1BPmTQbCU9gIDb4TBTgZaAccQCRj7BXnreCTRil9K74R3zm/SB0kk1dxIIsl3kqeDG47v4wAsRSYT3CSDQyMUI5PRE5Kh5dcMITD0fuikciJ8W0aFA/eEcQEvQrPSLuaPSJ14U2iQeTJnc9cV/09MYQPeZ/omviC+OiO8LLgtihXcLCCsqF8f7QB54TwkXZUqxIDwwixRphvvtMHLEZK2wcuzUMVszx9L4wRm3atJ8Ju6e3h4pqlaldIVAIFAKFQCFQCBQCg0agBItBQ1cXFgKFQCFQCIxlBPb80Cc/t/b6G77srNNOPuGi8/5y5lgeS/W9ECgEhheBl2y82Ra77vn+j97+n3/f8tMfHnzg8NZetRUChcBgEeiQn8L/s8h1AgSBAnmPtPedgCD0E+JdmdXDeBn4TiS4IgzxTkggIqwXRqyQk+KCMKGTXPdAq05tnRMmZJIwUClYEAi0JaxTiCATJkfeiYcib8VCC3Y9sVjskf42AgWxQD95MBAA9JcYQKRQv/4oT3wgotxPtAjBY/FQCRaKung86KtzxuIzoeFvYUSQlcMyH4WyNl4im4QRWYznklb7mcMDLtrTH/UQbdQLwx5vj5apVx95XOhnTzJvuSwa2yy5firHxSzY1JdCoBAoBAqBQqAQGCAC6S47wOJVrBAoBAqBQqAQGJ0IvGKL177+64f85JggGG++8Ybr/tlbLyXYfvcHP7nvXh/+1OfvvP0/t35g9x1f//BDD+Yqw9E5uOpVIVAIDAkBybMP+/UpZy286GLP+PslF5zXVwLtTTZ/zTZf+8FPj5kvto/uucubplx/7TVDarwuLgQKgWFBoCVW+P8VMZ/kvvBL6ZGAZCdW2IgOPCjsEe7Eh7XDiAuIe9c7psyLw14ahth3PSNAZKgo4ZR4WWiHeMGrwTXNXBjIf8IH4v9poQpMDHEB45/eGsoydamfSIHc50lBfED+66djRA2eHMbq2OJR14zw2CBy3Bl1piBj7Pq/fBhhQZ+7wwgpEoIrr951w54VBh9l1a+M3z5ECPk3JOjWd9/9hlIPrw39TVGE0KKv2jUWdWvXWJJXmEWw2I80UlshUAgUAoVAIVAIFAKziUAJFrMJWBUvBAqBQqAQGJ0ITIptp0igvV3EnF9x5VXXsDL67jvvuF1CbT0Wj56o8cWDfnDEa7d781vvuevOO/Z+23Zb3nLjDdePzhFVrwqBQmC4EHjiiccf32b7nXfd5k077brJq7ba5q47br/trjv+c2scFjama1KIE+tt8LKNP/DpL3z1vR/bd79JEydO2vfDe739zD+cfMJw9aHqKQQKgcEj0Aj/hMBH2CPNvd95ARAFkOY2IZdsjr8gjEeBBNpI+Q3CkO+Iep95PDDHCBuumRLGg4JA8cKw9KRQl2Tazw/rbl2DwEfo89hwvqeOqOSJsMlh+qcM01991x9igbnHMddql/FccI5YQWAgQKjD2ISKWjAK8aAgOBAOjFvf1e8zMUIfbAQZokp3mHH4rUPAgAOxgVcGgcI1yshjQcxxjqCjXWX1hzdKJgpXR+bhIN4Yj75kaK6e31y5lWDRRKM+FwKFQCFQCBQChcBAEciEWQMtX+UKgUKgECgECoFRi8CSSz/7OR/41Be+stW2O+w8MQSMqVOfeOK/999/33zzzz//IrGyWsetrP7TKScc95XPfux9d91xmxWItRUChcA4QGCByQsuuPveH/rELu9+30cImMTMB//7wP3Tpk6dutgzF3+WvDZguOryv12y/6c/+J5/XHaxkDC1FQKFwFxEoBECKnNUINAZgp5Hg5wL8lIQEhD3mYeBqLF+mHBHPvv75s2gHoIF4h+5LsG26wgOziHnHXMtMYBQcHerjsyH4fdE1umcjcjA24CngnoJJ+kJ4TwRhGBBSGA8MrSjTIaDsphQXwgCxAzX6Ku+S/StHIEkx5khn4RygsVtrbZ9J34QXYyJsDAlbNVWvfrz9zDjI2Yoc15Yhs5SV4aO5iPx1zBt8SwhpPDCuClMgm/jhKtwWPrKZua4qPwWoK6tECgECoFCoBAoBGYXgRIsZhexKl8IFAKFQCEw6hFY5jnPXW7TLbfedrU1133R4kssuVTwkVPvDZeKa/7xt0v/cvqpv4ugUUiC2gqBQmAcIiCR9iu22Op167z4JS9f+tnPXY5Q8cD99917w7VXX3nB2WeefvmlF50/DmGpIRcCcw2BthwIzX6k5wHCPol+QgXSPEn7G+MzIp1okYmnkfvIfl4FW4WtE0bYQLLzEECwEzK6wzI/BYEAge+8xQy8C3gOIPblupAvwjEkPcGEZ4Y+Ie95QhAbfBZCTv8IIvooRBIPDyKE7z5rhzhwcRgBQr3adVy/jVuoJ3Wm0EEY4ZXBC0K72W/CBIGAWJFiCcFBvzdq9cW1yhmDPhBlMmk4oUcIqLPChMjStsTc8nlcFMbLTBn4GJO64AMHv6Wc02/1O0e4IG6wHuGiRItAobZCoBAoBAqBQqAQmC0ESrCYLbiqcCFQCBQChUAhUAgUAoVAIVAIFAKFwHAh0EGwyP9R7Xk1INmR4kj/zEmBuEeSM+IB0YCw8cpWWcLAmWEbhiH+EfxCIKlPWdekyKAuhHwm8CZ48BRQnkhA6CAq+I7UV0eGRSIo6AOCPhN4Z74IZQgS2tYmoUR5RD5victb12lbHUQCHiLZVx4ZvCXUm94d+qpvxAFYqCs9MVxL6HA9AYPgor8EBm0TF+TlUJ5owctDHY7xKNNH7Rgzzwv7o8O2CZPfQ/2nhqWniD7oO9NGYmWvD8akjcxrMUt+izjeVUm5oVBbIVAIFAKFQCFQCLQjkK6ehUwhUAgUAoVAIVAIFAKFQCFQCBQChUAhMDcRIDow5La9kEkEAMQ/Apx4gTwX3giZz3hY8LzgpSCUE6EAue76K8N4WhA8UtgQxgiZj/gniiD1M2G3PbHj2jAChbLq5aHhHO8KYaL8H03w0E/ig2syibe+KofI1xf90E/kPWEDoZ85JzLHhnP6ok3eF8SD9LTQRgoi2vCZaOCaxIV3h/6oW/+Mj8iiXdcorz7X+i5nBVGCpwUBIz0+UpThQQF7ggbPDGKH9uCq78bLw4JAop2rwq5rtaEuwod2CCqZayQ/x6HaCoFCoBAoBAqBQqAQ6B2BEizq6SgECoFCoBAoBAqBQqAQKAQKgUKgEJjbCKRY0QwBhUBH/hMLkPE8A6z4l3MC6S5MESECcY9MR5SnsCFM1JQwHhKSS6vDngBBECAmpBcAgQIpn6S+cwQNxD+RxHHEPnIecZ/5JFJYSQFEQmzH0kuE94J+CdOE3NdPQoA6iAyEEP+TG6ONoKB/PBTUkfksMnG3PhmH65lxuJ4goQ+u1zfjghVPC/1RVl+IGsQGuPruM+8L174hbErrOqG2JBknABFtCB/qFS4KBvrH24Ow4V4QI85t1a8+7biPwlRliKj42LPNkpg7D9a+ECgECoFCoBAoBAqBRKAEi3oWCoFCoBAoBAqBQqAQKAQKgUKgECgE5hYCzVwVSG7f/Z+K4CcwIOWR9DwWeAUgypHmcizImfCSMIS7EEXIcAS5JNhEAN4YW7QGRixwHpGfIZqcSvFBDoz0IEC6K68uHgVEBm0wZH8mztZfZbJ/vAsyRBORwGd79REimO8Ifx4IPByMkReDttN7IvNdEFJ4kxAA9IcgYlNOn4gR+kLYUIYIASfniBuucRxOhB2iTOYBITYQFCTVVg6OvFm0R4Qw1tVadUq+7Zy+G6NrHYOlXBnafVmYfBjaJxzBCc7GmSG74mPPpt9PCRGVJ2tfCBQChUAhUAgUAuMbgRIsxvf9r9EXAoVAIVAIFAKFQCFQCBQChUAhMDcRSIEic0OkgEFI6A5DnCPZCRBW+iP5HROuSO4EJDkyXRmeBkQE5L9wUIh3xPmZYUh2dfIYQNS7XpvKEjsyxBPyXj3pCeGzLT0D/A/N24NlLguEPIHANekxkWGa1J9hnoRNQvpn/zORdXqHZD+6W/1Uf4oh+kDw0B8CAS8KYkCGn9IejwnHCTrGARNl9cvYbfCBAfFigzB5KQgq6pJ8m4CyWRiRg2CyShgxhxABN54UJ7fq5YGhTdjCmUCkPUIGPOzdM5gQKGCWobFKsAgwaisECoFCoBAoBAqBpyJQgkU9FYVAIVAIFAKFQCFQCBQChUAhUAgUAiOCQIek2tkOYSJJa8Q84h2RL5QTYpsI4JhyyHOeFUIVSVZNiNg27MIwJHp6ACDHeScg6lOA4JWwZhixAEnPg0AZxD8RgreDc8oj5Ykf+X+yvfYzxFF+j0M9gkAm0TYOwkLmllCeSOBapD2hAfHP84M4oTxCXzmiyTlhPBQIDcrqlz4SFrKfiH5jhQm8YKQ8ISJDYSnruL7Bz3iMX1+EpSImCEPlGmIJoQKO+vGXMCLO6q16CUMEIf0VVstx7cCf6MGzwrXCTp0Z5v4wuS2cz/BX8NZfooa6jJuHSFc8GxMi8XYJF8CorRAoBAqBQqAQKARmIlCCRT0MhUAhUAgUAoVAIVAIFAKFQCFQCBQCcxIBhHZzQ6wj85HcSHTE+ZQwBDvSHOFNpBDWyHmCBPGBYMArAGnuO8IcOc+jIXM6IPoR8q9unSciZF4JBLw2Nwzj3eAzAh3Zb0840AfXEAMyZ0R87DnPqyFzSBASiAzGRqSw6YPrfO9ufSYy2IyZN0Qm9s4+Z86JDPekbIa6SkEEBsr7rhx89CO9Ohw3Zv01VuPSns+EBt/hQggicBBpHCdKECdg2B0GH3VqjyDjegKPttYLc8/UYUza9Jn4o11eGe6X+6ZO90q7BJPEdALRIr53zGsRYkZthUAhUAgUAoVAITAOESjBYhze9BpyIVAIFAKFQCFQCBQChUAhUAgUAnMJgUxInYS6biD6u1t7BD6vgMw1wfOA1wXyGwnuOob4JhIIa3RVmJBEK4Qhy3kiXNay18Ye6T6lNd4UIRDwKZA4hZxPbw4igDYJCkQH7d3X+Jy5KIRD4q2ArE9PCGQ/Ip8nQfZLW4j8zA1B1NAP/SS+EGiQ+P4/15a9cTDCAqGA9whhQnl42dSjr67Rd8fTeyNDYxEkjN84XK9/6R2ifjjzinCtsFDGpq/XhLkX8M3cGTxahIzynUhxRRghZNcw90Jd7sOUljkHR33JJOc8PWzpuaIPTW+b1unaFQKFQCFQCBQChcB4RaAEi/F652vchUAhUAgUAoXAPIbAYbtv3BwR8qOZvNU5pMjUPQ7/S4WfmMfufQ2nECgExhQCmaMCgZ2r6xH8CHDHEPcIdkLD9WFECIT+v8P8/8qzgBjwj7CXhyHihS+yIeeJDMqqa+cwpDtxQ9gl1yLQbcQCZVcM877wjkiPCOIDAh65nwmuM9F2Eu3qVz6TXusT7wPCCvJf3fbKC0mVORz0kTiiTyeEvSWMd8eJYTuGGS/RgEAiP4dN/yTAJhQQSPRJGfUQPtSZ+Tt8J0g4ZwzpiaIf6iRKZEgpxyQ3Nw548GbRZxjxVuG5oh3eERm2izfGGmGEk7PDeFoQKQgqxiHUlM34jVsoKHXot7rTKyPFFvfaNqM8KlpI1K4QKAQKgUKgEBjnCJRgMc4fgBp+IVAIFAKFQCEwjyHgtw1iC7GDDELEvCcMcYM0+UYIG2KgP17CxTx252s4hUAhMBYQQFIzHgHIa6GGENuZuHmt+EyIICwgthHhVu2btxHlxIy8HgGOqEe2rx1mNT9S3XzvHeB69WS4Ie+DTIqN3Of14Foig73rbNq0uS4TRKs7wy/xECAIZMgpZdNDgOhBPNG2Y4h9ngraVUfWZ8zEBCKH5ODaMh7jz3BU2hFKiXDwulb5xM84iQmug4sN8Z9iivbUo51MIu473AlDPQJ+6xrt6ou21MWDwjWMQJL1a8v9csxnXhnw1yeCBDPGi1t1E5PcY14YN4QRLwhQ7rU+OGeM+qE/to6hoVrnalcIFAKFQCFQCBQC4wSBEizGyY2uYRYChUAhUAgUAuMAAWQS0uoNYRKBIkGQP81t8/hyXNjBYbkidxxAU0MsBAqBQmCuItD0qkBqJ8GP7CYUOGalPkLcdnVYd9g6YVb7++4ccQFJzlMg81UguRHefw3jTeBdYLsgjHcF4l1IpZeEIex5AdgTFbwnMgdEej7k9bwKkPDpWaFOggnRIUMyNb0tUpTQR2JI5qoglORmrMz1+Q66KD4T2vcIIxzYiAhEife2+qpuW9ND0Ph5S+R2aXyAw0qttvWV2KMuwg0MfGbp1WD88NMnOOtz3qtmgm6CEdHBefdBfzJh+GnxGbauI24Ig7VlGBwk6CZY6DePDPdYn7SbHhbG7PzDkc/CPfB55jjL6yLQqK0QKAQKgUKgEBhnCJRgMc5ueA23ECgECoFCoBCYFxEIrwlECcILuSM2lDjhNkRMM7mr0B8fD3teXPOu8LKwurW2QqAQKAQKgZFFwBztf097pDTCmiHPkeAIah4DwikRGAgFxAfke5L/RAtJnc3vPCiUQcIjz4kMm7XaEJrIcYQ+Ij49C4xQ2+Z9IoJ3gz7wQlCXTV+SiCds6BdPCnV4x/jsuHqVy7BWrjU2fUH0t3sKNPvQaqpn9+EwfSUWpCeD49o1Jlg0N0JDiiX6TlQhWsCWOEME0Ueb/vJqyC3zbviujxniyfccn7r0R1gnZVxjr28MbtrIfB+++yxfiP64V0JcEWB4T8BaH/VFOSGn0svDefdK3/PZsE8RSb9qKwQKgUKgECgECoFxiEAJFuPwpteQC4FCoBAoBAqBeQWBVt4KJJGVm98Le1NjbEion4ZlUlDklfjgwn245kVhZ80rWNQ4CoFCoBAYpQjkiv0MZ5QiABJbQmdEu7BIyGuE90Zhl4T9OQwhzlOOkCDhttX4mSgbye4ac3omxjbv8yZA6hNAXId0d8yKf+S58upQlz4h5BHr+snrQr3+TyZu2PSJeIBo13diBLLfxtsCEY9kTwFD24h5gouNAOCc8WaSbe2mB6Br2/8v15d2sUJdKVbk5+5WG3bGmG02Dvd4UxBSjMP7EKYpIGQ5IRNt7oXxGG+G1iIiwU0/9ct9gA2R4oVh3q1TwowBfsQXZc8L+0OrvXVj7x7xjPG+Xj1M2EZYwz9DfcE3n5fKN9VzS2orBAqBQqAQKATGHwIlWIy/e14jLgQKgUKgECgE5jUEECv7h6VYITyFRKXnhwkJYjUsQ4J8PWzPMCTJqiF4nBNeFoiV2gqBQqAQKASGGYEI8ZMihf87keaZ1FpYId4TSHvkN6J7k7CXhiHWkeJCEFnNr5xriQPI8wwp5TpEuj0hAMEu3BCCXjsZRik96ZRL8j7FBe8PZSXpJizwDLAnDMjVQBBxTXoBGE/WGx97hAhb/l+dJHsS/I6rP4/rf/smhBICv+kN2KHYoA4JN0XI4F1IAIFlhr7KvXbT6yQTYsOdwEMAci+ME7awcX8SjxR69N85Qg3BwrVEKOKIcFGbts6rhxClT4QjbV8bxtsCZuqwZaiqymnRAqR2hUAhUAgUAoXAeEKgBIvxdLdrrIVAIVAIFAKFwLyJAOKj6VlhBekhYUQKZFh32BlhRAqhRFYNkwQVufXsEC0QIlZ3Wvk5IwSMeROlGlUhUAgUAiOAQIgSvW1E4qZXBcLcMSIA8UE4qL+HIcBf1ZqbHUPubxomabN5m0CQ4aN4RRATkO3IdJ+R3LwokOPmeMQ6YhwhLvcCwQCJjlxn6Y3Bq0AZ7RMSMuyRNpHn3i36nOGK4mPPtYSM3Joigz7xvDAG7TfJduPubSNYNEM39VF0wKeME47egekN4uLMEeIzkYcHCnzhSmAQEioxhbn3JJyJRIQL4o2xwYenRIbzgp+y6nQ/tCOfFLwy9BZcjBOe57bKuVfMO1i78NZe4jpLPos4XlshUAgUAoVAIVAI177JLgAAIABJREFUjAMESrAYBze5hlgIFAKFQCFQCMzjCCA0MoGooSJ/EB4rhCFTJOJeJUyoCyGhrKA9PezbrWNW2CK1rAhFVNVWCBQChUAhMDQEmgR95phAcCOkkdj25l4CMxGZaGD+RZgjvhHezlt975g6CAhNwly5zD3henM4kv2eMOS3skSDzA9hFf/1Ya8OQ+Jnsm9kvXeEPrsu/0dGvmcIwfg4c9MXhL06tJH5JvKYggTwprDRvL798w59nRzkuUze3X65vsKZIJB770tYwApG7pPQUnDncZHJw9XlGvclPU2IF8Qn2GVejJviMzHIvXEfCTnq1bb7k6GhvKvXCCNkZD4S+/ScUV9XCGITIvF2hYcCRm2FQCFQCBQChcA4QaAEi3Fyo2uYhUAhUAgUAoXAPIwAogWpkhvvCiQXQoVo0b4hRBA0SBYEmFAgjlXoiXn4IamhFQKFwBxDIHMQ+F8TqY+0Rvz7vH6YORupLXE2rwbhhKzgF4YIUe4YEtvGG0NoP9cTFYgP6iVO2JDfwhC51jXqtsLfcR4X2s5V/jwEbK5HutsTTlxDqNDvZojA3kh/5RD33iHGlGGhmjknZkew6Mv7otXlWXY8EuDRadMn/UlBgqdFJgYntMCGG+FWYd6PxkHgIRJ4b8KfuEAAIu4TL2wSnqvLu1b9mZjcPkNkwS7zUqSXBUyYfvF6JBgRQIT/cn/kv+BlQ7hQRgir7jBj9E7uSdDOi6dEi9adqF0hUAgUAoVAITAOECjBYhzc5BpiIVAIFAKFQCEwjyOA0LJKF+mVmzjdnTYk0slhvwi7LgyBcn+EgSrPinn8IanhFQKFwBxBoClW+F/TyvhcgY/QPisMUf2WMF5v5mQiBMFCWCGr6qeEIdEJEAQHxDkC23xNXODVoJzPSc7zBkCMEyVcQ/RApHs/INqJD4hy/VO2OyxDQ8XHmRsx23EbwpzXRDNnheOZv8HYkPv6oK/N8FDGk6GUmvU3P/PgaOa06JR8u9O1xt5e9qg4tkWYceeW/WrWQYjYunEAHu4P3F7RGrv7YYNbJhWHtfuQoa4IGepy/+CUIgbBwn0Smgse/wgzzjvDvJdXbtVJfHJPPAswODrMfSEkZZ/gm3xFiRatm1K7QqAQKAQKgUJgPCBQgsV4uMs1xkKgECgECoFCYN5GgHeEpNvfDMvVoEaMaGH5ewf5cnbYd8MuCZGiGUZq3kaoRlcIFAKFwJxBIPNWmHcR0khn3hAIbavokdnyGKwTJqk2IjxDOxEaiMfmaULApq06ENrm8uXDzPFEBKS9PRGCwMDjgKiBKE/vDH3QrvBEPqcwcnl85t2RnhGZiDsOzRQrfNZX4zEOhkxvbs6pVz+aGwIfmZ+hlpwzRmNjmVOiPQH3QP83725rz1eJrZtiRYciHQ8RFdwfmMGkffPeJCTwRoS9/huX+0rIgb/xuD/weWWrAnXCL71feFys12pHCMb0TFHOs8BDxn0xBiKH45lcXR9gyio0VIebVIcKgUKgECgECoF5DYHZdT+d18Zf4ykECoFCoBAoBAqBeQCBSJyNHPpQ2OvCVmyRIYQMhNT5YQiPv4WdGnZFiBU9sbFrKwQKgUKgEBgaAo2k2ylWIKN5OwizZG7OPBIbxmdENGFCMmiE9Aat1k+LvVX4iHcCAPLein4bQeG3YeqViFu9PpvHM/cFscIxK/aR6plcW5+0yYMgPSf+GZ+7W+VbTXTcTYmjQiAhyYUmSiGkvbB+GIsNMZ/hpoQb5IEg9FKe76u9OXGOZ4Y+wckmDJRxuh/tAoqx8HRxP4SKsicswFN+DgJQU+zhzeK7NhjMMkG3z7Zzwog/vDzcG+9n9Xo/65f7+dcwIlOKKQSSzG0xvUJDtZCsXSFQCBQChUAhMA8j0HRbnYeHWUMrBAqBQqAQKAQKgXkZgRAgEChfCpNUe6ewM8KQVoiQf4XtGybJ9sUlVszLT0KNrRAoBOYSAilW+P+SIeh5PSDGnSNSIK8JCQh9XhbdrWPOK8s7gr0wDHme/6v6vFHr2hSiDdN1xASCiPZY5qdwjdX/Vv4TOIgVPAVs6k8vh9ahjjv940Xg+t7EChc2xQhCTeaMIGS4zrtobudIyvbdgxQrHEvcYcPzgXdD5qEgFAjb5Z4QeaaE8bSA321hvCcIHkQMAoV7I5E2vAg9vCXcBxj6rh6hG+WtsOmLY8QSIkbeW/fNvddP/YNvPlcTJeFuXV+7QqAQKAQKgUKgEJhHEaiX/Tx6Y2tYhUAhUAgUAoXAWEQgPCV0GzGB8BFCg+CQ+SVmCQcRwkPHIUYdrt017INhyKzfhO3fKQRUq6wVnQ9WiKix+MRUnwuBQmBuI9AikFOwyD2iXr4CYYaE+pG/4LVh14RJuIystpJ+hzBlzduEZ8IC8hvZj+h23N53CZuJHb57L2jLd+es4BdGSnghdTuHOG9umY+h7fCQv3rPtP9fbQzeX8y7C9E/0JBPxjIQQaVTx2HAyyFFgf4Gpy19zwTXmRfEPjeeFjB3LEMywdLnDJPlfihnn6GpnGc8JzI5t3vlvmjX/T4y7FWtPnipEzBOCfOcCCF2ZZiE37w38jdAz748LRp3qD4WAoVAIVAIFALzGAID/dE0jw27hlMIFAKFQCFQCBQCoxgBgoVVqsJoIEOY2NlWYF4YJln2wyE2zLJitSFgIEiEFkGMWNUrtESGo+iK65LkskoUmaatO+L4H6KOnljk8Vkf/E5C0CCOkDBWf/aIJ72JJaMY0+paIVAIFAIjiQBC2lxp7rQqnnWHCetk/kY4EzCs2Cc8/CnMynmr+ZU131qxz4QbStI7cxEJ+TQlTMg/c79yQhIhv70jHCN8eE/0tiivScJHsQFvnQSJ5sXp6dFsN5NQ65expSCQQoTvvUU7GKxYoU/eebOzZd8yn4d3Zb771JP9T+wIMXmvm+04RpRp5phIPIhQ3p/ey475buy8NHhxnBi2Wdirw7RzXphcGN7NznsG3H+WOOpHbYVAIVAIFAKFQCEwjyJQgsU8emNrWIVAIVAIFAKFwBhGABEhbIjY2cguxNR2Yciut7fOyUVxURgyA+lxb4gMBApkCRLMal6EiJWmiLIe4qTlUYHwEgdd7PRM3kq4eCDOi6ONEEGq5YY0QbQ0vT0ap+tjIVAIFALjE4HwrmiS7lbhm3+FezJvIs/Npchq5az+t/Lfivn0sjCHm+sJFMoSpZHfRAh7q/BThDCXI6+FDEKO845Ljzyr+AkWwx1BQPva6W/Tr6bQkCIGQUUfvVe827LMaAnNnKGWvCthLlG2e+ie2fS5mWwczgQoW4ouyiSvkPgT99PTxT2e0ipjIYJ3qWcBZoQJ9bjOPSVKeBbcY/3w/neNkFLe+elNM4FnT3hZzO1QWy0oalcIFAKFQCFQCBQCw4lACRbDiWbVVQgUAoVAIVAIFAJDQqDhuYDQuC4EBLGxET4EDCsvM3HqevFZTG0hKHhQEBrkrVAW6SFxK7JD/gpkykJR1/Kxf1kY8oV3BXILYWK1p7JyXyA/EDIINySLuN4IEpahqeJjbYVAIVAIjA8EGkm12wfcDANl7jRHm2+R4OZZ528K4wmxdmtONec6LycFAcLcbi4259ubu5HnGXIoiX5itMTPyGukvzk7RQ3tEjVcN9zbQMQKbXYSINIrgdcC4t37ST9H40ZssjVDSXn/4QuanEF6s6TQ4ZpOnEJ6bDgPQwIEEctx98l3m3bdW1439up9aZi2eVPatOl97B0MU8+EembEs1mhoVog1a4QKAQKgUKgEJiXEBjuFSjzEjY1lkKgECgECoFCoBAYJQiE2CD55jZhyCxkhhWel4XdHibxBZEBKYTkQHQhtQgXBI2jw5BiEntmOAmflUeIWOmJREIm/SoMGYZYkYD0hrB7QkiZGVJqlEBS3SgECoFCYI4g0IdggajOBNPmXR5xhATeawQJcypimdAg9JN5maec+ZpQbH4mBrsOGZ2ENfECqY2c5kGH8M7z2vM9BZIkxp33TnjRHAHlqY30lncCLkQcXnr67t3lf3DjntviBRGgPc+HkaXXQvadYEBIyLwcmc9idqDmsZFih/uaGOR91Bf31fuYyOX5mBLm3c3LRb4THhZELsczn8bj4WVR4aFm505U2UKgECgECoFCYAwgUB4WY+AmVRcLgUKgECgECoHxjkAIBneFaPGzwOHcsDeHESmQGIQMBJA9wmr1MGQYQgURg9TYKkwCT4QIMk34J8QJz4yzwxAmjiFKiBQIEuQSAqrCTYz3h6/GXwgUAp0QQGATC/w/ae713fwqrFOSz7zakPRyVPCyECJKeaQzsUL5/IzAZuZsYoW5t7mi3pyOQCcy89ZQT3MVv8/qE1JIe3N66y3vRL5DiBNECu8X3hbCFs7tjcDvvrRvhCOJ0t0L4bo2bOGtnGPug3G4n96h3r+rtCrxDl06LD02sm7vU9dlrhF7wpT76N1rs8ggnxHtuJ+epata10rIzWvSNZ4V93xaCGrq6viuDjGjtkKgECgECoFCoBAYgwiUYDEGb1p1uRAoBAqBQqAQGKcIWEUpDNSXw74VhtCQj+ITYVZmWpUpNwWhwvdMAOvzGmFWeCLJzgwjdiBQLg1DyAgn5ZgyJVKM0weshl0IFAIDQoA44f9IpDQi3lyKfEY2p4DMqwLxTXyQsyJzHyh7SZjQQ7m6H5EtHBTyPPMe6Ig5P5MuEy+0ZS7v5BWg/Kph5vPRtHkPea8Yi7Hz3kPuDzXEIGGAMNMbFu0YuA/tIkInscJ1+gZ3+SyIESnG2DvnXfnvVtswzwTprnXfm5tQT0Qs9zc9NJwnllwZJsG6Z8P7m3eMutSvr5kbw3teDgthpGBo7Lb01PCcKVvv7jbw62shUAgUAoVAITBWESjBYqzeuep3IVAIFAKFQCEwfhFAmBAebBK07hyGuBFWxOpa3hfIEaQaIgPJ4Zorws4MOyoMQYLgeCK8N5SprRAoBAqBQqB/BDKksD2ynEBhPkYeyxEk5JMV9ulpwZuAICG8Hs81czVh2Wp5382//ifl9cYDAVFtvmaOmb+zTd/bSff2Hpv7R9uGSE/PA+M1ToKAvuY4Z7fP6oQpr8KBbP3hxtOFR4P7SJhwb7vDmjktCC8EF54QxvD31j1SXgin3CwE8FzIOZW5KjLHB8FBWed54MDAZ+/vvPfqybBgBBN1bBlGjPKZWKK/+gKHzF0iCXe9zxs3oj4WAoVAIVAIFAJjFYESLMbqnat+FwKFQCFQCBQC4wyBRkLu5siRE4gN4Z1ujrBRwlhYoYv8yKSgyBHkBoECyYLkuLvyUoyzB6iGWwgUAkNFIMM2mWMzJBRC2zwsPwVvNiS0lfuZoyDDOyHAlX1xWArKPCaQ4AQNogdBAvmdoaZck8KIfZOMNu8r3741w0QNdbxDvZ4wnp5+RBz/e+s37LyHMqG18WeopUzU3d72+XGAlwEC37UEn+Hc2oUenhMnh/F42KTVkHZt7gXPCGMylvRscC+NqTuMt43NPu+bcvlZOWPxDKgvk6vz6iDueJbcS+9tGL4wTD4T5+VHka+EcMJTI59F4aG6SrRoIV+7QqAQKAQKgUJgDCOQKx3G8BCq64VAIVAIFAKFQCFQCHR1hViB3EKGIVes1EyiyKrM34QdH4YUQ7I8I8rXwo16cAqBQqAQGDgCzTwTyGuEc+amsJoe6WwetoqetxviWRg/eScQ3OZk8645meeFcnIhuAYx7hxCO1f48z5wDImf++xtJ7Fi4CMZ+ZI8KNL03fiI50RzIk4KKwh5pDss+koeLY+EcEspGoz0COC7Xdg6fTRkXOnJqBjhxXUpVuQxCbOFBTM+zwJhw5ZJuD0DxB1iDu8JdcLEs+CZy3BPjsOJOEYY6w7jnUH0yPBQ6Y3TR7frVCFQCBQChUAhUAiMdgTqH/XRfoeqf4VAIVAIFAKFQCHQLwItsQJJgmBBouVqTQTIL8J+FHZLGIKkJ656eFgMNYZ4v/2qAoVAIVAIzCMIpFhhOMh2BPHtYYhl86oV7xkWCIm8bti1YcIDCQ+1fhhiGlnv2gzvhIBG7GciZWJFEtXpXZEQ5vG5AWnmUxho20QY5j1jjBkK6tb4zHtAngZEu/cV74beknZ3ao/Yk6Ga2vt1bpx7adhwEff62tza2/NduEXChjEQHng+2Hg88m70XAgFZrzrtfBwPgUP13lXew68x7Up3BWPCosPjNVzluJXYqduHheeJdezCeFlUaGhWjegdoVAIVAIFAKFwFhFoASLsXrnqt+FQCFQCBQChUAhwKsiCS0kSHpXZEgNxAlCzcrOm0Og6MlZUbAVAoVAIVAIzDYCGXYH8Y5kZ0LxyUOBkEYuI47Nt47xqEA0O2c1PA8D3m3IaHURLszfyiD0XZve/447354o2nECwNwI+zTY/5uN6d7GGAEPw0xc7rvcEbnBIsWLzNnQON1Dyl8TRhSCxbfC3hWWXg08GAhFOzXqyev1o+n90Kx3oJ/bcfB9tdbFxtH0fFmzQ6U8TPRD2QwP5X4SM7yjXe+7kFeZ38MCBM+PkFiSrh8bpm51EUc8U0QcHj0p1NSChIHe0SpXCBQChUAhUAiMQgQG+8NrFA6lulQIFAKFQCFQCBQC4xABxI7VpFuFST6KpLDq8vrW3grX7cP+HDZlHOJTQy4ECoFCYNAIWK0eF7NMjG3OJTwIAYVE5jmxVtiFYVbD86yQVFs5RLM9EZmgISQfASNzNiConVMuw/0godNDjujRvg2nWEHQNpaR3ngXGBcMEfVEhwyf1S7AwCM9SZD4zS1DI8nhQJD3XeitM8K2aBWUv0nYqE4eG0MVK5p9aXpSNNsythRg3G9CgvHzIjFmXjbGTOwiuhhv3lMCjU1ibYIYHDI/RiYENzbjFh6L16RnicijnHd/j6dFPLeunVH5LJq3rD4XAoVAIVAIFAJjB4HhchUdOyOunhYChUAhUAgUAoXAmENgxowZE2LrWY0Zn3tW4f7q429Z5KF7bn/zjOnTXxFfhYhAlCGETg87PGzzsF3CJkyYOPHwpVda64jXfuLbj0c9PQRIs84xB0h1uBAoBAqBYUJAouJetmaSbcQys5qdOJwhiV4dn5HkiGlzs5wWxAxkNVK6O4ywgVh3vVXyCOb0MDCvI5ntEdlIegR4ihrDnXORcJCE+lBDTAlhRBTvbTN+ZH0zkXYKM95DzTwWxp542zsHhwzBZK/v9gh9mzouaGFG3PEePCLsrWEr9tGvgZ5yD9KzpnnNQD01XA9j4xcyLJOpEypY+waDzPFB2IKD5wbGvntOjN+z5rMwUeeEedZuCrskjOihXaa+Ei0GererXCFQCBQChUAhMIoQKA+LUXQzqiuFQCFQCBQChcB4RSDEg05Dby6smNAq00OenPXD/1vk4fvu2n1C14TNQ46YHPZQKBBBVky4aYGnL/Sz1Tbf/vZ/XXjGffffdtNKoVYsN2P6tF3vvvGaR/5z9aVHRz2IDERP1pltd+yEkyFyjNdbU+MuBAqBeRyBWIXe2zaj5WHhvPkR0U+wQDZnuB85GeSo6G6VMVlaRW+ORSD7f9N5QoUNeS3psnK5gj6J+6YHwEgl1W6GXxrqxN6XWGGsxuydlaJLvmNggGTnEcArhdkIOT5nvQh34bWEPXIMSe+7MsahXsKEvbJMcu52z4xW9bO9y/wQ7Z4ZTQz7qjSFGkKKawg8nosUXPLa9LAxDveEF4VnQkiwzI+RAo/zBDDPneeMd08+T1Pis/e7fvds5WEx2/e8LigECoFCoBAoBEYFAkP9kTYqBlGdKAQKgUKgECgECoGxjUBLjGj+LkmSx2pKx3u+33nDlQvecP7pS1x95gl7TJv6+OtCjHh6aAmPdE2YeO2iSy2737Krrz9ljS13fGShxZea8NhDD8x3/i8P7p5y0Zn7TX3i8edPnDjxxqVWXHO/8LJAgKRogQRBIiHVfM7wEwCdKWCUYDG2n6/qfSFQCPSOQD8eFuZGZLkQPchxHgMI6A3CiBaOm0+VscrfCnmr4ZHSSOV/ha0SZi73mQeG80hpc7sV8Qh2NtzeFKPxtmduBSQ73AhATQ+MZp+9jxKfFDWIFsJr8TwQFgnu6ZXA88D9QOgPV/inZuinweJpnO69Z0BoKGPiHbFCGO8c3wlUngmb8cDJcV4mnjnvY9d7RmBH7PH8COtFGPtbGLx4WsjhQdghkEwt0aKFau0KgUKgECgECoExhEAJFmPoZlVXC4FCoBAoBAqBsYpALx4UhtMMgYGI6PF8CEPg5Apc5XriXJ99+FcnhwDx/icefVjIi+kT51vgwfknL3iDkE+v+ehBZz3zuStYkZnlp06b+sRyv9t/763vvum6HePgw5Pmm//6pVdac78tP3IgEgYhkkm4s60MYZF96YmDneGoxir+1e9CoBAoBHpDoBfBIkM2mXuJD7wqiA3IY/PkpmESICOakc5XtY6/MPbmV0SyVfJWuyPlM8QTkh2ZjoDXBlLZ+dG4EQCEvuqU/Dr7m+Pqr/99hZ9q5rFAyvO0yBBcvdWb+UCc994kDhExMtG5dyERKIUOydBXDiN2OE40Gu7NMyBZtjb7wsU9J7wQL2ztydSJD543zxARQzn9JV7AKj1RCBfquTzMNZ67f4bdEAYLz55+EC2aixGGe9xVXyFQCBQChUAhUAgMMwLjYRXLMENW1RUChUAhUAgUAoXAIBFoihPNGN1ICKSXlaJW8zIEFkNs+b1i1eiSt/3zb+tNnz59ywkTJy04/4JPv2uRJZ9z7gs2eOXP3/D5w84OsUKd6hB6omdVcAgUk7f4wFfPDo+Lq+PzkiE8rHH7df9472MPPiBUhzrVrY1sL9tXjz7p2wIhuEyS86LN5MHosdoKgUKgEJiHEEivNoIDopghmc2JCGM5Kl4URsBACP87jGiBMEYcu055hH8mS84wUsIbOYdQN/+OBHE+XLci83S0hzBq1t+bd0SzDI8UxHr7liQ6vAkVmcfC+6e/ehO3JP/dk9XCCEoEifTOyHZ5uWgnBY3ZwUjfBrKtGoVSIOmt/wSFf4TJvUFYyP7zirDpr9wfrl8+DBZyZsDQM+OF6znM3B6eJ2GheGt4nozdM5nPrWdxYiO02UDGUWUKgUKgECgECoFCYC4jUDks5vINqOYLgUKgECgECoFxgkCKFYaLQEA62COzkDSEgTyOUGFCPlhF2kOQPXTPHV2T5l9g2QWevvCDUx979JEQIB5basXVf7bBjvv8Jz5bgel3DSJD3T2hIFz/tMUWv/MlO73v6GvPOeWhyGmx+IN337Hi5acetcF62+7xr4mTJlmhiWBBbiA+EGwMSZIrOfUrQ1TkStC8baVWjJMHuIZZCIwTBHKuRhibl82NiGAhdoi7m4WZt30n9Jorzb/CEAkR5bi5G3GMPEekq0u+gZznzbvI51xhP1Avhdm5BdobrlwOs9Nup7K9CRC5eNBeiCR4JuGvHqKD91A7+Z85H5SB9dKtRl3L0yJzgngPwry3TXhEQsBL+xmgd+uUMO/U2U3m7T7rr2fm0jCeHp4x4oq+wSY9HfXXuVe2ymfC7kz+nQsKlOFlYVMGBvKkwElZ72v1wlOdtuk8iSo8VAuN2hUChUAhUAgUAqMcgRIsRvkNqu4VAoVAIVAIFAJjGQEeCdH/zEeRCTWRChnHG2Fh9SpvB8SGMA5JMiEcnF9mxvTpS9102Tm3Tn38sQUmP33hayc/fZH7F3/eioeuv/2e14dYgaxBWCBFkBgMsWKlJrLtieetu9Hfn/7MJbvOP+rg9f97121r33L5X5+x9ta7LDVx0tOURXBkDgvhJ5By6kT+IJGEA1EXEohl2KjMeZF5MMbyraq+FwKFQCGQnm/maPMfwjdXrZtTzX28KK4Lszo+KOCele1Xts6tFPvVw4gF5nLhodRl/iRSmCvN6bwtklSHen/eBIO5M5kPYTDXDvc1/Y0PLt5BTbFCHzJklvdl85zvKXZkMvPss+PeWcQg1yDse0uS7V7NTFDdz6C7O5z3/tT39n43izpnEYB+8ZjwrvfOz/vj3Z3il+fL8wGLDKHldwDhC4aOew6vD7OYQYgrgstlYX43OOc6iw+U1T+flbE9EaLFtBItWmjUrhAoBAqBQqAQGMUIlGAxim9Oda0QKAQKgUKgEBhrCLQEiux2ihV+byRhk6EckkRBWhAHxDXPkA9EBgSXa3haPDh92tRFnrfOyyddf94fFoj8FddEGKijVn3ldrdPXmgRq3fFzEZ4IDsykSsSBnmBQLsx7NrFln7uefMtsODDEydOWnb6E08sPO3xRxcMD4unhdeGlcFCTiDUEDtIDsljkXVINX3RX6s2kSLGkGE2euJjx7hnES0q58VYe3Krv4VAIdBCIMMUmQsRxQhnRLM5ENmMLCdGEJjlLDAvnhuW87i8A+lVgaRGIKuTEJx197XqfzhuBMGEtZP57XWnwD23PTHg1FvYKe+0FPiz/+0CiPcdnN2fC8POCtsjTJiufK/1hqv3X19b05ujvdxA76P3uPexZ0k/JeAWPsq4jwtTz7Zhfiv43SBxtnLdrTIpYhhnhnz0zlbOogL30W+AFH3WaV0v/FR6W6anRz/DrdOFQCFQCBQChUAhMBoQqKTbo+EuVB8KgUKgECgECoF5AIGWWJG/LRAHyAjkfib+9NmG7LKqEqll9SRCBiFmxaTkmVZNIkkIBstOe+Kxux66967nTl5o0VumXHTGcxZ+1jJTl1l5nXtbQgOyDOGC0EFM+GxFpVXACArntdcT6mn69GnLXnzsD5e7/7abl3vB+ps+tPhyK1wauS+IJcojPGxWbyI81GMVsTrUfUvrGBLPRrTQBmLMZ33OWN+VqLsFUu0KgUJgdCPQSrrdDNtnXkb2yw3AG8Icbp5eN8zqfXO5udZcmF5xyHLEsWt5VphPM6eQ+TGTSQOjP5J8dAM293vnXeN9mblAkPdE9hTf3R9a5IDlAAAgAElEQVT3yzvYO6ovD4hOo1GvNtw378Fm3kttEZ8Gu3ku9Mnz4vkwjuyrOrXrfew3hOPa03/PoH4RMtIbk4Dh+fT+V4/cF+rk8aMO5wlofw+TbDzDQ80oL4vB3r66rhAoBAqBQqAQmDMIlIfFnMG5WikECoFCoBAoBMY8An0kl24m0/bbIkMn9SS+DuMxgVBAPiA/fEcsiDmNUOABIXlrJtkkZGRs60mRr2L+Rx+45+HwWpive/3NlogcFgvGZ2KGdtUhJAmSQ5gScbERG+J4IyqssJRsdOOw88K7YvKLd3jPgnfecNUtTzz28CKTF36G67RrJaqVmxn/GrlGVLkmzMphK0QJF8QNoTacy8SeCBSETiYBNVZeF46XcBEg1FYIFAKjHgFzWOatMMfJVUBINldbxY5gPiFMGCE5DzJMUSZCJlKYdzOHkPnSnOp7ihWZE6MJBs86c3aTFB8psEZTXouhjDE9V+yJFN2Nytyn3IhLSHqk/kC9IVzr3ep93QyrlSGavK+9xwe78FFfmpvfA7xAvE/V673tefMMei78hrA1E5R7TjNUY4ox3tOEmr+26psSe8+d3weeRWKa93aGgWz3WmnrVn0tBAqBQqAQKAQKgbmJQAkWcxP9arsQKAQKgUKgEBi7CCRZ0Z6jwm+LDK+R+SmMEpEl5MUaYVbkIlqs4EVWWa1pJa9jSIuMRY2ImDbf5Kct9Mxll58wYeKkR+ebvCAiI0NGITKQFAQSgofr1YXMQEog2wgbxAgrgREc/9aPJZdf9ZHIi/Hi4NL0AYmRq4O1jQBSt/avDTMO11ttKvwU8eK81nUEE+XUnUlAkWJw6clx0RYuamaS7hBd4nRthUAhUAjMdQRyHjd3Io3NgQhjq9QJFuYtXmcIYHOq+Zwhn835CGdlzOdZ3lxqbu4RcFv1dfrfU339kcfZVn+5IPoDsj30UzPckf6b42fXG6G/NjudT/J/dq/Vv/RUdJ9sSeT77P3J0yDDSynbW6gp5YkPRPj2rRMGnpHst+diKF4W7e15TjxDthxX00uT6OLZ8hx5/3snM89OChfGod/dYa71jvYuVsaz7B1vDDw2poVX0fTysuhw5+tQIVAIFAKFQCEwShAowWKU3IjqRiFQCBQChUAhMIYQaHpUEAmQBJl4E/GAcLCy1jkEP5KJsMBzApmCmEjPCKt1rah0XSbWRIoQFuyXjdBPN4dpI1fnImWs5kVCJHGRsdW1hUghOKgzc1o4vnbrnHonTZg40TWu50VhIzg4R5BwPbLj1WHG47OVxPqPBBJ/O4k9/RGT27VWcsICAad8huRo5riYKVq02q1dIVAIFAJzBYEgbs1R5kpzrHk7Q/T5zhDe9kIOmavlBTJHmi+VFcKPkOycedPcThjI+dC4/M/Z1/+dzQTcnXBQt7bM+f1t3i8DTbht7r8izCp848sx99fGUM8PVq327kmRJb1Fmt59CH33IsM4NXFA+hsf0QPe3onI/9nZiPv5jhvIdf0JM3mvmrh7htKrQhs5Pp/TE8c4PWfpaalPxgIfeS0sYFgzzHtZXbmAwTs580892krA3RR8BjKmKlMIFAKFQCFQCBQCcwCBEizmAMjVRCFQCBQChUAhMNYRaISDSrEiw3dk6CZEQXcYwgsxknkdEASIEcfElUakILhSxEAyIPyFhuIJYZWkvBEZXglBgpSw4lcdPhMNEBAEDsKAPmR5YoXvCAxEhbr/FrZZGELKimB9U0fGxXbc9Sl6+H10WZhVvVkfooRIog8SzSJaXI9Ayzji2lW/MWh/SljmtrBPr4v42NWKGOVjnChviyeBqK0QKATmGAJB2DZzDpm/cmW9VejmP/O0uewVYUhuXhbmVCSvudy8aB42D2b4J+fNvekxZ75FXJu7bc7LJ0DAHihxTzTRjxQsrLbP+trxGqhY4TrzsveOud91ObaRDE/VVxLr9rF0+p59S5GnWR/cvYMI/ulpqDzcvPMyiXrWC1fv0HbBCC7yPnW3dSCTZmcib9/7uof93d/e7pX7kMK+59LvC/1Mrwv1GpPx6quxOedZM0b9EwpS7oqrW9/TM0Wfve8ZT4sJ5WnRdpfrayFQCBQChUAhMAoQKMFiFNyE6kIhUAgUAoVAITDGEOjxUAhDUCE8ECLIBMS/TVJNx4gRPiMXeCQojyywMhL5hEhA7r8oDOnvs98mylshyTsDsUX0QGBIeo3g0GaGJkGsTQlDOmXuDHviiDjr64VlHg31EEAQHOoSnkp/rEhFgAkhpb/6ZsUtEsuYLgkTXmL9MCQJr5CMoW3lL7ElCRXEifEROpBG6oeDsBXq7S/0SRSprRAoBAqBkUcAUdvysEAK5zxubjSvEWiF6hM27+WtufD62P8+TH4Lc5z50ZxtXjPPCTFkM+8pa1503Nyfm7nT/D47W3vYouYK/Nmpx3ukGVaKANO+DacHnDkftu3/czf7kWJ7X+PwfoRxM6QVjIVXtPde9B7SnvfOaWHedxYHbBHm3hJ4mv1I74dO3i3uG6/I9i09btzPwd6DgdyvXIiQZY2TV48+EyPgkL8V3E9jFYqMyEao0Hd9JWB4Js8Ps3DBQgfvcHi4L4/H30B5WAzkjlSZQqAQKAQKgUJgDiNQgsUcBryaKwQKgUKgECgExjAChAS/HRAEmZAzvSf885/JsgkCCP/0tlAmV9MiZ5BVSCyhRdSD+FIW2UKAQCqIkY0wU45AgBxxLXLFceeRFNolLCAw1JUeH4QKxITrGRKHmNAdhmSzz/ASRBEkCGJOWSuHNwwjbmhDvfqXyUGROVax8vpQh/FoC8kiHAXhAyF1cZix6LvzGevdOWMZTmIsqqutECgECoGBI9DysDBnZiionN+RvduFCavTDPeHODZ/IYXTw43AYY43F6rLnGkzH5orlesv5NPAO/1kycHmshjIdf15BcxOX5tCTV6HLG+24T2Q74JObcNfv5t5JdwDG8wJ7t5f3jUWASDtXxaGtGfePer1nvNu9t6y9ReuqTdBgnDQngukN0wI9X3l0MjrPEN+I+SWYyU4ZF6VTDSeCwSUhY2xdbfG5jdEhqn03rYYwjNsEcHhYYQfz6T6ezCLv4FHy8Oit9tXxwuBQqAQKAQKgbmHQAkWcw/7arkQKAQKgUKgEBg1CDRCPrX3qUmgpFcF4t5vCKQJz4buMMQMIQAJQmBITwYrcZEoziuHmJgShvBCUCDuERDEBCEorIJUhxW9iBUiQhI2uZrXcYaQcC5jeSeJguBAkiEunCOIZHJuZIW+6D8yRT08Oex5WTiP+MlVsfpLfHG9eNi+wwGZ4zuCxPU8OrTPk0Rd2n5lGIJkSpjVxvqr/szj0fS2KPEigKmtECgE5igC5qkUVBHbSFzeDAjeJLYd42lhM9eZUwnLOb+aG83N5uJM+qwuQq45rzexIufZOTrgtsaQ/QTvOb2l4OA9433VPv9nziPYwbk9RJXj6RngMyFCncQB9wr+8HXMu9g727tWuMW8r4MNe+Ud1tv7qv2eDkSsgL13vzrT84bwn7h4L3u+jMNChUzmns8aHHoSabfGm+GqjJN44zeMe/ySMAsXWC4ggJs+l+eju1BbIVAIFAKFQCEwihAowWIU3YzqSiFQCBQChUAhMMoQSLEiwyf43YCAQGYhD6xS5InA20DyUsQCc46tG4bgQggg7hELyHqhKRBZCJR/hF0U1h2G7EfyO0eoQEyo76yw9LZIbwr18YTI8FNIN58zEfd1rX6lAEGkIIYgM14VZiz6gtRAuBmjuvVR3fqgrL6qO4kXfdIOAkg5ggw8kHiXh1ldrM8wQagIO5UxtZEj+odE0Y7xw2Z6CEaw7lW0qBwXgU5thUAhMGwINJJtZ4g/85b5iMBr3jM3Z94Ac9k5Ychxc6P5ypxsvjOXmdeQxsRnZZRXT19CLLK+v82cmbkHvFO0YS7uLX9Ff/W1nzfnt4eJmt06eiufq/+dbwr/mTOieazds6I/MYFQDhv3DPaZTBvJn+8q572X0iPQ4gL3yz3Rt8F6veQ9z3aanhoDuaed8Hpx20F9zdwcRCWWHpbuF+EiPSq9y42R9493rUUF3v+8K+DkWu9mz4zvzuU96Hn2428hMXlK38L7orZCoBAoBAqBQqAQmAsIlGAxF0CvJguBQqAQKAQKgTGAAAKFITUyzBLCADmCTBBeAgGAMEGM+IcfaYIAQmgg8f3OcAz5cm0YggPJZQWvY74TKTLEhNWVrs0Vj+k9oR/K5GpdQoE2mc8EBdaMa+1axIW++6xN8cr1w5ZhUBA6Sbwge5AbVqFqLz1AjM3YiSgEjvQa0VfXGmN6YRAj0sPCOMTPtrdClECiDkII4g3JAofmCs/ytGjdoNoVAoXAiCKQ87s53pxl7ibsbhVm7pYTIBMaE3uJz+Y+hDFhIhNhy3fhmPqIv/bmXoKyeRlJ3Ck00kAGl2KFst49mXTbd7mFhP4b6nZBVMCjb7i3dtEhBQzvEudm9/9w98LmHQF/Ao53cIaUIqKnmOB+qN97rOmJ4Z7kfe803vRW7HQuc23wTPSuZNoczhBazXYTPx6bxpM5VryfvaeFlDR2z1iGnSREeMd6D/ttkqKM9z8sEpcUMjy7ypSHRac7XscKgUKgECgECoG5iMDs/lCai12tpguBQqAQKAQKgUJgDiOAiEhiP4WLjFOOgEqviq3jM6LKP/08CzIBK3IAsYBEQegTABD36kV+IFKcc636EPoZ/9zqXCQE8oGnBmHC7xbXKYtg0zekmfaQ/syGxBFyCtmF2CEOuJaIgrDRL9d0h6Uw4ztCSP1IDJ8JJEgPZdRjVaf2rOLUNrIkE3nbZ5+17zsSzKrPU1rXI1hcB0NjMP4k8nLlaxyqrRAoBAqBOYKAOdbcbk6Se8eclvOeY+YyIq95mzjAu0xIHYKEeducaG523Nxq/jTHpVhhEIMVK/oDYLUOBfRH27OzjYRY0al9YgAsvJfaCfIUM9LTLkWIpheEe+U6GNsTylkuFtCm4+ogJKSHgnZzQ9r3tfWVmyJ5A89Jc/Pe9swQFAj0hC/fB7Nln12bAkl67Bin+2vTB+9oY83wWcIuErQ8sxZGePfmbwjX+n1gfCmqeeeqW5n87TCYPtc1hUAhUAgUAoVAITACCJRgMQKgVpWFQCFQCBQChcA8gAAiAAGBeCAO+Icf0WJlohWOzRjbSATESYaDQjQQBZBcyCxEPRIBkaROZBdhw14eCJ4PiBZEmHJJwiA/MsSTOgkC2S+rKhEO2s5VlogS9eub87kKlVCRyVaznSTVjCljcuuzPgolgexQn9jaBIrsf65OhQnCzCpkdRI5hJrQrtWdiJH8nAm2CScwgqHxJ+GinwiTJKniY22FQCFQCAw/Aq1E2yo2l2W4IHOUuSmFYfMgsVgZc7DExebEi1vXmP/Mx+YwK/29JzKRsbm2e/h7/pQam0mo8+TsihXtlbYnfx7qMIgFGULL/93pNdAejgn+Nsdhnu8Gx7wX8tp8l6R4nuUzf4Nr4e8d6H4mHs3QWkMdU/v1xJHceDIMZWv3SknRwnNJ7OHZ6d3KvP8z7JV3rcURxpw5rry/vbs9nxZLKA8fz7Hy6vYe9u72Tk5PkfJyHModrGsLgUKgECgECoFhQqAEi2ECsqopBAqBQqAQKATmIQSQBogQhBBSCjmQ/9Qjr6a0/tHfPPb+uUcMCHNkQ/p3hyFpMqQSMj5DhKRQkCs9XUtQsKV3RSYK1XZ6bCAUMsm2z9q11y5hpEkyZIgqbWnHikrnlUVKqPPSMGLDq8O0gwxRHvEj5FUKH/qn/0mkJNGhDYm2M5k4zwsCC2JF+BREYHqDIPtcd16YlcjaQ6LY9C3zZuT4M4RHq0jtCoFCoBAYNgSaoq/5i6CM2M5wQN3xGQmdnmxIYnNt5o9AAiPMzVNp5jr1+t9ypEIEDRsAfVTkndVpy5wHzjW9APrrk3dnek/05WnSnvshFwd4R7k3BHN9QLb7nOEPvZfcF5grl54O6b2Y3hb5fmzmm+iv7wM930xcTjAYrvwiniXvSb85vDONn+ekseXCA+9MoSTTyyQXRbgONn4byCMljJVnWP+8iz3rzsErPTszz1YJFgO981WuECgECoFCoBAYQQRKsBhBcKvqQqAQKAQKgUJgjCGQRJN/9DNUEnKAlwFCSmxzZL9krEiJtVr//CdZIHk2ogUJgPTPME+Z6wKZ0AwXkatD7REIWU8m1LbCN5NYIyCQaEmMETUIKulN4TtSwnd9cM5KS8RGrqxEWCinnpeECSuRIa+MWTn1I4Dsr2jVI/QVwkT/X9AaQ3p1uC4N8aefQqjoQ3cY7JJk4UlhTAgUwsXvW+cRKIm3uprkUnytrRAoBAqBoSPQ8K4w7zEErvnOZ8Ls9mHmb/OYc+YxXhVXt8qZy4jAyhMyCLXmL/OZeTw91tKjbXY7TVR2rbncXDlcW67UH2x9TY+I/hJit7fRLJ8hm3Ke9z6ypWCRgoLzRAliPnHcvfF/e74zHXePmnkxnGt6cHjXNre+iPimIDMQjJrCR5NPuCouXjnMu9LzMdR72AwtlWEpCQy8GT1zvDMz4bj3uvIWV+iH797X6W0Ja+dfE/bTMGNOr8dcrJC/FUq0GMhTUGUKgUKgECgECoERRKAEixEEt6ouBAqBQqAQKATGEAK56jZXyep6hltwDPkv3IO91bXnh1lpi3xH7EuM6XeFJNpWRLo2k3UjVRAuCJZMxJ1kWIZCQnSpDynh+vTaQPLbkgzzGamQ8bvTQwE5QRhJ7wpkRIZY0t/0FEmhQz2ItyR5EFrCU2U8d/3cOAzBsVFYhr0yliTj1m71Td2uJ7o4j9Qj1sBNXG118cbgefGyMCtCM9QWwsR1+p3Ch2r1PcNutZqpXSFQCBQCg0dg8qFdM1qiRVOcVqEweOZcgrS5B1luXicep3ghL4A50zlCrNX/64eZM5k5z1zX7i2Q89lAPC/Mi9pvJtce/ID/d2V///NOaY0tRYHhaLNTHU3hI8M3NfNZpMdKvmPg4d2YSafh4hyMMtRUCvf67lzi3MS7P+zbQ1T1N/5mfc0wXBs2Lsx72V/bndoyXmPx/kzPSu9J707H8/3q+czfLM7BwMIEool3KgHMvRVuMpN0e8ZfF8Yz5OSwFHkqJFR/d73OFwKFQCFQCBQCcxCB/n68zcGuVFOFQCFQCBQChUAhMAoQyH/akSBIeHsiBEFAGCWrE18blmGbECw8LZAAyiETcnWo4SBCkkCw2lKdmZw143T7PcIy74MVlMplUkyEBXIhE3UnSYHIUX/GXU9RA5mTeTTUa4Vl7vXXOaafjqcXhhWbOR6ESIbwSOEFNkku5apibWe4CuKD8RMyHBMGywpQdSJbkHvbhMlxcUkYkcdxq0Fdpy+1wjNAqK0QKASGH4EQK5qiqDm7O4xQQYg2x5vPzLfmLyvkrWRHBKc4y/MhcwcQk4kWhGZzo3nXHJyhiwjAVrgTlWfHK0Fd5tfczJHqbBcxMlyQcgSU/hJKN6p8ykfj9z7pb+vPU6O38ylAwyeF9HZPxgzF2C4eeNcKBcWbJRcWEPyV887wfnHPvKea4QS9z7xzHcs601Njdu5Hf5j0dj6FhtkVQ9QnTxYvEr8V/AaBwUlhFhEQHrrD3DObc3D3Ds13e4oonh2ih7qYd7Tn17PuPggBpv4pYZ7lxKXCMrbArV0hUAgUAoVAITC3ECjBYm4hX+0WAoVAIVAIFAKjBIEZM2Y0V0D6bYCo5yXgn39klc/IAaFBCAfCPVlJ6Vh3GKIHOeKffV4OBIckUpBKSDDeGUgnRL36XMNrIUkm4kUKEYgyZL+2MmE3sspqyfRMUBfyLGN2qyv7rh+IGaYd4yOaZNiLFDOSnFAv8g1Jh2BD/CQmGa88v2csdxhp3zWuVyfiT/kMhYUUkZg7vU2y/UzK/eJWu8ojS/Rf6BVt6LsticDW19oVAoVAITAkBMx75iJErXmZUGz+RhKbz8xhjiOIzWsEiZyPV4zP5mLvhZvCEOfmrRvDzIPmc+eJsObDoYgIOUj9a25C6XWHeY/Y0uOurdiAvuac3Ewc3bxQ3Rn+z/H+/nduP5/5FlwLywz/p90mOW6+b4Y/avZBHcQlhHx6DnpHZVv65z3XLkJkmCPvKffQ1sn7ZUBADaAQrLSVOak8G4P1lOEhYWvel83iu2cKjnBQv/cmQcJvkVe2MPLZ4gp4+axPnlV1EdEuDyNc+E5Mg7vfHHlPSqwYwM2uIoVAIVAIFAKFwEgj0N+PrpFuv+ovBAqBQqAQKAQKgdGBQMaHRjD4Bx5BYnVikv9ICOQTYss//PZIkEywmd4TiBNkANEC2W5lqLLKIVYQYkib3OeKU3uiAzICwY+MQPYjq5xDIqQHQ/bJ7xhED+JBGZ9T9FCWCGEFJQFAP/SfOJCChVjXSUh1x2dJOLXnvBASGaJKmfS2cE2SPsQNKzlz9ax+Iz5ssHONtrN9uS2sklUvTwvjIF7YG0MmN1c/ocd4muFCWlXXrhAoBAqBQSHQ9KAjMJibzZkXtOYyuX3MXeYg86/jBGpzlPB/SRhnGKgprTnK/G4OQxLbI4+HczO3ereYi827SWhrg/BirjRnpzecYwP5P7e/1f/qGWw+gxQrMuygPqYHRrNvPjfFBmNNT0Xjy3dk5m/yTvBu0a/83BTnE/f0QGgXfIbzvjTrglWKFY7nu9Fzlp6D3n/N/BcD7QsBQh3G65lcIYxg5blrhpOEpXG/NMyCBzjCs7v1OcMv/j2++73hWXJMH/Xfu3owIawGOo4qVwgUAoVAIVAIFAIDRGAgP+QGWFUVKwQKgUKgECgECoExioB/0BE9iA3/4DMrZP2jL7Y5gp2AgCywstZqWysbkequzbBMSRIlqY+csFI3Y3ATNZLwcp12hHNIsYSQoU5EBw8OxzPhqM+usZJXva7TZ8JIJnrNkBiIIp+V0ReEnD1Bwuf0XkBoIEHkldC28hnWxPidF+ZK/TnWDGmlnGu1nytfiRXqcFyIEuQNvJCC+q4+Qk13GDHF7zDYWiEq9Ip2En/3ApGSgkp8rK0QKAQKgcEh0MhdkSvykb3moDXDzInmGyQwstf847z5m2DhPA878zHxF8HuuO8IYuftzW8jsWW4Ju8Yc2JuCGZ5CMz35vbsk7med95wbHAxL2t7oFsmxG7iATN9h23mJ3Is81aoO8UNnzO0Yb5f8z3nPex9kqEG9S/DbrV7WWivUwJ0uKUIP9AxDaZchqtybXqQDEYQgIEx+h3CS8L99Q61MMHvAeKaZzl/D2TCb5hZhOH6FDK0f16rDs/+hWGedXUTLpwvz8bB3O26phAoBAqBQqAQGEYESrAYRjCrqkKgECgECoFCYKwh0AoHheRAxhAKEO5W0iJVCBO8Eq4Jy0TaCBCkFs8ASVl9VsZvioxfLqcFsiVjS/9/9u4tZr83r+/6TDzgxMQDT9TU9oFCW4FShj3MADNA2RXa0to2pWmNCUmrJx7oifGsJ3pgYozRg4Y0WqOxQkSqUgq0DJthGAaG/UYQ5hlAo2nsSeMGE+fv9Xq83/+u/5p792x+z//3+/++K7ly3/da17o2n7Xu77XW53N9v5fykfLIm2asIhaEasijwv4PrWR2rvORMpEPxTOXN4+KoG72qd/aIMmHsCBSJESYkZk3CFICuYWsKMSGzxbO1hbEl1mdBAeEz99eST+ERCG6IIl4TOijxWhrF1EGGQRLZAnCplBWZgW/ZyVYFAIKnvBDrvEGUe5PH86vv8U8X7tnGwQGgUHgQQgkLrN1CHWENfvDfn3dSj+30q+sxPZbs4LHAlIYketcn+wd28imJSaz2ewfW3vJY+FBDd+dZGZ8Gxv7TSsZK9h8woW2ILJt7Hzjx7nQUXlwOIe99dvm0ziij9eEt8p7QH72Oy8In9v3br+1M5E9zwv4GW8KS9Q124eLyttCOYj4zolsPzT/zZCI/e4TJq5t4ab2xx/6u3ZvhZj69NAyneeZwJipr8Zn1+QzVip0JRwbJ117zyfywsl47Nr7/KWVPLfcrGR9qdvDb8f8J5qwkKD0mDbPuYPAIDAIDAKDwCDwCARGsHgEeHPqIDAIDAKDwCDwKiOwESualUlQQAAhM1rA0gs8Ap0nALIdYYVo+YKVEEfNPEWCIbGQWmblOsZrAHHf4qg8DVrY1axGzyFIA5t6I8mQM0gOhFprUORRkSjSjFu/HbP5VH6zT3lH+K4cJFwzO7UVgZGgQiTQTu1HfBFnEBj6JvY1PMzuNCsTBo5L9iHEYHS7knJsiCCkSvHg7YOftiHV5IMhgtD5X7VSi4aqi0iCKOOR4dqsS/XGWQLl3e9+yKTVQ2vnYxAYBF4HBBiJwg+xhzzAzE5n93w3Sz3ym736tpX+3krsthCByOFCQbFxhFt2EgHMZisLcfyYdRIuLWrtOln7p0171J3HALtcKD22/HYlAov9+sG2HtsaT/Jq8DuRgaBzamOXjREJJey79mmXcY8dh3meFpHqjldHIk+fhRiMPFd3Yak637U0NiTG3I0TKxlPjD2N6fuBYbsmk2t9KdyVcbwFrM/A8Oah2mGH6+DeUk/radRux++79ojyXMt//dDH+s7jojHVPsnkALhrv4kAxm33pwkHnk/cv465dwkfJk8oozCY7sPZBoFBYBAYBAaBQeBtRGAEi7cR/Kl6EBgEBoFBYBB4uxDYLLSNQEBwIDIKPYH88ZJPcEDqR7YjYngpWMNCSAbxnxE0hTIiVjSjFJkvr9BIwivx2mgWJKJL+cI7yUdQUHezWAthgTyw36dnlkilQkIoD9HgfCQFQiOSSfmd2yxLn/LqKxJGmc2+RCwhtWDhPKQGrwd9UjZSg7DQbFF1IcCQYvqgT7crIYwSFwgjyv+xlXhzOIakQQwSI1qQHMaugzJ+/ZCvGbPF1V67J0wFEGYbBAaB+yFwCAcVwc32sd8ECMIzW0eU/tqVWqGgcuAAACAASURBVMyYgMEey8smmdHebH/2zdhwsxKxAPlb2CQ27NgWUX6p4efeTdlJdnFPwptRz55qKxvOJrOtyvqclSLvCyV4LESSdiW4522Yt8S5Niu7BbGVa3wxNigDNmb6a5O2w9YY0BiSV19hoPSrBaXt0/6td526ylOfjIHabYyy71iYp20/9iGj9lgaT+HUdh+xonP0S9thYKxuAgIMEhnkvU+ILflhB5992DG4w5kn6Fdv6pNXfzw3aIP6e17Q74+t9A0r+R/4rs28iggZruF4Wbx5G8yXQWAQGAQGgUHg+REYweL5MZ8aB4FBYBAYBAaBlwKBNSvfzH1tyaMCsWI2KbIf8YGkR9gLx1C88xY1bWFQZAnCCrmFqJDPvmaQIj8cN1P3S1ZC2CsPSYCwEA89YowAcLsSMi0SB2mgLcqOCFF3ITyQEZEwWzKrWb6INPUULsr+bfiMvCKU0exjZIXfytafFjTVJoQGIgQuf3MlMz6/9ZAfKYIo81nYFeSZPAhAJImykCbIF2Gq5CPqwFq/kTE+kYRmQSNZiB7XkGcr22yDwCAwCHwKAs1sb7Y/24bgZd8Q7uzy7UpEaIRt4fSy5YRpHmvys9nGiBbaZs/ZWHb6lHfFnii/zyVib40hbGkh+thEtlM/2FKbsYJt9dl4pd68NvZhlfZtcFwytjTWsL+VS5i2/dpKRHxjW94nlWV/bWGzYQJfYyyMhVlUJmGn9ZuaLNA4k5fCNrxTIZaU7Rpqn/PK07n7Pvl9H/c7OG8Fi2PlXdq35ReIYcSkPDNdCxMB7uuF47q6X92PnlGaSEBQ+a1Dee5P90K4uk/V7Xra755xb2vD7UqFiSK+Kdu9ZPzNy2LWsbh0pef4IDAIDAKDwCDwAhEYweIFgjtFDwKDwCAwCAwCLzEC1IrWrsi7AYnQLFQv+17ovcQjpyQzWeVBUCF2HOc5kHeDfcpEniDckRWeNQrJgYi3IVsQObwuIuKde3M4v3AMeWTIj0RA8kgEhwgcYkdxs7WjGanqjSRB/BduYxsWynktYHq7vgtdoa3N/NQO3xMNCn9FfPH9G1dCUPU85XsChzAhvsMPyYYIsvmuDfoDR5gSOWAGc/kLraJvjmlDoacuhfA4VDMfg8AgMAi8BYFC5bFniNxmkbMtiNzblZDB7LS8yGF2mrDKTiGN2Z+859gqNpRNkw+JvA3pdK1XhUZu15rYXzb2VZ3seF5223dY32sDUSNR3fhkTQ523fhlq02OyUtMsDUOwYYdJtAIH5SXA6GBXWb3taX6O3/f5sZW7c1rwqfyeQPkEVH4J/kQ6nkrwqMQXpXd2KVu45nr03iQgPEQYSgPRGU+ZqHy7TogtVmZrgchAObqarzeY3buN+z/7ErEfefDSf89D3iOgAnMJGMmfF1318o5TUIwcSBxzj2fR6T/Q+uJJATdp32TdxAYBAaBQWAQGASeGIERLJ4Y0CluEBgEBoFBYBB42RE4hIMqZEOxpc0URQAgU+wTtggZgBBpgUsv8r4jfxAkQj0hSG5WQrb8xErWpEBSNNOUECGUknzKRb47dzuTMyIHGYTkRyRUlzYoD+ngfN+RC8h8fShsA8JMHRE29kutXeF7dasPWeWYlDeFvhZzXD2+q5PnSeUhQ4TGKowTIs93JIjzEV0tCqqNhSvRfvvF1tZPBAxskIAIQnXJI6Y2cgXOMNWOYpK37saIFguU2QaBQeBeCLC77B47YzY6jzeCc/ZQ+J7vWUkYJR5f7NMXrlQYosL7sLX2Kcsixghj5DBb55jvtvuQ59tQQac6dcpDwpiRyMxmstc2+/St9ti3Dcm0FRuyrcaWD67ETiPFC7EEp0JJ7UMSnWqvuuFkbP3nDuUR8Y2zxq5wzbOv8anxyLiSrTf+GJst/F2/GvsSaPbtMI4QxvNy1McmDcirr8Iyag/PmlPre5zq336/9iYo+V4Yx+2zQIuZ82iw/1osq0v/90KY/rmu4QNj/dJ/Y/DNSsZt/XUPC2lpnE5A6Znlp9Y+zzTua/+V2QaBQWAQGAQGgUHgbURgBIu3EfypehAYBAaBQWAQeJsQKDyIF/9mjHrhR1QJsYAY+sBKiQARUYXEQKg4T75CLchrdq6X/daHQLariyggH5IAQYGcMhvXOcpBHNh8R2gUq9sMV/uQB4kVeXDIb5/6im2uP8iLwjEhT9RViIhmkioDqRVp5FM+4Z6El7hZCZmi7YgOG2GB10TrXBBcfufQVuUi+PTvQyt9+0pCXukzTxMCDGKPR4XfCCJtR6YgBPOeaIat48gj4oV2ES9gFC4jWBwuynwMAoPAVQiwGYXpy5OMrf3NlRKmCdHysKm/sRJvM7YzO80WId/Zd/booyuxtfYTDcxef8ymXjbxvhu7q63sI0J7u7Gv2y0BOC8+ttcYw84j97VBiD92fhu26FQIo7wF9uIMsty4oj3KNAbAGVaNi+pm61snQjuc1/hsPMgTQx8a+/K8aD2mU+OBtgl3hJA3fhmjtluhroyzx8SK20Pmm915fv7codztIeMjYSZPlO0x2HoOUGdhoe4jaG3Lcj7xATYJHvB1XxNz8g7qmGtrvHZPt94H4QY2rk1ho9xDvGv8L2DaPXKk+7NrEBgEBoFBYBAYBF40AiNYvGiEp/xBYBAYBAaBQeAlQuDgXRHhgUBAVJghi3gyq/RmJURCcc2RJn4jzZENjjfjH9HRLMXCKfCy+LKVCmvkuPqIHggD5AlipnjSyBp1I8bUg8whhMhfHPVipedRgZiIWEPwKKMyERLqRNAUrgmhRbxo8fDWx0BM1D99MysTSeFTecpFavzkSi1OKz/yQ3nCZ8BQXcgOJAgMkTbaikTR9/cdjqvXTF3kDQEDYbVdIwPm8sLjdiXknXPkRQY5L8+OES0WGLMNAoPA1Qi0pgIbxyYSjdm4m5XYnoRmNgnJS8A1PhAi2Dn2DcHLBiLfeeGZmc+uFnLv6sYcydh6RteW0Uz7ROprCPA8MXoHhoUxAx7Gpvtu6jw2Gz+BwzG4w7S6EO28XPQX8W+xc2KRMSePR+VqY94XrXuh/fq9xftUiCXjm+tm7GjM3PaPKPOVKxVqat931/g/XOnfOQKKMGH7zf1g8epja2DA131UeMWHCFPVB6NtKEb74WzczWsFnnC2331uzDZGw68QjMZqzxpEOGO++9o1IgS1LsqRbs6uQWAQGAQGgUFgEHgOBEaweA6Up45BYBAYBAaBQeDlQqBZpkgqpISXdmR4BJCXd6QAwqNFV39mfffCf7N5mUc+RAggW8T5RsAIAeV8xABSBpFgtqNQSq1LgcThoWAB00JQIRiQHXlCFGsdkbZtJzIhQgfx05oWES9ICfm13eZ3wog8ET6EjcrSHnhIyKUW5lYPcoV3idmy+shTgmCh3cXGTmxpoexCYLWgOe+VcI9sEhbj5tAG5WgLcglJ2LVwbfTFMbgUd/7QtfkYBAaBQeAiAuweuyOxI+wXgv5rVmKb2Hq2DVnLpvMQ8114HTat2fxsZnav/c5VJrtpQw5vwzBdbNwhg7oSZK95R02gUK/xq5BN2/ryrjsmZiCoHd97Uzj/2HoMp/oRpo7v2533YAJ26zex68YaHiCR74kp1VMILNeuvjXGteZGbT0WUsv1EfrrmCCxDd8Eu0I5aV/jkzb/+ZV4IBiDtttWcCDM5yVC2D+1FWLrMWJFZW9xJkh4vqifhXV0n+qn5xZ9ck/qi7Fcn00e0Cb3j3M947iP+5/YNxMDzlzQOTQIDAKDwCAwCLxIBK55GHyR9U/Zg8AgMAgMAoPAIPBMCBy8KxA3XsIRE4gDpIbfXviLk43oR5A4RkBAALxnJbMqERPyifWMYHEeMl15kfq36zsCBWGA6FBO4Z6axYisNyNTG7RJGUixQpc4x9ZC3ogHxAhyQr2eYewr7jeSQRtaS6LFTCPSmpnqHEKK8vULKeFTn7QFgVFoEn1A3OkjskOZRItIPX2xKU+5tyvxCoETkeaHViruu99w9aktykKeyNtCoMQIdZvZrD3qtU9btQ2h6Dx4Fb/80IT5GAQGgUHgLALsIxtKGGDPhfBLmP3x9d0seHYFkcveINTZG2Hy2HH2jm1CALPtjrOXbKhyEywuiRX7NQhq9GPeSxsv9gAcEzHKw463RsVWoNa+U14HpwCGU8kYpDxjUmK6Y4nbrXnEjsOyBanh29jg3HDSlgQn45nrKCVwbNu6xfac18sWly1223OUz4vw0pZYcSwfYcA4ahKEsa81o7bCyKXyT4UK+4V1ovI9I8CXp6h7qPw+HdcPyfjLm8J5Nu35wEqw8F+AnfFaW2cNi0tXZY4PAoPAIDAIDAIvGIHHPBi+4KZN8YPAIDAIDAKDwCDwAhAw9iNpkE0IE2E+EEyEgBbc9gKPVGkxS8Q6IgOJlUBgVuhPr3RzKOvn1ycy/8+uhDzw4m92JxFDWcgCxAryAjFgwVfkRWtTIBaQCa0tkRDSwqXqJwxIiRPaqe2tRVH86WaxItmaWascooh+EhWch2zTNjOCi6vtXASMY8Uah1GCif6rV3uFi0L+1UbHvmglBIq+3hz6SJwh8NivrfqIvOKpYdNuZJ86iCcIE8ftKx64a9MisYgtx2cbBAaBQeAaBBKp2SpE7u1KbDIPNZ9sOZtGRGaf2CH2M0GiEHmF3HGOshK977N+RSEGWxPpmvY/R55m0x/zxtDXvAW1JWFd6EJjVR52jrWOgu/Gt9bGYLd9R47DdrteU2XmAeh3IRDzplCH8IO2Fhb3nUCSeHGq7c/9zm+MT1ixyLWwVzbjd6EOD7sufpzyyDA+/hcreaaAp3yeQRpn3aOw65nDOG9sd020yQQA46tnF+Or5w//jUSh8a64eGkmwyAwCAwCg8Ag8OIQeO6HlxfXkyl5EBgEBoFBYBAYBC4hgMyQCAVmFyLtfXrZ96IvPJOXfrGdvdSbTYsgsTAr8oE3QGEdnGeWLmLCd8SXF3xlNvuzRUSRAAQOpAoRINK+MEfNzkXgFDIKcYOURyL47vzCLCH25SsMRmGXEGDyFKpKPxM31te7thb+onO1IcFDe/VPvog9x1o0nJCgLS0savapuhAn+qj/2pWniJnKvjuWSKIf6hAeC9lFyMgDBQll/Y9fWQkmroNNuxKYtLcFuGcW6AGg+RgEBoHjCPzed7y5iDO7IyHOeU3crIRsJ0i/fyW20z4JmcsOfcVK7BN7yC7mAaYcNo3tO+XdcO6SPEVYoKe+5HCpXWxzNrd6WiPB74SBFnbeeibsvTPkRaIbCwpl6LP1nWDqfGOSc7fv51sBwjH15Z3gmijD2HvOy6G+PDVe58rrWcOYtl3vIo/Kh7bFRAhlW6MiTxZeKiYKeIYxVjaBwH0ZXiYNENVuDtfh0w84uvflIaR8ZKXtQufKH0/Gh16pOW8QGAQGgUFgEHgkAiNYPBLAOX0QGAQGgUFgEHjFEECMIE4K7SQMSDNp/9j6bv0ERBRCCmHu5R+Jjuhv0criXRMgkC15NJit6Nmi2Z7EDmUhehIOEiV4OkR+OYboR+o4biZkMdPtR9IjXQgYCI9COSET8oTQhsgKbVaWcp0jtSi4T20khGhn4oZ9zazULuSHzXH7kSQIj+1sV+XDJeGgcFJIFeJJYTxawFOfEmwQfdoCM+1wLsHI8a9e6fZQv74WqsU1q4zD4fkYBAaBQeAiAuwXe5SYzOazJezg161EXGV32exCzrFbv7MSkRWxy16x2/Zb90IInv26CxcbcsjQGHJt/sfkuxR+KJvegsytaZEw7nxjjdRi2ufaIz+swzFvAwR6IQjVaYxCiiPJ2fbCNcpv24d0ajzJy0U9xkVefue2PPMeg+Fjzt0KWvpNHMhDBMbnwnbt6yU0dL2Mx8Zp1wQOPCoKAVVILvi6x92zhfpSJ+9Gkyt4Wgjd6L/gP0HI87ywvX6P6fucOwgMAoPAIDAIDAIPRGAEiwcCN6cNAoPAIDAIDAKvIAIIEEQRYsYL/O3hRf196xOBQFyQEFdEBnkR5ggCYZF6bvDi34LcykIK5JmAKCjsknx+S8iEkhmNFudGHCh3OzOymZmIh9Z5iEDQ/gQEbSReaJO+2N+aEr43M9WxwmwUcqpZk/IRJyQCgva1wHfeFjwd1I+wa3HUFuZMqLg54CFkCBJKfm2FqVATeVc4biueeTHOI0fsV59ytV99yB2ChdnO6kncUMd4WBwAnY9BYBA4iwDbwu4hj9k4Nlj4J/aEaOoYW8qmsHVsXEK272w6ghf5LbG9iGI2tdBO8l37bnlufYWnvpT7un55VUBwacsjgs2PSIcP8ab1idhjWJ0TLCLSYanOwnD5NMaEDdvd90JtydPC4VsvAW1zrPHMmLWdFFBIxafCzLU3thuXj22n1h85Vb+yej7Iw7LFxJ1zH7Fif72M2X9ppf9sJYKFUFsEjZ4D3Muwks8zRuN4+/XFvc9TVBt5YTSRw/0+IaGe6q6acgaBQWAQGAQGgQcgcO1D5QOKnlMGgUFgEBgEBoFB4GVBYC24HeEROYOQIEoUSsILeyEUIq68sEe25LGQR4LyhLDw8p+oYU0HhA8iIA8FxA3C3qcykBZCTX3GIW9rRqgfWWLWpHYgb5p9idRIZCmmOnEBAVH4Jp+Fc3AewkE5yArftyJFzz/IntaxWF/vCCr9dVxZHdd2pFzkin40ixZ+jt+uJA785x/qRFAh+PTDDNhmgm5n3RajXBuQfZLynEeQgasNccjLRT1Ej65hZR2yzccgMAgMAm9F4NO+811vrLBQ2fK8B8wo501nDGBHW6iYDUfoI38dJ0yw84jg1s1hGy1czKYSU61PkHj8GPgj/O9Txn1Ekso19lzalAujrQeJ9kXAt07Cts1b4aPy8x5kw21strEDplvxo/G38xxr/NuGmMpLoHynCH/tMkbm3XCt0KDe2noMo2NrZJzD0tgmpCRxbItJXo+XrsOl48bLf2MlnhEt9q5OExV8wse9afwmSFivwnhsn3tef3gXuY9db/33HyFU9Z+51IY5PggMAoPAIDAIDAIvAIH7PnS8gCZMkYPAIDAIDAKDwCDwTAh4eY+E8TJvUWwzSQkItyshaRAcZtAiSeRFaOUp4HgiBcIBcYUE+OGVkCPOQ/oXm9sLf+GdlIH8QeAjRG5W0p5fP9RLVJDMlEQ2IAwQ+sUUj+DRbm0ibCCP5G/9CG3+4Er/zeGY9irnt1fSXn1tZnCzYJFH2tZCs/IXG1t56tOORIXW6khEsV9+nhTy6+/tSt+50k+u1OxefWpBbbOSlRlp07od2mLGZ2tgKMe10W7XKu8Yxx8yM3WdNtsgMAi8hggk2LI7wuEg7VtjiG1iU9gX9vELVmLLeXi11k/HC4+EHP7Mlb7pcM5TQLpf++GaMh8y+a4+7ctnj9l/Y9TWi6F82md8Y9ML27RvM5FByrsizxV19t7N3m/FivJUT2Ufs/Hbcs7ho13bUEzXvvMT+O+z1VbnnPJIMH5990p5PhivjY8/sJLvT7G5n8PUuA+77g3Xq/W6vnB9d4+7193T7n3XXX5l+G84L4+kp2jblDEIDAKDwCAwCAwCD0DgIQ95D6hmThkEBoFBYBAYBAaBtxkBL+0IDC/lyCjkOfLJPsQTov03VvIiT3xAVnlpb50F3gN+W2i6sCGOmblIgEB0KBNJ77t6CBCEAOch6dVbCAwECo8KJIZ8SB5EQvG5zWBtjYrWbii0U2Gh8thQJuIBmSPxctCuQmloj/6rR73NvNR3fYhI0dbCMyGuzDDWV9/ljZzJuwJOH1/pY4c8MEN2JcIoayt6aKOZnPIQXfTforaRUNpIoPC7GaOIFoIIbKXffzjuex4m6+tsg8AgMAicRKA1LFrTh03ZeqHlSVCopNbdUSC7F6ne2gCtHbRdi6KwfIVVeq7LcV/PDH0x014ooM7VdraXzd++H7Oz9dF5xqJTgof+JjLI25iUyGMsgLu6WmA7D5GtoHCNN8SpPl9z7lNdl8ZhfdbH/bokxH1iRUK7cbQJE1+/vrcm1VO0Z9tv16/nCLg2acAkh63HjO+eDbTDf8G16f/Rc8CEXXyKqzNlDAKDwCAwCAwCD0BgBIsHgDanDAKDwCAwCAwCLxsCK+TTuSY1C9SLO1GAwGAfwp8AIRETvPR7gUeKI9/l98Ivn99EB+EUEifUKc/vrlRoJ+Ug4pEZvAUQ80j9FrtGWCD6bdqhfEQRkguJg8CJjDGbVYgS4ocQVs1aRSIpBxmCaLDuA3IIIUEAaCFTQkTxwH0v/FPkm0/nq0PIpsgL4o269NX5rSsBB+0zK7R+WCgbiYX8+pmVProS/P7llfTfWh0/dajbIrXwh5XFbAsPsr7etU0YFsIIrxF9+yOHT+0kJqkTRvoXCVOMc2XMNggMAoPAWxBY4aASThG07Ad7zUax08RT321sINvK/rHZbClbxbb6lNencoSms9/YoXz2yP7nFiu0my1lH4WmajsnYmgv+7rNg6hubaJNMXd4eF9uLDwnVmzrbs0L5yVUwCfhaBvWb1uf79d4Q5zyRjn7ILCv6IG/P7zO+5KVjI3GJmNrXgraLgSkT/dRngzGwkIcqlY7hRl7zEYAganx2LXzrFHZ7lPjNvxb0LxwUIko2mn854FpTFWe/4ZrrFzPMDO+PuYKzbmDwCAwCAwCg8AjEBjB4hHgzamDwCAwCAwCg8ArgkCEUmsyIBeQ4WI3e6EvNjmxwUu/l/Vm1eYh8KVrn/BPiAGb8wgKSAjeAEgvJAVywD4EkvKQYDw4lBcJgCTYkh0RBAQBosjtoQzE/QdXQjAgz5SHEEPqIxMQIr+0kgWprfFgHyIN8UC8cDwvD2XrW/1FaCAsPrKS9lt4HKni2QhOhIWEDfUleCBgeFQUWkK96tA3s3PF6kaAaAcBREL+qRsuyvKJrCHC6E/kyvp6V4a2Igdt8vrtWslHINGGFlu17zlIqkNz5mMQGAReQQTYiEICsilsN28vdowYzd4VXo/tYsfYfvbQTHniMjvMtrJZLbQNCrZxO3OdTXrORbXZbW07t+mz/icY3Owys7F/8NDn7aE8SS4U/+bhiHs72HAis3GksH/wTJSX55jwcI1gcaw9rpvxRZ37bespcm1fTuUz4aC+Ea2Mn+4dzwjqdj8YA3k61hbPGzCAj3uxxcMf05bEse9Zhbjn/sJKhXPS37yEWtvCc4ixWN2FvnTf6o/JBj3PFHJxxtXHXJ05dxAYBAaBQWAQeCQCI1g8EsA5fRAYBAaBQWAQeAUQ2M7qNKs2coG4YHaql33PBAQBBLsX98JfIJ6K2U1Y+MWVkFVe6gsz9f71vZBFiC3lITESNfYxuxH1SBv5CAvap04kSISPtsnH6wARwwsjAg3hYCYkAkpbEBPEiWayFg6itSCUI0yTNmqT/AkyCDtES2tU+ETgKVu9hAblOQeph+Agwmi/vNpthqf26gv8zOz8rsN5ykb+JZQU1uoTa1+LfKpLn7TJPvUjfeCBIFQ+IQNBc7tSIakKW1GoqnVotkFgEBgETiLAziNwEbZsGaIeMWs/0t/+PC4qRP7Ebnl6f2R32GvlREKzV/tFmxHCRA+E8YvYjB+88FqkWh1bIaC1jNjrcx4gW6GA7c3jT1nbNSdOkf/q2ebTHra6MFq1CW4wMSa0uPde4Mn7A77yuk7K8T1PyC2Wjbk8Xo4JFvtwTY+5DrwJYaM9xsSblYxZef65/u4JY7QxseuRYGRsI9g/1TpM6tp6HcKya70VHdzH0vY+cbzQku59/XAPzzYIDAKDwCAwCAwCbzMCI1i8zRdgqh8EBoFBYBAYBJ4JgTwlzEY1k9QLPvEBAYKEKlxIoZwiWTQPQcOLABEQMeHF33NEIUN8b2ai8hEZyHvl/uZKiH/kAOIKidFM3RYp/aHDOTfrU9lIGaSDcwgE2k8cQC4QBBIflKVNPA9+dCXEFWKMEKNvBBptK+SHfiGVCBBEAMSLsrQXYeWYPPCpP9uY2NqjTvkKq0XosTWjUxv/4kqIP8eILYVTUScBRXuJOuqwL7LMZ7NP9ZNYQWDyXZssiAtPs6NPhQU5NGc+BoFBYBB4006w32wbwjnPim34PnaQrWGr89xKyGCHWhOIF5y8yP880cDMJmYLt7Czh5fEivuuQ7EtP7vN3iOdC4EVWe24cS/vwM41xuhnYa7arxzjAjus7fvtGPkvrGAhjlp0GzaNE/a1noLrkMB/Skgw3rb2kjYkhGwX0tau1jEyzqrvdqU8Cl6Up0uhEwuTpV7jWOJMExSaHNCYCn/YSsbAp9r+9Cro76/kXnb/dT8oP1FE22zaZHJDYaH+l/Xds0jPLPD90CGf/BMS6qmu0pQzCAwCg8AgMAjcE4ERLO4J2GQfBAaBQWAQGAReQQQKCWXc90KOLECmI3QQ/LwUEC5e5IkDERGR6M3+R/AgcpAsCHQzKRHxzZ4t1BNygGCAXEekIAeQFMpDXOXRob5IHZ4IyBekP9IMweRTGCptTLxA3hAMEksQ9z9xOE8/f+FwzhevTyQEUUC79bdwUsrV38QB7ddOZZoVKp/viLn6qx5rUfCW0GbHtQV28BFSQp+FltJfxIm+NFsTmYWwaWFw61k4powINqRgRBm8kC2IRZ4eYaIvQlmpv/jo6+tsg8AgMAgcRWC7sHTr5rC1BGCeYQRV9oiN9dvGtrBHCbmOsWc+EdZsVp5h9j00jFENfqj4qh9sOTvcGkPKRJKzlXnCsZf7917navt+pn8ixX3CWhmjtqLz/lz222Zcq6+t77DFTpv9hrsxQF7tzNNRGa4DLwXChGuoX8Yv3ojWl2irf4+9Npsi754ZJG2DrXvBb88B+pMwoB9wddzWBINErqdsk/KJcIR85au3+zOs4QVTm3s8oci973q7PvDS/p4L5J2wUAfQ5mMQGAQGgUFgEHhuBJ76YeG52z/1DQKDwCAwCAwCg8B5BCLDfTYT0ou9WM42+Lk10gAAIABJREFU5LpjXvQL7YGMIEgQIGwRKEh4eR1D4MtPPCBMKBuRkieBl395kF7yIQYQCZJjSH7kPELjZqXPWYmnhDLMekQUKPPzVlIvceRfOpyzPu7IKHkJGoQChFuiRKKGzw+shMzSBuQOkkVff99KZoWqg7BByNFPIoVyC7fUrFzt1OafXqnFvItHbqHtHziU3cKiRBD9gGWeJtpMfICJshBOyBN1RQARcRwv3Fazg9euu2vm2tXu7bV1fLZBYBAYBPYIJFjbz3axIZ9YiTjNbhKL27ZrUUTwOpYnQuGj2El29z6k/qUrk2B9KZ/jbHlrL7HfbLrxZCu2s8/27d93I9X19aFCiTZsyextHWGS96G8xrZCDTpeuCm2vvYU6k9+5WlfaxUZh1w7XgTGEOOHjTdMIbiMrQT1tkIwbXY9+qsxTPvDO6+bcM+7IhEoXAgC2pyXz6MbsgponSdlEYLgZe0szxrG4XB1fHsvb+9x977/gP+C/4T/BpxtMyHgKa7SlDEIDAKDwCAwCDwQgfGweCBwc9ogMAgMAoPAIPCKIIAwMN4jGBAbSH3kx28f9vUsgExBohR+wst6ZIT9XuL9Rkjw0LDPVtgJhDsCizhAqEAYqFtdyASiBrKDVwHCRRgkmzKFOiKCIOuVj4TZhpFopuZ2rQd1ISzeuxKxg/Cizp9bCakTKZEHR7NNC/NBaEH8a6P66/uXr++EhmZpKqvQULwk4KDt2m1/Asi/cuhDC3AXI16/ml2rHh4fPgkmW4Iq4cj59rsO8qnHtVCGa0a8cc2QMq5pa4FsyZm1e7ZBYBAYBO4QiJRnA29XYoMtiMxW28eWmJ1v1jk7cyysEztZYnPYJzZuu2bDY+G+T1nsZYIAG6lNhe9JSKjfrRnBphsX2HD9LnRSXg379htf9iGYtnkuiR3sdn3a5239h9a52HpQVEdjs2PGAv2V3/i4DSVljPrllf7ooW/GX3me4j2feN9Yr13ugTx2YC4lRNRHx1vfpLWu3FPbcu5zrxj3hFD8+t1J+3Bd+m9CgUkA58JhEdt6XjAJwPOM/4K+/NJKeVuo7tI1vk8/Ju8gMAgMAoPAIDAI3AOBp3iQuUd1k3UQGAQGgUFgEBgEnhkBL9zIDWQB0sDLPLIEqWBmIQIHSd7s1GatRgZE5iBvmllZXG5kBiIBOUJAQAQRI+Q1cxRxos7ioatHQhgQTgoNhYyRioGOiCc+FEZK+yN01KkOMauR/nlLOF+Z8jnPMw4ipbBOkVuECu1sXQx16rP6IpHM2FWOMiLp4IgYujnkK9QTHAlB8EP8KRfJlYBAMGk9DPvhqSxESSFBfKqrECaF0/BZKAvXCsbK168IIOd2zdbX2QaBQWAQeAsC7Ag7x/7w9iIgN3uc7WCj/OYVxlb5zcayfWy7DZnLlvqtnGMLOz8E9nPE8rny2FA2k/3TZm1NZC88USKGcrS9UH5stnHPWHLOy0If92LGdsHma/p7zAMlErwxbeupsV1rofJdl/BGphub9ZfAb8xJ5HZdEfEJ5Ne071KevciQKBSH0KQG4yeswkvfus+0tfOqL6HjGhHDuC7tt2NigmcC178xsvHW/dxYbex2zxhD3RP+A3khaXPntL7WJYzm+CAwCAwCg8AgMAi8AARGsHgBoE6Rg8AgMAgMAoPAS4ZAYRiESzCbkBeBdRC8mCN8WjjVi34LVHuJj7D3co+styG+inOe94G8iAchm5p5izQpfAQvA99bGLR1MhBfPYsgDJRbvUIz+I6oyMMBKSIfUueLDu3RN8RTs0/V8SMr8bTgCYHoJyioh1hhVm2eGsWs1id9QWhov+PKzetBVa33wRPFd/3VXmSM8xEwNyvVJ20qfrq82p1QBAuhrNShjdpGmNC/2lSscO1xfli6fuKUu5a1U/tmGwQGgUHgGAKFt2NHeYkRZNnBiHIiBvvDjrHNBF+2SN7C3vnMoyxCd0sYF6IpgePaK3GM0HeusSgPuHNl5YnHbmYzEfnGAWUXOqmxRz8Ks+ScztuGCao+tt1YYn2KPAJ/fn3/wZV41BlPtps2G+uQ5vfZtjj2Pe87n4lIhYlqTSn4fOZKRPs259fnU23Q5/t4syjHWLYdq7unHCscVKJE90feGIUTa1Hs1hd5LA/BE9K9aw0TGLhfu68Lzah9xkkeFJ9YSd9vVnKPuOdbQNy941yeR549jK+Ejb3QcgrT2T8IDAKDwCAwCAwCT4zAYx8Unrg5U9wgMAgMAoPAIDAIPCECkQqFZ/CC/7sreTn30u6FnSeEDbngBd2sQy/4CChEP0FDOQibPADysCiMQjNci5ld6A2iiBmgtytZjBqpgNQx21XZ6jTzMcEksgap0IxZZEhrXiCD1I1k0J7CmUTSfOzQF20Xy/tLVtJGIgISZxvOAomSoKAO5FNxwpEdrWnRLF0CDDKudUASC2CoXXlI6BsMfUbyOV4sbxgjtISvaDZqRJQ2IaHgCSd91W4zaJGINyu5dq6ha+m8uzLeeOONo8TKu999bBLqOmO2QWAQeF0QyJayR0RYAihS1sz9P3awM+xJpDQ7vSXBs21I/RZWZreVY0a6rc/HYpp3xO0qiJ1MHD9WbgKFYwkPDB5R2dZ7LrvqOLuq/dl5tpO93XuLsP+FvWLvEeIJFkR5x/dihfqMGcdCSBVCqT5svUr2xwqjaFzRF31ApBcCqvCMjZ/asg/btCXrj+FmXJFnG1bqWL7tvi1n0KCije6JRCD5uybywDfh3n5jceXcVzA51r5fXztdU/c0scJmXHbP3B5+V496CXVtrXHhOro3CFH+E/BVnvwJMfox2yAwCAwCg8AgMAg8MwIjWDwz4FPdIDAIDAKDwCDwjAggCSLmvXx7kTdz8BdWQoIgwRHiXuoRJWbzt/A2cr5wDcgHIgESZxu2SPmIrkJryKNM5D6iB3nwWysh6ZH2jhMTxIlGcCGK5Le+hdmXCR+to4E4kL/wTMQV5f2RTTuQDWZLan91fu2hLwgZ+XkltMaGtljzAvEED33Qf3mbuZqAoN8wIBjYp/0+iTCJQYg7i26bmUygkV/5ypNf+fYjvPS3/a0/EcHjmUz7EXYJOAka2qX9CCJhoVxD+MHjbg2LJUxsw4qsXbMNAoPAIPAmAuwEG+yTDUPUZs9kKkTeHjI2iG1hy9ks39kqNvWhmzKRw+zc3iODjUP6I5cv2bSIZP1JWPd9G15Pf40r2p43hzFOSsDerlXBVifq6B9B52c2HTXWnPIKOYXHXjUudFXXopBJna9fbL425i0hb9chgaLQR43N2kYUOBY+ad+2a8WKvaDSNdGnFrLe7vPdWFX4rcJqtQj3Q++ZY+cZA43j+7L1rTW5thhvy4BR7W5s958wGWD7X3nK9k5Zg8AgMAgMAoPAIHAPBEawuAdYk3UQGAQGgUFgEHgFEWjGJtIGAfJZKyFBEA6FIGqBacd7wd/O2EfYEwYiRpBNjiO5vPSbgWqGI5ICMYT0iWjxGwHUbEV5vuKQT9sIKtWPgEC4IGSUry2RSZWjHiQIIUO933+o98+sz+JPExTMHlaXMnhetA7Ge9f3ZqwmzkRcaYf8hYIiCBAzlLslZ/SFUONTu/7U4TtCEM4IN6QNcaR1K1oTBDbbcFPyqNczWfVvFzFtdnDhsBxDtvzKoa6uV7HP1+7ZBoFBYBD4FAT2AsCWSC/k3P6k7TjwFO5a2sDeGof2GxuWd8S5tQ2MReyr8SjxoLB8hTuqrXlU+M0G62ceDnmoZae1h9huDGpTPk+9NmODeh+71T52vb7CRvuMIba8FLRJvfrik3eFbe/RsW33f7mOf/uukZVzn7Ybfwkhf+DQnmP3Q+s/JeLDOaGjdTr2de6FkHNtOtYX+YldiRV7r5Vt+afu2+09v89zSSy7D4aTdxAYBAaBQWAQGAQegEDhCR5w6pwyCAwCg8AgMAgMAi85Ar2EIw2Q82bFmv1/s5LY13/40H6ChLyREXkVICvsi0CX3fdPrITkcR7RwixURJHZsYU1Iiog+r9wJd4FP7FSIgKSH9GAZCIESNpihqN92oq0KYyE/FvPBG1AkihX/X9yJf3RbqSMvPop7BJi7JdXMnNSfqSOtmkr0QPxtfUaufNYOOzbLubqmUle5ziufmUhcvSTt4a2O0a4sIbGD6xEfPlDKylXn+GkfVLrfRBGeJgo377ixq+vdxjbeJXo481K+uZaFqf9XUJCreTzLelw7nwMAoPA641A4aDyPiDqsuF5KRBS2fX9xv63FgTbVXjBX30gnOdEj2s9F9jZRPBtM9heY1YkeeOZTzZW2yUEfAtTs+vKamNn82TbhwIy7sDgXJiqa2DJa0U7G3u24a1cozxAfBpnjG3yhFFts884VV+J+MTsvVihXX/3msbt8hibbw7ld2h/DRMNth4Ll8StS8fDRZ1/biX36n7T739vpa55x42ZnjVcc1geq8u97p63qUv5/hO+b/8rD4BsThkEBoFBYBAYBAaBp0BgPCyeAsUpYxAYBAaBQWAQeHkR8LKeOGD2KjKGx8EPrYTMt6DozUqFmcgTooUynY/gt7+1LYgEQnYg2D1LmPGPxIkMiyBC7vNmsB/ZrkzntAZG+e0zW7Q1NZBI6kTSbMl7hJGQSMSArz+USehAXDimfwgldfokAgh/pXxrWigXUSEfYaA41upuYWyERZgpp8kdeWEIAeW4PihXEnZKe+1DhGmTT2RT/W9Bc6KJugkW6io01G+v74g0cdvlzbMCJsQWdSCjiCPO1wdYuCaXYpavLLMNAoPAa4pA5C/RlF1iQywuzI6zZ2wR+5XHHZuD8DU+sL9sERvbuj1soVA899nYNrbwRW7sb2IC8tyYFvnfeKYP7Od23Yr9GhaNd/uJfcaO1rLY96NQUcomGHzeSsdm7TcxoE91tWZThH8ho6o/YUO58rh2NkK88TvvPeUYZ09tx0SMx1yPQhYqQ7vylry2TONcAoE+bsNU6Xv9d82Ms9t1VdTxIys5tvfGae0n97PngjwXeYY2YaH1WKw1JZ//Auw8W/iP+K8UAvPa/ky+QWAQGAQGgUFgEHhCBMbD4gnBnKIGgUFgEBgEBoGXEIFmxHpx78XeS7sX9e89vKxbJDriBClupmFkvlmKXvibRYnIctz5/+tKxdounJT8jv+PK/30SsgvRARCQCgLhFLxpSNtWosB8YLUKuyF0BvyJGQgzewrPnZhrsqPnJIQN+q/XQnB9FdWIqo4hvjQ1sIwbWe2Ik2Uj/CIgBH6qX5+fH23/oYZnMrVT6QG7PRNUoZ2+eRd0uxdszkJDMpzPoILloXOag0NvxErMFGua+NauFYwL+yHa9mM3/1M4HVotkFgEBgE7hDIxrF9tyshZdmfCPXEVXbGcbaIiMvebNdOyENBmcjm+2wvWqzQlvqTB0NhgtjibLp8iO/E8lN9OLbGA0J7u984Ax+b/hnbjCs8Do/N6s9OO5aA4lzv42y5VHmtPeW4fc4hEumHctTDg9AY4fq5Vk+xkPUWD2PQuS1PRO2Hsfur9p87z3hu7CSW6Useh8fOKU9hsLZ5CDDCdRlTf3ZzQLsSJOCmTfBposDt+u5elydPG/n8J/w3HNeX7bPBBSjm8CAwCAwCg8AgMAg8NQLjYfHUiE55g8AgMAgMAoPAy4fAlihB3H/6SgiAv7FSngJe3r2kI0IQEF7okVKREAgZ5IhzeQFEsHupR9wgIORH0EcMECbky9uhmaLyIeXlQ7qUP2+K8iFMkDgtpIpo0peblX5+JSSDEB7OiyxyHMlP1CA06A+xoLUkEP7Ft9Zn/ZcngaLQVmHAS0T4JaQH7AgVzYAVDkpdztVWuJjx6lxeFj6FmkC6wM5vxMlPrqQd+iNph/MRObbW4mjB2BZFt06HOgknwk7ZRqw4ADEfg8AgcBSB1gpiy20R5uwW28I+IXmtCcCuEEP3ngTZR+eykfKx25dC+5y6JHnaJYQ/1aUr5B4bnddcxDOPC9/VzYbqY6H8TtUvf+H89nnUtffO2OYhXBvnCA2R+o4XWqtxxzF5jQGFCtR+16Sxzzmw1t6EIx4ftyu9/xHX4RzulwSQvPsScXxewy0Y70xgODZx0vio78ZAm/F1G5Jyu0C6fF+5kuujXufKX/naX3vU1wZDSbnK8x2+8Dbeu7fdI+Hvc7ZBYBAYBAaBQWAQeGYErnmoeOYmTXWDwCAwCAwCg8Ag8MQIRCptF6Lsu89mpHppR0J5gfeS7jzPCnlAyEe4QK7kIYC08OJPHGhxaseRCHkcFGYJQcGrAFEkRFMxueXldZCoUIgnhAThRJIXua991nDgrRCxpp1Eida/cJ4yERfaQEzRB9/1S5+QV3laFO6kEFTr0F3f1eWcFnTtuDJ+fSVhnJxrv89CYiBBnKMdreUB2+KoK5f4EdnlPPn1U7tsebhsZ3kWMkTbtt8Pp8zHIDAIDAKfgkC2go25WSnRlVAhtN82rFCLXu8LibRnw7ONDxUrlM0GsvkE3WOz55HGROdr17WovYUbbOwyNul/ggCbb+MFce49uPFROXtRRZmwg4Vje2+MCHTlEyysYbQl5+3Ps67xt7FC+8LVGJCnXWNFXhjqhc8Xb/Lvr9ljfx/zMtmXqd0tdN46G5fui3MRHggOeT10DfIqUfcxgci1dQ8l+Cfi5/25b3P3uHLd+9or7KK+fO5Kni1+Y6XW0XosjnP+IDAIDAKDwCAwCDwAgREsHgDanDIIDAKDwCAwCLxiCGwFC7MyzUT80EqFi0KSSIQKRBGiJKKGiIAcQcITBQqvAYLCTBESEjkQLAgJ5AFSv1ALzo8Yk1/opcSI4qRvZ8cWR7xQE8rTNiSD79qLNGqdCTMjtVMoKG0gnvCMUI5QHrwaai+ix3nKs0/925m0iJdmJReOIxEF0RZBY+as8rVH/xFw2iEhqpBJ2tGM3sKAILDsV2beJWaACm2hTfrVQqvF33atvmel9x3qG8FiATHbIDAIXEQg7wgZ2Ssixc3B3rBd7NM3HEopzJ6fxITWDWCH8sxwbLtQ9cUGnMhgDMiObbOwn+zpKWJ7K7zvi05Qsd/31grS9jz+9kR89nxb1inS3djCzrPPxiZj6V7kaTxR/1estBU8tmsjqEPK+yKPBdcoXOxr3NDuPCzUcUzoMXGAp8xzbds1ptTpftKfwk8m3tynPVvPjsJ6dS/4/LGVeFbYhIKCkTHeelWuS2ETt2LX9l7e3uMfWfmNwcbdm8OnyRg2dR+7P+/Tl8k7CAwCg8AgMAgMAg9EYASLBwI3pw0Cg8AgMAgMAq8IAl7wC3vkRd1mMWov9e9dybNABDlxwss7AqAYzgiVZjh6qU9sQLB7mS+cReQLUQMBZK2Hjx7qu1mfSB3HCA3q5yWhPHUhXpA0LcDptIgKBA3yA/GhTcgE5SPMkEcWo/6slYgfyhMyCeGlzIgpYgnx4tNXIgo4zyzjPDryWJAvcq9wJ4WkKgxKJBjBI1yt+xF5pd2EGXVoD8ybRaw+glHkSYSK+uV1jnOV3axgs01h9G0rqQd2sMorRBsKZ7G+zjYIDAKDwFsQiHxnR9jYRGeiKTvDNtqyoQhvdqzZ7PKwMb03+v1U75DHhAFeZuy+9hyb5X9uBv8xjwz59eVUiKNzoY/0lVcgPIwZ2sM+13/tPLUZKwptlPC9XasiYcP4pt2Npa0DYf9+QWn1bceAPDO0wfhhLDeOIfBtDxEMnJdIcszDZN9f7XbNtNU9tsXzIfdJ11zd2+vZM4EwkG0mH3RdTAQw9jtHO/YTIDrfWOv5QT3ufeOx6wSrwlEmMm29Gff9nt+DwCAwCAwCg8Ag8AIReMhDxAtszhQ9CAwCg8AgMAgMAk+MAMIlkoRgYHat9RW85CNeCj1ESGgR0WZyNrsTGeHF3Ut9+7aeFjwpxAQnYhAVzDpVFjLAeT79JhYgwxAqnkG0oRjdfhfbO4IMFEiEBBPtQDxpA3JGWQgLM3V5O3z/SkgTfSRsCC+hL8SL1ooobJV6wwb5T0zI0yQBwPFCO6nHb54TSD990R4iiPARQklYwwKZ5BwiinU2CBDaYZPfDFhiCMFIu/LkcC2+YCXt7ZrI5xx9E8JEn4SrEIrKtey6zizQA8DzMQgMAp+CQB4JCFs2w6x0Npi9sWhx9ikyXgHse2RxomnvjWzyNeGCrr0UbDlRgM1UNpvIxtp3c20hZ/Ilut+nKPXXln9hc+Je3Nj+hu2W6HZa9r2FsiP3KzJxwtjjWOtGNSFAvkTzhBrXS17nFAZJPmPU5+06+ZB3feNf4pax6NI6I9rgHoHTpXUvTl0Dzw3GO9upNnc/dr/KmzDjuzEcBnAp5JYx02SJbR+Mtf3WZt9/aqWPrWQsd27rVszYeuqKzf5BYBAYBAaBQeAFI/CQh5gX3KQpfhAYBAaBQWAQGASeCIFetr18I76R7L98eBlHRHiZv1nJbEMESCRFZH+kfus+FF/bjMRihSMakCyFgkDEIxSIEcQBAoLjSClCBoIGGaOsYnlXTzNqtaPZp+pqlifCAjGCLLs99EPYpcgJZMWvHsq37++tZFFvMyqRFNs1KvLYgAnBwuzMQp6oXz3agETxHYlDJPg7Kwk7RTj5UyvJS6wgypj9Ki8vCiKKcwkM6kZYETMcJ56oH85EF/Xok/7Z16LbzpEXdurUD+39tcOna3pHrLz73e8eYgUQsw0Cg8A5BNgds/DZYHaP/Ubo2s/OSOxcnl7KamHiiNxzC00/BH12O08xY4H2sIV5fjykzMeek2fivpzs7H4hbnZYqCj90J82NprNb3KAMYAd17etuJGHonFRaCN233gY2Z6AshUEnF/ILvWdC5V1DI+8PvZeKU0SKBzhOSyrs/Wqtnn1u9Bhp9qWyOOeeog3yDYEFmzcqwk/MINhm7GVR6ZnFNdIgrv/gP+Cc/037rtuyjl85tggMAgMAoPAIDAIPBCBESweCNycNggMAoPAIDAIvCIIFGapBaYR6GZhIhDaFxliH4KhsCGFZPBiT5AolFFeB0h2IgRiHjHgPPu8+NuQEGY9Iu99v10J2c4DAqkQUaCeQmskjjQjtVjmhWpC2BND3rNS61Zoj2caYaYSAMycJF5os3RzaBvhwW9tRpYgfJplqU4EE6KGuIFwaUFwuCGkCBvwE5YC8aG9H1oJCaVNEUr6pu/2I0l4tei39ikHXupQH4IEBvoAa/WHofL9dq3y+NCW9jlnS8qsn7MNAoPAIPAWBNgX9o4dZ4+JomwREpctRNgSMVo7iHfYB1YqNFThdfxmd1u34b4k+anLknjN3rYw9qWZ/U9xie/T/jwAGzerXxmEHkI1L5E2Y0DrGRlj2Hbjnutwu5JxrLHUOco3NhA3jKPGh8bivYBif2ED80w4FyrrGFaneICtILUPSXWsnFPXybNE60Ukdu3LS/hJsFF+oZv2dW33Gx+Nr9v1OrTD/Qxn+Mivvtapck8bhwsXyYMH3k0c8J+Au33OuS+ex7CZfYPAIDAIDAKDwCDwQARGsHggcHPaIDAIDAKDwCDwCiCQ4GC8j2j6qvUd4Y6ML7ySY/Ii8pHniABEixd/3+3bxi1HeCEEItkRM0Iz/P7DfiKGEFGR9wh2oZN+5YBZpHyeBUJK2exXF7JAmcpHIERiIYqQ/gkjCBEEXHGzlacusy710QLVyHyzWbU5Dw35EBnEioiNFj5NPIBJRF6hUj577YOZMosXrg3qF6ZJ2CZEChwQNdqGBCm+NzwKCeJ8/UJS6WdklTa5Do63xoby1SvpC7x+9FCWvvxTb7zxRgTW+vlPtuV58Zbf82MQGAReLwQ+7Tvf9cbvfceb5DZbxI6xM4jbwvi0UHFx/dm17PtWxDYOFPIvL7v7ALoNm+S8hGj2s0W4tUHd2c37lH/fvNcayMTiffkJHoR1ofvY8TZjSOsztUYFe81W89Qjvn/+Suy8cvJ4MDbVri1JL89WwDDGPDQE031xOpX/UritxCftPOYFuG1/ng2nPBy2+2G23bpX3NfG2O3YGd/xZWv/VozpnjcJwbVwrrCOP7MSbLV3PBef6k6ZcgaBQWAQGAQGgXsiMILFPQGb7IPAIDAIDAKDwCuEQARHszOR517IkQwEBSIDkog4gBjxkl9opy1pgkhBNCEXCsmEzE8EsRg0sh6xbnZi3gD/7fr+LSsJs5AngbqUhXjxieBBHCCpKlPehAh1yJNoou3IhIghn9pFRFDPH1gJwWb2KtI/T4T19W5D+Cuz8Fa+56GQcKDuhJtmaMJQO+VB2P3PK+mLGbVfsdLfXolYkWcEIlB7YOc8GKnHjFAeF/a3cHZxzrW19TMShexzXfTFNesaKp+odBfvfUJCLRRmGwQGgVMIJGiylRL7x8awZ2w2shaZ+0sreT+UR1goWyKuMmzs60OJ3P1s/Ow4wr/xhejMjueF9tRXldfbucWy9/UlKh/zJNgKHnnMKZ/43jofrU/Re7d+fvnheEJ516UwRepybFt+ExBqX2LAU+PzIsprUkReIQk3xvrCRj2m3jw3jI/GVdvWe8VvExlcS2OvMI7yufed678Az65Dz06PadOcOwgMAoPAIDAIDAKPQMCD0GyDwCAwCAwCg8Ag8M5GoMVWkevCfiDbkU+eA5BCiRQEg8JQtAZDM0i96MsfuYBoQMiLyW2GInLGd/mUkWcEUcIsUl4HFngVZiTRAUEgb0JFC122doO6lNOsSech1bSt2b2OIYiEdfCJXEtkKMRT5JrP1upAWqhPntbhaF0P60XwcoBLs1gjqwgH+k7sERaqOOIEEnXri7J9Eiecj5zRPuSI3+ox8/ZmJcKDdumTtT9qf6JPYbNaiNa1cw1dy+3ioOvnbIPAIDAIHEUg8pttskYC0TQRmr1k6/Ic+8j6bsa5kDlsnc0xic3Mjj4F1Ox7XgTZZvVrz3Z9hqeoqzI+vCtMH9nVU5sx7RqBprBZytEn5Rpf4JvnYAuWE2SE1XKc8xxrAAAgAElEQVQN5GuBb2OcficSnet3ov82j2tENK+9CehPid+xstRrMsOpzb2kTfIZWxvrPTMk3tdm4+R92r0NiQg39xRsEi7g+7uH5N4yhvfc49p4lnAd/Cf8N/J0GZ7kRd81U/4gMAgMAoPAIHAGgfGwmNtjEBgEBoFBYBB4ZyMQSeClnWcAUt8LuU+zab90JeR6MzkR5RH5EVNe5pEMtuJD24ccMAuXsKD8H1+JN4EkPEahLrz4I2HMapUvjwnPIYVnQi5I2rLdr12t45B4QiRAOiAafEdCIH/UiTRRRwRdi2fL1yzjQk3pjzLVWYgr+4gJNn10TD8L36T/LQhOsGmG5nsPdSonjw9tKCSIUFbNuEWSEHBgUtiJiEDtlNTtfAINXFwr16wwLa6lfiJeriHTDl06/vGzv6Mbd5s6a2eE2Cff8y/SU2YbBAaBVw2BFQ6q9QG2Yf8IAjwZ2BHiJ7vGprJ3X7cSgZVX2M1KhQg0ez1b2Az51mR46HoTkc3WGyICs5eJ2teGa7rvJfmm3Qns8bkFvvfhh/b1bUP+tWA1nIx3eRY4p3HD+ECIzruiscdvbYFlY922LmXbH9Z55m3zsN3Zb/svtb01Ju6L4T7/vt798TwgtB82+qwfcE+M73pfM9i4d+G79WRxL7mfnQ93Yohnk7wT3Vvd2/Y5lzDyiysVwrE1rrb/mUePr48Fd84fBAaBQWAQGAReRwRGsHgdr/r0eRAYBAaBQeB1QgAxgOggOHiBFyscUZDQkBiAfPdcgEDw8p4HBsIDec5bIE+NvCkQL477RB588eFcxIAXfwS78hAUH1qJF8Knr8RDwDHlIhmcixRQfuFI/NbuNuUV/9x+JFGxzoVGEpcdOYFwK5yG44gwdRE0kCaIOG2OTGqGpfLUaSZm61IgLWqH78rVRrOP9TGvCR4mrU9RO1sPRL3K4ElBFUCowFY+pKFNuXmnwF77hK9A5DhPndpE5GhmtPzqgEWhWg7F3e9jiRWRa/AiWBVqpFmz8J1tEBgEXl0E2C/2hJ1jDwm51hSy3yLP7DRbwhawWQh1do4NIKyyP9m4CGefCN9r1lFQ9v69kw3k2cAWWzeArfO90HradE3Zl66KxZaFLNxvkdaXzr90fLuQdBhFvhfKsDUc4NAM/7xLWqOpPI29+3qPvbc/VCiq7KcMK+Ve2Yol2/bDwZgVVoVDLP92rO+8Y6JNx0yKcI/aPLv82ko8Ht1Peajk6el+L7yYe7tJG/4PxrafXUld/hOObSc8XLr2c3wQGAQGgUFgEBgEXhACI1i8IGCn2EFgEBgEBoFB4CVBoBn8PhElSPIvWOlm85JOjPCSHqm1neHYzP/ORzAgSRAMyHfPEggC+xDqnziUFQnjfCRUYaEICsiD/20lpD8C3gxf+c10/KqV5CnWdAttJhZovzrNjmw26zcc6idoNKO0mbvWlyikVOIMUgKJhfTQNsQ/kkiZknOV88uHPGYWF8ccTtrOY8LC3kQL5RIYIvL8JszIK7wUAo6nRKKQsp1nc44+JbQkEDknwSTBQJn2fWwl13J7bQ/FXfexRIptDHtCkmsgbMftSnnPFCLmukIn1yAwCLysCORdVmgi5DG7c7PSb6zEpiFw/Za3NXz8zquiMHqtQZRgfU2fT5Ht7KIxhYj9wZW+daVCBD2FWKFtx8QK+9n67UbAIXzbjBHq3y7SnDB8LlTQvp/OiSxnr401bLs+56Xym+u7sSTR3rhDRGKXX6XtlFjhOcF45znDvZQwY5zsntpfC/02fhbiaY9Da030fOHZw/3s3uzZw7hNtDDWmYhg7HQ94G78990kAqEYb1fyn2jse/REgFfpwk1bB4FBYBAYBAaBlxGBESxexqsybRoEBoFBYBAYBJ4WgYgQL+HIErMQkS7I8WI7e7H34m5DPHSOzy1Rg3Q327bQUL++viMLEAde/hETZsYqD9FeWAb7EAeIfeIDMgahQBzRFgQ88aAQFXlbOFZYq+Jey0uEQFp4lkH2qxcZRITQz+9fSX+EF3G+2ZjqbW2OwnE4Xz6kkn1iiyPv/I7wyOtj7borQx191yaEjA0OykD8I08kxJc6CR4wc672wg0Zox/a27oXiRTOgfVHV9Iv16pr5zOi5+pwFUuk0HYYuxbCr6hf3wqRpb15bfge3nedm20QGARePQQ+7Tvf9cYKCxVx7tMscx52bKJZ5ezWDxzsC8L+y1div31nj9kExH0hibbhfR4atklZeW+wQ2wjIZad/H0Hu5SIbp92aPdTb0ILJQwkVqhjvyi3NgiRZbwkgl8KtaSMPAQSifw2RhpfjYPGF2Miz4CEefXCt/UX9l4GxzxVrsHklNfGNec+No9xx7Uz1ngm0KfCRcKi8I37ehKLzrXdse9byThbiCxluqfz4DQx4nNWMk4LrfiTKxGntOHrVyJe+C/4T7gfjLuJclePr48Fac4fBAaBQWAQGAQGgbciMILF3BGDwCAwCAwCg8DrgUCkP8IAAWVG/R89vKC3LgPyhAiArEYWIRoQUl7sW9sgLwKkO8KltR2Q2xasVD5PAMRM62TwokCSI6KIDe9ZKaI+9JETZsJqZ4vBFiYCeYNQUGdCS6E2mlFpRmrxsZX9LYf6C5mB2EDOEVuUkdeE+vWxWZnKMBM0HJodm3Di2Ulb9bdQTZUR6aQsopDfBBDnwhy+eWpoh6SsQi85x0xjpJW8hJQ8P5BqQlcg9dR7cu2KzXoU2qVuGMAe7s7VFmUTeSTtFP7FTF9iyKNCTKl0tkFgEHipEGDjEijZ+5uVEOVsNfGS3Uais13sZJ5nhdFje9mkbHOEbjbvvp1lR5H/7J0yvuTQJvvZKKQy0ZngzSOQ8PwiBAshEonIl7w5HLdGkrwtwr0Xa2BnX4tth7fPZvfrA5tsjDXWwLW1kBKwC2Wknn27Hvrufs4r5L7X7r75jXFwNq4ad+GjX+Hn0zXvXtqLNPu2J2AYrzxnGO89y9yu5JlDXZ4HjHvGN3V5hiBkmEzgOrn3tcczh2vw8ZWElTK++i+oI6+k9XW2QWAQGAQGgUFgEHhuBB760PPc7Zz6BoFBYBAYBAaBQeDhCPTijQgw29ALPtLayz1iComCRECYIxcQU828V6vvrc0gP7IFyVLMcR4JyPfWpkAOIAV4CXzhoXykgfw27UEqIMgigJAJCQURGUQKRAYSXVsRbcgLZJk2yIewUB9hQF75lIX0Qerrp/46l/ASGa89iAkeDEi7PDa0u1mfzo+kQ5yZgakO53zloW5kh0RMUAdSSx6kH5Egr4U8TlqcNIKm9Tb0xfdIFgKCWaIRWvqlLzeHz9v1ufV+eddOqED+ECX0zea6E43gBXfhtwrVAWcYfsps0lls+4DefAwCrz4CbEL2m71iS9kon+9biYCQJwX7yKOAXWVD2E5jRGHtEhbYLTbulMdB6w4dQ499Y2ONLY0xZrgTuH90pS9diQ3j0bANzfSUV4IQfEms0Af2Wj5E+H7bhuaDhzHDOJOAYd9W8NZXYyXc7DduCAPlNyI9Yf6YYPGUfX/RZSUsJP7nqWgMTMSpDU1AgNUlr50PrzzG2ZtDOZUBU4JEExPc68Z196znDWtNtfA2rLv3XV8ej/4T9juP0GH/bIPAIDAIDAKDwCDwNiEwgsXbBPxUOwgMAoPAIDAIPCMChXdCgCCIEAhmFCIJeFogEBIhkC3EB+JCsaa9uLcQd94IyG5kC1JCuQh9AgVi6cdXQoL/4ZUIEq03gYRHBjiPOEIwQKIjpSLswaJdknYgfQgqzUzN66IZqvIh87U3IkSbtB3J1CKcyrVFIuWp8WVrnz5HmDieKKIP+uR5ySccHYMFYk3sdzN/iRH6qh2FflLmNmyT7z+10hetBBPtb9Ypsk/bCTPEBPXCBqFnv9/qcs30K5JP/+5Eho1YAUek2tcc2gQ3fcuTQl94uSB2/tESJCbkBQBnGwTe2Qg0BrAZibk/d7AfREw2hm1uIWpr77BF7EXrC7BZ2TR2zpb33Sn0Ti0KXeg/dolQwtYbZxD2n7uStSw69ymJY+OBMaftmACx7wv7aTY/wfqYuNHsfVjlHeC79sMp0dzYkScf3LLFvvMw8VtegoWtz1PYvuz79dd9ZUwy5nlmMJ4l8u/bf0moKL/7kafGfnNfN6mhyQrGVNfOs4fngsQI18F4qi0mIAgL5RzXwPV8c2x92UGe9g0Cg8AgMAgMAu9UBEaweKde2enXIDAIDAKDwGuFwLvfffZd/421wcNLOEKKuOBFHZnwqyshFhDkLYzpuBNuDse89CONkPBm2XrZR/QUlghJgMxCCPCScNxMRuKFl3/fETcIMOep2wxJ5FEz+xEZeT/I67dOJRIU87z8PpVvBmXhSQrXlOeBY8ppLQaCgroLaxX5pN7CLCkz4sn5MOr3+npHQol7rYy8POzXL4TJJ1YiEtyspB95fcAQMUUogJfzfVeH8rVBGBSYwsu1QBoq1zWyX33a4xrWp63goO1wNTOZZwtBJC8VhAzixr4RKhYIsw0CrxkCeUMgbdlpIoF9tysRU4WGyjOLnTQDnS1iX9luoil75FznsS1s2UO8H9gjtopNbA0HdWf3t5cmD4xrCe1zl5Xt3G7XiALGR23cb3kQJNxrPzttnCHCs+uNTXk5bvvQmOdYHirGg0SPp+jvdpxQXmPfc4WIMm7frkTQt/ltDK2P8JHy7EnQOXYNjfnGbAuU7zdiiGcTmPOUcG8SSXjQuBawNsmASOH5Bi48iAhFcOFJxDODeLYd14+1Y/YNAoPAIDAIDAKDwDMgMILFM4A8VQwCg8AgMAgMAi8BAoVWEm7Di/3nr4S8aAYiAgNhhYxCICDTEVsR7ogqxEphiRAryJ9m+3vJRxrcrOTl3zHkuPLNhkQatGYDQge5rzykPDKhRU4jVbQHsaH8Yl5rC9JCu4kneUL4VJ99wj8IUYXUSIhZX98SDko5ZhXL7zxkke+24mjn7YCwi5SL5EG26Kt+NvvYuUSGj6wknjbiBRkGJ+f5RI4gRSThKwgbvtsQMfrLU0Rem37ASlu0D07EC9fGvsgoeeGGnEH8WFiUR4hZpa6bmdTa9X+NR8UB2fkYBF4vBNiHRFl2Ku+uP7i+s8OOI2vZJLZDGKjWKWIT2X157Ov9sXB2D0GSqLrdmtHO1kvsfiEErxEVrm3DMeHh2nP37U1QMB6wx+y2ca0QUPLnZRFJv/UW0Wf2ertmEBv/lFtt3K418qLECsLSf73SN6+UBwQ8jO3GMc8WtoR8bXKtjcXuKYKC8aqxWF7YekbgFbMdax1zH1vn5E+uZByX13MI8c2YLr/6m6Sg3NtDPZ4TYCOP6yZEov+EMt17rk0TJtQ12yAwCAwCg8AgMAg8MwIjWDwz4FPdIDAIDAKDwCDwNiLQ2g9Ify/lyG9kgoUnESWIBMQLb4u8ExAN8vuNXPdCj8yKdEB+iP+MGEBIILycjzAo7rkXf6RMs/3VjUyPFPBbHcpCKiB3CkOFzED+I/TV4dlFfmUiKZAeSB9lO4cogrjISyNhQ5mIC+dG3ihLvyLs1tc7wkM9ykOe1Idm0cqrLHmQMs2ild8+ogQ8zEgmCjlOrNE2bUbC5emAGORVQWgQX9v5hBDnSHDWXjObXQfthpM23hFfPGtWOKiIRPkdQ8LcrmQ2KYHqf19CxSykDbDZBoHXFwH2g20glrKr37cSG2xRa/uRwrzH2FrjApvxCyvdrMQesU+F1GvdhuziKRI8L4RrUFcmW37JY0M+45C2m0V/aisU06W68367lI9HoPFE+xDezoMbm16b9oR74Rbhzd5vvSZ6D4ddHgeX2nDNcdeostX3FJ4axATj1LnNffOVK23XM7GPsO9atOXZ2DjdxAfPDQS07abtp0QmWCuXQPHZK7kenlFcE8kY6TlD2794JeO1thlrf2Al1xNOFtr+eytpl/+Gdrle2wkBu2bNz0FgEBgEBoFBYBB40QiMYPGiEZ7yB4FBYBAYBAaBlwCBRWx/8hAWqhBCXtZvV7Kmgg0RgxRP1EBO2JeXgGcGhBdyxou8c5H0hS/iVYCQyWMBqY8ckMeGjGhtiTwkkArCjvjULvuRBggXs32dozxlIYkQ/+pA6iMqtKXZmPJ0fgSSNiPe7E9gKXRVHh7Fq5ZHv3o2QjQhkvxGmiBCClliH2FEWbY8UvTXuhOIFLM1tVk96viZlWDqXJ4T2sMLhFhUyBNYR6LASl8JFkJY/PRKN4f67q6ha3r4DbMPrPRvrQSzD6+ExFEWnGadigNQ8zEIvMYIFF6PrWS/2B02rlnw7Atbxr62HpExgbDNlrEzEntmy1aeEyWunc3PtiYkR94rly3Thj9xqNNse+GFjDuXtjzVLuU7tWD4/jyCTmEQEdtEC+NbAkEiznZmvu/GEpgaX1rbqLyR94U7aqy6tBD4vm3Od13VtxUsXM+tQPBQ8cLYpaxTa5LUHuWrzzi0XWfi2LVoIoN8ziG4X7MRq1pryrXzW/rESu5l3jvGPaKDexf+njF4cxgTPRPcrNQkA/eo+0kbjPMJSNe0ZfIMAoPAIDAIDAKDwAtCYASLFwTsFDsIDAKDwCAwCLyECBQSBLnhxd6sRF4RCCEv80gUv5ENyHgv/QgaeR0vHrcXerMUEQJIpc9Zyb4IiG04JwQBMkE+pIBnD6QHUl9+dfhd+CdtjBQprAMSB0FhBiUiDeHgNxLNscSUCLnihUeW1a5IIcSEvkR65NXRAqGOq0fbfSJbIlxaS6NwU4QVRAuRpHq0Bwnjt3p+ZSVeF8QMfTKL1MxPwoW+JExoNyLMrGGzQnlpwN81ca30L++Y7exP+/UBPgQe1/ObDvUhbP7T5YXxu+NlsZCYbRB4PRFgI9gX9gspy3aauS4MoO/sx81KbBGbygbJT0Rlj5H17JHzE5HtZ4e24YYegy4Bhe0ttI92GWOsx9PWWgiPqce5bO8574xT5cNEghebzx6z90jxxh/nsvtsd2GJeBmEPdzgvBVzjLFt58SKrRixbaM2NAaHofFn+67/ULGiek6JFX9jZfgLKxkjjXGu4zbsk/OtF3FzaGPPFPabhNB2bfuMcx9ayXUwNn7GoQB99TxBHNJWbTEWwsV9DHMik+/awtPRPeY/4D77tZX8N2DcM8SmefN1EBgEBoFBYBAYBJ4TgREsnhPtqWsQGAQGgUFgEHj7EUAwESO8yLeAqlYVIkoIIaQQUuBHDi/y2/ASQisg9okQZv4jHMy+JGggbRAGza5EGiDgEfpIrQh3+7XBOTwRkD/agmhAQCARItUi8/NWcA4CAhGEeCgGuPzKQl5EziFA5I0gaQHuZr2uQ3cbTBIAkBX1Rb/1sZnF8hauCaFxs5L+bmfowg1Zo0+JIvJaV8KnkCvw+cHDufoHI2KO8uSBO1LQorQ2mNyuBHO47UNVqMdCo9+6EhIt7xb9RsqJ8f1bS7TQNutZ/ONZy+KA7HwMAq8BAp/2ne964/e+4862sG3sN7vF1hFOEbZ/fKW83NhiNo89ZocIBuyIcH/seOWwJ74TZ59CtIioZ7MTx7/20JZTV0l/tmT/qXz6gZAm0rDXDxErlA0juLHDxoKtV0WEO0y2HiPtl7+1iK71PNn359S7e22Rf1v2Q+s5heN2v3vH+PXelVpfAs4/tpJ7w/icZ0xrn8Bmu05H2NxH+CL+SCYBEPxdT+cbV13fBAfH3MMfXUm73L/ubfeW6yYUmlBQxBTnKk+7C3M2nonX3AWTZxAYBAaBQWAQeEEIjGDxgoCdYgeBQWAQGAQGgZcQgWaHtqC032bNeoE3w9BLPbJdOKEvWwmRjpBABhADblYSSsTL/f+wkhf7bzn8RoI5F8EvecYw4xJ54MXfjFb1WjBavbcrIQ+QTcpEVsmPbEdoIPBbq0L9iQbKs6m7MBjaT4AhCviMWEOkIUq0TZnalFCyjSeu3YiTvCjkV452aavv8hd+qrBZxBJ9Q4poX54osFSe2ZwfP3wKfSUVG1vZ8NBP+4kS+gt7/dUm4U/US6hQR3HT767jIcTX+vquN37ud/9xs5MLr2UxUuISYu6vrqTv8BJa6t9d4sXHR7QA3WyDwGuDQGQ7+8LWI5zZNmHpfLemBXthHR627XsPtofIamN/2Be2JNt3u9l37Qz5awFn4y8JIdeIFerTbmK2/sKBXX3Ipt+wI/gow3hijSF9N6M/AV0eIjq7buxh2/WnMIMPqfvSOQkll/I91XHPB/rNw7KNeAAb49HXbPYb6wr1dew+4alIhLjPllBBIIHrdpIA8YGQYkKFcZSw9W0ruVbGWM8j1pjyfGCShuvomnm+aHLFfdoyeQeBQWAQGAQGgUHgiREYweKJAZ3iBoFBYBAYBAaBlxyBQitpJrJc2KPiXAv74QUe0ZI3QgS4l3phiVqcG8H11SshDZyPzPLCj7gXLqp9kfeIAgtM36xkFqRzlZWnh/MQGciC1nJoxq2y8iq4W2z6UA8SxPn6QWwwY9Kn81pcu9AcfqsPqdEin4kX8hA3IsgKpeF3i3LL4zyki77ovzUofnElAs03roSkIS7wYvjllQg7xBPEiHIIBoXfQuogUT5rJRgjm5Bv+q4tiSYEJdg6TrRoVvP6+pZNng+uxDuGUPFfrSRsBlJJWeJ6/8RKwlPx3Pinl2ihDb8zoaL2UM7vQeAdiQDbxY4mzrIzwtOxTT90sC0fWJ/WI0K8F/LI90RUwBgfCK7Z6uy+3w8RLdhhddjUw+6yhds1hZ7ighDIpYduCf7GF8I627z1uDC2FhqqcImteeGc+qicp97OeQNcs/bEQ9qzvdaw4KlgTSwCV2MaHExSMF4a605tvCGu3ZRn7HKPJJC0DoZjrYvVJAfX3LMN/N3bxtCPrGTc5j1EcBEeyn1ozHbfjXfFtVdj8g0Cg8AgMAgMAi8IgREsXhCwU+wgMAgMAoPAIPCyIbAWaV6T8t/YhqtANHl5N6sWCeWl34t9JD9SoJAfiHcEBVIe6W4WLmGicEiR/Uh4JA3iHkEgLyILwUNQcI5Zp5KyEBotNE1MsA9xIMSRGZdmxSL6leu4evK4QCrcroRwQ3hs141IdEgE0Sff9cdnfWkxbZ+wQMQpHxlCBMjro3jt8mjzB1ciBmgvIUf9yBLtU9YnVoIRQqQQWIU50R/fm3GLJEF0qQvR4xogf5QD39amiBA8Fl8b5maNEifU988sIeLjS5RQxl9fiWjyFSshlISAUZbr8++vPN+78u7DTK1Dsw0Cg8A7BYFDWKjWWWAv2DEkO9G1xYiFTZLnPYfjiFxks3fGQur4dN7tSjztiM9sV3b5vqLFlsjPo2IbNsglYNeIudsN4XzN4tv7sFHEZGPLtYttV+fWQwIZbjwyvuk7Utxs/jwp2nfsXfupwzQlmpzyRtGmS4tl76C9+PO7Vw7CAE9M3hF/c6V/bSVjt3WTjDHa5ZrByLh/bsu7cZvHOHcMK+OuMj23uC+MacZI439CGtwTlG7Xd88bBH/PFTwu3KPuedfRvey/kEfnrF9x4WLN4UFgEBgEBoFB4DkQGMHiOVCeOgaBQWAQGAQGgZcLAcQS0twLPGLey3zkQGszIAMQSQgIRIh1KBDy9iFqEPSOecl3TmsxtD5G3g/qEB9dPuRAIaa0wXlEE8QTQqVZkupDREUcNKO1MFPKimDXdseRI8iL2qN+ITpseW/IUzgThJj6kBWO+63t+lZ927jakVU+kRvw++GVzBq9WanZxkgSZFjtL9QWgiWxSB75iRktBuqzWanba6FP8IGjOk8JC/rGswOBiIz5Q8I+rU/71W1dDKEwzJp+30p/aSXX/utW+u2VF4mjrjdn/y4RY/2cbRAYBN5BCDRznC1hc5DsiHuiK1vMDvpNiEXssxEIaXaTbb05nJMtQkwbC+RnS9nx+woWwXuOyN+LFc65RqxgzwrlVz3bEEaXLq1xJGEjLxO22PgIk4R62LDThRoUQpHwfM27dqGSLrWl4wnfYe18+J8Kj3VKmDm1gPc17TBW/q2VhB6Ei/ugBbR5+cEh0Yl336lt23f31PZa7e8Hzx+Nl8Z9eeFr3IK3dsDEWMYj1P0BE/ncy8ZbWGgX70jjbc9Ayv2dQyPHu+LMBZtDg8AgMAgMAoPAcyFwzUPUc7Vl6hkEBoFBYBAYBAaBF4zAwcuiGZnIGC/pyA6zUBFWZvYTJd6/Ui/7LdB6u/aZlWhmpfwWs/zmlRAACHhEv1n+ykBaWYzbfsQAAsMxBH5CgVmVZl46T9nyIymUZz8CQt2FMkG8a1PChOcY5TsXgYSYQJpEgrRALJJC3rwr1te7PqtLfkSJchNInGcffJpJu/W+uFn7v/1Qpr4hfmCnfR9eCfmhD0gT9ThmprJQTGJrIwDNUoaJc7UPXsiTH18p0SfCsPU/Wg/kFKHiWgrtAruvXEkIKHW/67BehXL/pyVOmDFN3LhZyaK2f20l4aN+cCXH7kSLlc95vs42CAwC7xwE/L8Ru2wcTzDELsGi8FDWtDBT3fpEjtt4ELBTCd3OR8izKewo+1U4pKdGyhoF7Nm5Tag7fbCxly2qnUfepbUwtmUbo3imse0+I8blMUO/9Q/YW/3/3EPf2c4777aViOV7oeSUMHFfgeeYt4S2CLV4n+0xPACh+6+slOjheaAt4eJSW9xLxkJih22P1/Z8XhtEiW847HRt/PZ8YO0qZblW7m3PDbwufNrHW8iEC/d3oR+d5zo7l9DkfPdIa2RdavscHwQGgUFgEBgEBoEXjMBjHlRecNOm+EFgEBgEBoFBYBB4QQggTprFb7ammYte7i3IjOiJzEK824+IEvuZoODZ4WYlRIPZ+spB6vtEWiCxzDZF5CAJkPiId2QB8l7ZBJE8FnxXD9JC3epzvvKRCM0ORTBox3YRU/UhR7QJ2YHEqFxhI+xXhnqLPy6fOgrJpD3w0EZkBWLODNHIC2SSMrRJ0l790h59c34hneTlXSEQIcEAACAASURBVJHoQlixEQ1i/vWzmbf2EQ60T33yI960DSmWd0tx3S+FqshbBOGoT9ay4AXyFoFjiRD/5xIjfn7tJz65pvAXCuZPr4QE4qVx58kxosXhCs7HIPAOQGCFhfrk733Hmx0hkEpsuxB+7Bf7yg5J9rFX1uz5BysJKYfwZf/YLDaCvWOHkb/slfPZxFPks3z3VUH33hWEVV57tmblJ1bYl1jh+yWbeSjmLR/aVxv1t42N1lceAwQdx2Bj/POdp0ltPdb/+woTx9p2bF+hDq/Nfyqfa6ov12zGfltcwt67Y1vWqdBOMHJ/XeNhQuyX2kwGIDa4d9+7kvHbuEt8I0D8zGEfTwrjufHUM4UtryH3t31CorX1nLDZNV8HgUFgEBgEBoFB4O1AYASLtwP1qXMQGAQGgUFgEHgbETh4WSC3CwGEnEG4mJlvnYkEC14ByASkgPzIGkSF5wczSAvvhMhH3suLzJKfCOIcxEVhmogPyH2EvDIQXMgCHhmIBZ/KsW6FcxAaCRGICOcQLZBCCCPERGGmEA15XGgHcsmnhMhIVCmPNmhbZAnizjktjk2YgIM88uZpUYgRM1qRImZyOq/QIAi77WxTGCDQWsBW2xFMCBRlEVxgYB9RR9/V97GVeGMQRlwnZdaf9fXk5prpg1nJrpF2w/It28Hj4h8uQeI/OeTjaSFUipmz2vLfHdo3osU5tOfYIPAKIbDEikjzRMxCwLFlbN1fXokHHZH1ZiWCBFvF1rNHfrNZbBQbzB77rjy/CQhsvHzHtvuKFTw89utZbMPinZuVX/36GIEeeb5d6Ls1DLbixKmrqq/yqRfxLRmzCpXovESUFic/VdZT7uddsQ1hWNld52vEkmvFisrerw2y7Y/76csPO9xLx9aoKL92X8tJGA/dQ54lfMLffSc0o/uOCCEklOcPzwxEJNjIx0uyMFDGt/rbPbHFasJCPeXdOWUNAoPAIDAIDAIPQODah4MHFD2nDAKDwCAwCAwCg8BLjMAbS7j45FqEu1jmSAWkjpd+hBWCwQx8BAHSSLgLBLhPpDhhAtHgu/BGiHokASII0U8A8JyBoFcO0klCxNvfwq3IL+cgP4qBrh4EBBGAKIEcakHtZswiYCQEEuKiBbmd06LhiRbao86IrsQF5yR0qE85SAxEk34jPgg4SA8LcDsvjwwiAKHBzF4kiD5ojxnE1qjQb2UJtUSwIGwoV0gRXhzaw8shUQfe8ikHQVgoKW0uXvw1pJN2CislTAmhw3UprMv6+tbNYttLtGhtEqKRc/7tlYhX/8GhfZ9y3uwYBAaBVw+Bw8Lb7EheXS1UjHBnL61J4L/PHtmHGGYDkc9ssfGBjWicYLfZQjaQnWSvEMj33U7NsmcfzZ5nZ7N/7NS1m7YSwtli44p22vKW850tvkaskBf5zcbyTNMepPj3rfSBlYyb6oOBsaXFxK9t62Py5UW4r/OaMeMh9X7XOukbz5yYWCHLObEi/K9pQ+s4KS9PSuO06+c6ENRMDOCJ8f6VeDLCxT1sHDS2es5xjxMwPI+4V4377md5bU8uVqwxtucV/zH3hrbcPY9M2MVrLv3kGQQGgUFgEHgdERjB4nW86tPnQWAQGAQGgUHAW/kbb0RmRDp5+bfugdmxSKuPr2TGv7AXnhmQ+ggfpDtynZeBMFKIC4RQMxyRP4QI5XkpR+Ig54VuQAYgHuRXr3IRCsikFsJOFCAmIBTMjMzLIHICuRBJQwBInChWeSGckAPKI2JI2oOg0Hdt8FnoKG0jFthPZCE6RGwggrSjcFraxhuhNSiUof8Eixba1ifCgRAmyCybMngy+ISr84k/QlzAFOlCYNBmeZoBfZZ4QnoI33TIbx0L4aBcLwttC3uxnZV8aMr//7HO/b/Xuf/x+iocFOJNyJO/uJLr9J+fO/ctBc2PQWAQeBUQYMPYA/YXccoOIXpvDvtuD3aE7UwUfv/6zm4aEwiv7J1j7JQxQd487ZDD991O2TdeZ9J2KxzRtXUQGIguiRXOe4io4jwkOAyE0EOMs9n/6qYhxp/6svcMuba9D8lnzDq3aPlDyjx3Ts8Cx/LwOCGyX3MfnAoXtS/XWGgMNmGCWGRzHxij87yEt8kCxnnPBPJ/ZCXYuOe1CUbue88ct4fymjBxcoy8BN5h7N1ma3JDa5p4JlK+thBN9MezxmyDwCAwCAwCg8AgcAKBESzm1hgEBoFBYBAYBF5DBA5hoRArvch7gfdCjaD3om82rWNesM3At9/MfUQAwgA5ZeYqQSNCCflQ3HPsufIkxILynfv5K1m3gacFsoHo4OUeESSvOhEKiAft6DhiXz6kmecX+32XlzCCKFJ/xID2Kd8+5IDjrUuRN4cyWk9DHvmJDBE/iRwIGIScWZw8SgoBgrT5hZXkM+sTiUXogRmBRXkW/CQY6DOCC3ZEBOIGjLVFjG399lt7YK392oFMacbntTM/CQ0/stJfX4lgQlRyXc5tsP87KxVyw3X98ysRTz64acOFYubwIDAIvMwI8LLQvhUeyic7w14U4g+pX4gktoeNZefZPrbM+jhsAlvleIJzCx4bK3jP3WeR6xcJl/60UPNT1IOAZuONAdsNjsaQ1nF6UZ4Np/rQmMV+X/JoeAockO36fEyUgY0xkcfNpZBd2k2EuCRC/fDKw2vD/UYwUq+x3ThrHC/EpfvUBAATJjxjGPuM055HjK3uZ/dnExXc+/pxTbjFc7i5L4zbJiYo33+j5xvimGOtGaMcx2cbBAaBQWAQGAQGgTMIjGAxt8cgMAgMAoPAIPCaInAQLbz0R64gnRANZo0inJpFa8Y9ggAZgwyRmrmInEcYKKNwB8gMsxl5akQmIASQ5ma7eoH/spWQSQgWMw6JIUIwCZ30mStpF8JDOQiA1p7YLqzd7F5lO+4c+7RJQmIkRMiDHNFO+/QBidDaHNpeiIj19U0PB0ILXBAMyBEChfRNKyEkzE5G3n3lSkSXiBD5Yek3kgRZgTxBukRs8YJAlnSO/DDmuaIftrtFQF2rw++THxsvi8KoqAe59s+uGaD/6LBuxbli1PXBlVyjf/Nw7l9bnwgoXjWzDQKDwDsLgdbnYSt4eSF12Tm2kB1I1OVxxhYjf9m5Fpgu/B47yXax3cTP7Ndj0HrONSDu007jFduvvzBCUhtbjCmtNfTcgkXtfw6xQl3GcPfGVrAwlrtHbu4D5sp7SaxQHAHdGEiQyCPCebwCC+vkt+M2nqKeN1wn47O2yufe9nyiDPe8e9U9fHbbeFA0Vve84RlCiLJCinnuyMvGtVCH5xr1EvPgUxjIS9XO8UFgEBgEBoFB4LVGYASL1/ryT+cHgUFgEBgEXncENqKFF+k8CX5pfUdeF5scyY6Qatak2Y6IevuRV4V+4n3gZZ1HAeLAy71jyPpChpjxXygoL/fy+fzRlZBg8udxgfRCOGiblMdFpIAyESbIgBa+bqZpHhctjqo/iAuCR2GeEjqUUViJ9fVuQ3a0LgaCA/Hwz69kQXGkXJ4ff3x9zyvELE7EPoEFFspVhhmfPCqIPPok7BJypbBPH17f4Yl80f7CaOlza3bUrms/lfXdK8GBOOQaIAAvbfryKyv9Ryt980rugW9bhI1QVXC+2ybu9iUY5/gg8NIjUGgo9oa9YyMSmInW7DevMDYYKYsEJly04DY7x0YZG9jmQvLkmef8Qkq1btB9QHlo2Kb71HEu77FwRYUVbJyLgG7GP7v+HKGZYHxOFNHOa0UjBPp9OYEvOQDH28H4ZjM+bMUHRD3vwafYblYh7tMmRbhPPQfw2vTcQoAw9uZ5CZ/3rWTM0z9inIkAxvKPHs5trM2z81w7Ye35xPOOZwDjooXFCXjq4TWp/yYnyGf89Rzkf+Wz8I4XJx6ca8QcGwQGgUFgEBgEXicE7vtw8jphM30dBAaBQWAQGAReFwS8RHvRL3QSsoOw4LdnhRYZReAgKJBTCC2EiBd35DziQBktOorYQmg5x/le9JuJqkzkArFCHi/0wkoRQORVFhKBeIEsE96h8Ezaqg7n9d1nnhL227RL+1qE1HEbsUJZyo7UIWLUbqGokBPOLxwT0gOZh5hzPhEibAo7hZiQ9LfZm4QZ4S6ch9CCmfYgTpA8CBNECjyIIPIRi7RL+fB8KMGhDd+zEkEFlmaAnhQsNt4ZK9tdnRa6dc2E8OIpIzzU3zqUJc9sg8Ag8AojsEJDfXKFhWIb2DufZoSzg+wEO/felRDQPArY0q9eSTgo4e0cZ7eJwIRcoe7YxdaziFBuRvqD1wd4GyE+JjzAASFtM379/UP/7X8OoSI4LnlwXCtWKO8xfEBihXL2nhJPJVYo2zjrHnIv6nshltyrxAHjq33G3JtDcp4x1T1J6PjQSt3byvMMcHfv+y8E7IlP5fzllQge2mBMNPGAQKFdjfHKNKbfruQZ4u65YwT+C+jO4UFgEBgEBoFB4AgCz/lgNRdgEBgEBoFBYBAYBF5eBLx0t2hqBL0Xcy/yyADhDP77lRDpSPC8BJBciHjPFMI2RA6Y/Yj89wKf9wLSwPk2L/LNYJXXDF5kvoU6fTYzFymkbEJGIamKjV3YJ3UiDAoHoXyke14XfhMB9EM/tQe5hsTXfuQO0k25BA8kRH1pLQ9t4iUhLjZhwrn6wjPCTFL54FedYsJrHxJHHT5hBjvnwRKmzcyFdV4QZowq694k344YIST9yEq8V/6P5SVxluTanYtwNKMagQkfobrenPF8ZJHRdXi2QWAQeMUQYINbB4hdY5d5U/3kSq17g9zNswIZywOrRY0Lg0eEdW5jxpYEZ3fOxew/FZKHIHJsu0Quv+hLUP3GnT+xknHjOd+p87zr2hXaaN9vY8x++8G1Q0jDp9pcd+05thn/t5sx7dLm/pGOberhxai/xvfblYyRNyu5D43h1pFyj7qn3LPuXZt72T3t3naf+u3ZxL1/9n5aY51ra7wX9vEbV7KAu+cD+/Tx765kjP2+lXifEvuNm02SODRhPgaBQWAQGAQGgUHgPgg8ZkbFfeqZvIPAIDAIDAKDwCDwkiKwWYBbC1u80ku374QCZBNBAGGAGPCC7+XfS/lXrYQ8MOMQKS9MArKeN0XxtBEViAYEvnNbL4LAIJ8ykRTIBJ4GrVNBOFC2WY2IiBanRkTkeWBWpa1ZwspPlDgcuvvQF/v1AYmhTdrfs1CxxwkT8vidwIHg4eWBmDKjtFmVv7i+I0a0S5lEECSbRWotUKstt4e2ITTkMRNZf+ErFBTy5VdXIlZoi7q3QsVDPSxWMXcYwS1xRn9OkUvy380E3YgRhCukF8JGP/TfvnsLKXeFzzYIDAIvFQIW4F5eFsRJNp6NZCMQuURKHloIaSIybwv/e3bQMTaLgPs5K7Hh7GXrB7Ve0LavbOap7Zg3gDYRwo9tzykOnKq/8ETH2v6QEEuX7otCQPFwJEQbd40vjX/Hzkfg77c87oy11jd67GbcKvThvizj+HZzv1xakH1/TucTBmDAm8KzhrHUp2cMXj88NvMEUkdjPW8g51o/ynOE8do5xn/32P/TIvRngPBsUUhM97GyTCogjBA+/t81br7dItqZ5s+hQWAQGAQGgUHg1URgBItX87pNqweBQWAQGAQGgReFQAQ5Ytt3n176za7/cyt5MUdi8zQQwgkB4AUeiYTARx4g5W3IbaKAc5EViAMiBa8ERIdzkelm6yIQeCogUZBA6pGfF4JzkWYIc/kKAeG8LXmlLp4Onm+II3lebL05tAm5hsj/oZWEOUFwCMWkLQi4QlvVLm0gLBBi8tzQJpv++G5/RL4Y2UQVsa4JO7wTzMYkUCCYhFkyS/O7VtIe58KiGZmPESn2ogMcYaaN+nWfTTuQY9bCMLP0r670/SuZRfpJwsaEurgPnJN3EHi5EFhiBTLW/5xtYDeJyQQIZDc7Saxlw9gp9oyttLaNPGwD22hfNpOtTzx+zHsm+33fLRHhvufdN7+xSx+3Hn2VATPjyFNvecch6WHuml2q5ws3jdiuaeEaFyrxse00ju231nfa13FMQDlXf+I6AS1PRPcX8cB4nFhEPLBPf60pYczjHeh5hIdhHpvGXdgR5+S5C7noP3BBtJBXfZ4tYEfE02//ARM0/uEaC4klbxm3Z2x87K015w8Cg8AgMAi87gg85kHydcdu+j8IDAKDwCAwCLyTEPCyvZ0lSAhAiCACkDBmEt6uRBTw0u/l/0tXQqQgsjxTFMbIPmRA6zogCLzQIxuUS0gwU1dYBTN1CQG8M4gSSAEEg7b8/EpmTqrLbwQEkogg0oxHwkBhoxBW6iQ+WBND+UiNhACfwpk4RjggJCDbiAnEF6SEPPrR7EkkC+8QZSN94FR4FDM19YsYAKNCJskXAQgb+2ElD+wIIUgvbYWbtsC1UB8JHw8WLnZkifLOhWRZh//JtvOygLu2arPrhKw0yxc+d94YQ8y8Bb75MQi8MggcPCzYa3aPzWKD2F82CyHLVt8e0mevT+I1W8aOI5Kdw6ZJhYdixx1HMkv7rfUtnhonZPJzbMauxgP2m71PYDnn8fAUbYMrYp49P4btqTr2niCt9ZTnxmPatr+eYcGjIS8Z41vhmY7VRRgjNhi73XfGG4KYRd95NSQI5JFozHbPeW7wzGC/66+fHznUe3v4vDmc37OLe1yb754LrvSwUL5yv/3QJnXq29ev5D9hEoV9b647lafijI9Qnm0QGAQGgUFgELg/AiNY3B+zOWMQGAQGgUFgEHinIhBBjqRu5i2CBGmPfPgHKyHpzbZF2iAVECcRCvZ5YUfM87RQjmPOzeNBfkQ9UgKBgXCQD+lDiBBOyW9lO6YdwkR5ZkESRYYh1RAQYnIj1d63ErKCeIFQs6/ZvgSF2qkO4TD8dv7NSgQKJIY2C4FlH5IeAaI/ZlMiTAgX2oOoI+YgVBzXF/sct2m7diAx9Ot2Je1Vr3KFjZIfJkgP58E+0ejBQsWh/kd/7EQL2PBG0S9C0f/X3nmAWVFkbRgTqGDGnDAgIpIFUUHABAoqYl7FVcw55zWuOYA5JwyYc44YEZCgoph1XDGnFcEc/nrv3sPfXu9EhmHCW89Tz73T3VVd9XZP98z56pyzQarX5ec+w+eyAwlIYNYRyCffDm86BoIhHEESAzLP1PAgQ6jFyIuHHMbZyOWDRxnPUPIQsY9nK+8MjLzxvM5OsDLeEzMjvFIhbJ7tPM8rk6iad0MIJJWZT3VcaK5PoTgT75OKCiaMmWuG11+vSg4q663BPUG4wy3yDLP7siG9ygsjiJcm73Lum9Xz1wIBjL8/mBNj5e8I3tG8h3i34z2BtwPvZP4mYUEDn7yvGBeVfdyDbOOe5p3P/cnPv1VArECQx5uQ8/O3D7V/qkflx0leC/5OwfuTMI94dpSkyr2fWwCiqA8FiwQkIAEJSKDyBBQsKs/MFhKQgAQkIIH6TiA8LfinHgMARgMM7mEoaZG+Y4B4LFX+Ucegj1EAww/GBFbgY6znn3b2hVcEBiEM/OE5gfEAgwIGfP7pj9WSGF+65I9FeAjxhBX+GMxLUsUzA4PaeqnSL3/TRB4Kzv1JqsT55ngEgVh9yXgJq8E5GB99Y5DD0Ea/jJW5InowfwwiGPM4FoMH32PlMas/MaBwPgwuGFYYI6s/EWNidTKrRglbgaDTIlUMJhhcMILQbxhZYFprYmFnVoZisMHTBWMSc26VKiIS3ioaZIBgkUDdJhBiKQZnnlX8zCp8BF4qwgHPaZ7fPNcwKvPM5znGc4DnJm143vKM5T3Ac5VnaPy/WRXDfk38r1pa3oSKXlGe2WXl1agOL4YYS4T1K2TJOysruMCexQJl8eN93qvIJHkncR2LFe6P7DuKdxp9RHiq0kSfsnKY4CmxfqqIAdw7UXj3Mq+YA+/WSODOGBBEeGeumirz5RrwLqbCh78naEuf3LuIbLz3c3OoiFiRGQvvbEJUUvk7h7E+nSp/w+ydKl4v3PPMk78PrkmV9354d2a68qsEJCABCUhAAhUhUBN/BFZkHB4jAQlIQAISkEDtIhAGLP4hj7wNGAQIs0RIJTwFIl8EKyExXEVSaQzwiAnsZzteCxgU2qeKYQNDCT/zHWMCBiP+JmEbRn8M4/zMP/8RIipCNTEGxoRRLZLEYsSJONMY2TBkICQgnBDqicLxGDLYH4YFxoloQFvG0TVV5ooBhXEwboQM5sDPz6eKoZ65YfjAiE/BaNMt32+EvoowIXwS7gJDC/1wLJ4ZiB+cN8I18X2We1bk51Psg3ngZYHYxD2AUYY5lJnEu4z+3CUBCdQuAjyDeJZSeS7h7YbBmGcWBmye7x1T5TnNsxVhluci26k8Xym0xWAcOQx4lkcOhpqccXUKBRUdd7FzVuc4YMm7DPbZUigUcBxG8xapEraovJIN61SaWEEfhefhOsffCmWJNrwnSsu5UZjbIvKA8J6O8JKMj3d0/IwAwd8N4R2JyILHD+/YzVLl3Ry5LnhPcS9H6EbmUal3bd7L4sHUDvGO93/PVPGYxEOF67FLqvxu8PvA78vlqQ5PdViqLJioNQsRmLxFAhKQgAQkUBcIKFjUhavkGCUgAQlIQAKzhgD/1MeKTv4RRyDAMBBhn1htjzgQhn0SZmOsQmRAxMDAwCfGCjwQ+JnjMVDwDzwGjPCKiMTY/PPPOfhk1S4GEYwTeFTgMYGhhu0YIzCQYEhn9SM/I4Twtw1GBYwGEfea4xAhMG4wD8bBOTBA4C2AYQ2PDPpgzoR2YPUw2yMMBOIJiboxkhCagpWWGEHwIGGO4YVBP/DBowODBu3JY0EbxsM+zs2YwytketzrtK02F8bM9UWsgU3EHK+U8ac2T9CxSaABE4jfY4zCPJ95bsfKdERKvvMMxUMNERbRmpXxrHx/OP9M2Cbfluc57SOvD88N+uVZXFPiRWXOU5qoAAf6KauvrKGeeVbX/9cY4DHaZwvn4h3IezPCP8XYEeARkngn8b4i3wIiO+8kvA0o2XbZfqvi/RLtOT/vhLjWBUPO/VhegvBoE145jJd3bSyWyIVwyvfD9rtT5X3K/YeI/mSq/F3A+5wk8SWpwidE9cgPxXn+rKR3RYyN9zThzwiJyO/AvUnI+DR5H+JhdGSqeB3tmyp/G/D3C38X/CvVp9Mx5L/gev5NuDDHReD1UwISkIAEJPBXAtX1B5VcJSABCUhAAhKoXwTCeBVCAv9o83cDhglW0kbOBkQKvBYw5iMeRDJpBIY2qSJQ0BciAgYEtmOwx7jBP/Z4MISnBNswWCAW4EXBP/z8k4/RBQGAEBF80g9eCqzyR6TgZ8aGQZ329Mc52Yehgu0YTDBwYLyhTwxQEW8boxCGpkh8zc+sJEV4QZRA4MA4j6EEox0rJjGoMD640A+GIoSO6AvBBCMQhg0EnfGpYuzD6AE7zhc/hxGjthv+GR9GMYQjBAsEnrgX0leLBCRQDwiEAZ7nJs8unp0RKorfecQLnvk8x0nEjccdhWctz2Ke+TwnEIkRbHmW8rzleJ6xPN8rWqrTOyHOybM3ckDEc5h94RGSHVtWrODZDZvC/595jvPOYZ4hcET/jL8sz4OyONAX/CNBduG4GDtCONeG9wwlKxpwrRgT7+QQLCqa46Ki14d7BG8G3neEUZzRghgT+S4ir0jkr+BnWMA0vDVZDIB3zwv5fXDnvY2gxns7wi0yTgrXorx8Gn+bQyTQTjt4d9M/510ubedvGMZDnwgnx6TaL9XdUmVhxgqpHprq0FSfSvW5VPk9qPQY/jYoN0hAAhKQgATqOQEFi3p+gZ2eBCQgAQlIYAYIhLEoVttiDEAQwEDC3xAYA8ak2iJVDCEYSzBQsbqTnzHus/oQoz/GkxAE6A9jPkYevDQiATbGFwz/nCeMZBgrED4whiFcYATjfGEgQERAOAgRA8EAA0YIFuHNgOEGsQLhAMMUyTJJ1M2YY0VxSX4seEYgsNA3IaAitATjYsyMl34RLuiTeTFXBBSMcRhVMIxgbCKONf1i2GAMrLxEOGGl63SjxWyzzVbbxYo03Fxh3lzTtVMl7BZ8xsVOPyUggTpNIIyvIaLyGeIEz3ueYRiCMYDzDODZyzuBZzTPXhIdI9yGMEt/PBd5L/DOyOYoqAgozs9zt6yQQhXpJ44JsSKE5vD6yCaxZh/PdgRvanhX8MxmDoX/PzPHyPcUuYpglhU7suPPCiZljR3jPR4CxQQL3sGMB6EgwjTxLiv0csADgfdNsVJVMYh3MO9Ezk/h2vIerK7CPYS3BAWBgHcrXOGOWMD7HS8H7jsq9+COqWbf9dyrHM+1pC33I39LVNW7grHAi79PEGgI/0QYKP62YQFEFMZ3S6r8DbFnqtxXLVLl75x1UmVc16X6SH5c5oDKwPOrBCQgAQlIIEtAwcL7QQISkIAEJCCBRslgXhqFnCH9zz9zH5FvAWNJxC3HKI/hGgECAz/GE7woCBMSyS7ZzmpD2tEHRiAKYRII4cCKXdohBvC3CWIFhgB+RgygLW1YzY9Bhv0YwTgn+yPPBscwHowTiAqMAfEEowV9YSxgP3ktMIogKmBowTiFYQSvDYwf9IOoEeeKnBP0xz7mwTkw2mG8waCCwMHcmDtGCo5hRSXHIaYwvxhrcKgrIkUjwlZkVplGyCzEGK4xTDAGWSQggbpPIJ5LPKcoGLx5fmFA5xn6WP7Zt2365FkcoW54ifBs4LnK8xlhk+chz+CeqSJoFOZeKI9WCAkzErIoe47ojzEyz/D+4NkdBnw+MXLz/OfZhocCz3CM9NEeAZp3DO8mxAjeA3gL8q5jniHqR58cQ1vOlxVHypo/x+HZV6xwHgz0pSW5zrYpLSdFZUJm8Y4PLw6uJ/zoN7we4MF7tKzk2mXNlX0Rrop39cT83BBsECV4H3NPcR7eNVyXyEHFPYVww/uW9zlc2MZ7P8Iwcj1mRKyIsXMdub6INB1S5W+XrGDBcYyPsFTMAZHi2FT599zeqgAAIABJREFUW4F7ASHmoFS3SBXPC/52sEhAAhKQgAQkUISAgoW3hQQkIAEJSEACFSXAP9wYE6gYePjEqIIxiZ/555tjCN2EuMA+tvMPPsZ6DEAYDjA2YHjgn3oMQxgBIs42BiD+4ccQgNGBc7yVKoIC21nByPboj+8RcgMDBcYKjEdPp4pBjXjeHItAgeEpVoYSwoqEmRgeCGmCMYR9GDiIRc24EFRY3Up4CcaAcYi5MF6EDwwmeIVgsIi5YgTCuMInc4cNc2b8GLgiJ0idESvSmHMlI1owB67Xxvk5wZyVpxYJSKB+EOD5xPOUZ1gIFhiFeQbzzORZj2cVz0qe5zw/ESd4xuN1hZGZcDg8cxF8eT7QF4b2YmGVyqNW1bBKZfXL/8GMied6bvV9qpEbifcKz27Oy7wp8d7jWc+ceQ6yjeMiyXgY7NnHe4JnP+8MhF3eQxTaF84H1hWZI+8czkEfjJXz066stpURJvJD/MtHzCXGGJ4L2RBaZYX5CoEhOo1QjIXn4l5hUQDzwhMycnIQaio8dAjFxGIGBBS8Fvg7g783EM+5J+NaIjDRH/cu1/iPKuatyI0x8+6DwV2pMiYECRjMTlJujsuI+txLvBcR9whXxd8YtMEzgwUT5HohnOYeNEuV62iRgAQkIAEJSCBDQMHC20ECEpCABCQggcoSCGN8rF7E2wIDDqIA/8DH6k8MFS3y2zBYYdBiP4YGjtk6VQwtrEyNFasYuTDsEA+a7xjAWHmJMIBxgu9UjACRXBSDCkYJDAQYhhgPcdQxZGAAoT+MH7TDgwJBg2Mx/GAIwViA8Q3DGu3YxspOxsQcWUnZLt+en5lH5MXAswLjSEmqGK0wtiB2sB/DTMRtDw8E2NU5sSKNubDAAKMe82mWDDUh2OSMOxYJSKDOE4iwSTyvEFwxBrNCnOcoq+kxEPN8ZhtGV56DPLMjATNGWo7h3YDRn2c0z1m8BnjuI2ogbsyqEiH+OD9jD6Nx5DcqzGnBMxwjdZdUeUfQhmMRJjgWQzrvQAzSnfPbsp4hvJdKKxURK2gLW86BUEThf3nef9nzFAoEM8qXseFJwTXnPHzyjlu1SMe87wo9OsKjMg4vzSsEphTuOzwSWCzAJ+957jHuF87LO537inuOvljEwM/s5+XD/clxsMqJSjMiVhSZI15EV6TK+4+/C/i7IecpUeTdlxMu0vuRRQ8skmChw5b5Pvm74vZUj0n7H06f/I0yvfgeLULeTRKQgAQk0KAIzOiKiwYFy8lKQAISkIAEGjKBfFgoEERs7oj/jTEDIwOfGIH4Rz68DDBgYVTACwHvCY7DwMAnBi2MOKyExKBFe1busw8Rg1W7tEV4wOjBqkuMShi5MNgQTopCe4wbGCoQHBBDMCJgtCCMRRhQEE0w9pTkj6U9RgLGi8CAkEHfzAFDCYaoGBuiB31ivMF4wifHR/gP+sY4EYm/Mc7RnuP4ZE7sj1pWGK50WO0tmVWkiEPEruda4y2Ti5WuoaX2XjtHJoHKEvh5t9wzjGdi5KDgeYkRmdXiFJ5pa6QauYP4OULxYYjlGcF+noG8MxA5MGzzvC80Zld2eNVxfIRtyvZVLGdGeBcybgrvlxDKmS/vEraVpMpqeuYW3iSVVXF5TyGuFxY8C3gPElKoJgvzGpnqevnrVtE8HJUZY9Z7kv5hh0AET/KlwB+xJArv5LGphj0DAQM2IWzkPGKSWJHzfqiOkn/3cT7Gc3CqXONrU70n1dx5ir3/Mu9MfodIVL9TqoSEosB2RL4/ru/04ru0Oq6afUhAAhKQQF0loIdFXb1yjlsCEpCABCQw6wiEh0AY3xEKMC5gZOBvC77zT3iEimKkCBFsY/UpK0BZjYrhh+SUGPkJkYChIRKJEhIK8QEjOH0iaGD0wijEqknOjQcE/WIoQ6SInxE5GAP9sqoRw0aLfBtEBs4byUoZMwZ3BA9WzLLKE5Ei4mZjSGA/4RvYjqCBwY5wUiWpImxQOD7CPXFejCUYMKJmmeWb1PkPjI4YbLjO041CGGc0tNT5a+sEGhCBJEqUVrKL2/jOs43nMc9CjMmUjfLbeB5G/goM9BiXWYGO8MxzluczffB85plNP8XEguxYKhoqqapXi1X4vB8itwbjZ3y8Ixgznn2EOwrhId5zjAsRh3dGPNuZE/PjXcQzkX7ovzDROO+K8nJ5FBMrmCMCPH3CsqwwTFXlQbvIJcX3EJmYD56RIdZUJA9HedeW/uMYBCLmxLkJ78SiALwX4cTfC4wDrpGEm2vDAgjev4RdonBPcs9xj06/b9O9PVs1e1gw5vi7gjHw24NwggdoeUm0Iz/Hv9OhL6eK2MHfF91TvS3VvVLFu3R6iCnfpfmr64cEJCABCTQ4AgoWDe6SO2EJSEACEpBAtRAoFC3CsMF2jAYYNDA08A96hF5iH+EUwugQccDxvuCfdAz+GB0IGcLfKBFaCe8FhAoMFggK9IshiX5YlYlhg3NyTKxqpS8MSBxXkipGjMi3AYAIaUJ7VvxiAOEYtuPdgaCBkYaxMRZCORD2gT4wODEXxoKhhTYILRHjPPJ75ASdlNC8PoSAglmuZOJ5M1+uDSFSMBzx3Vjc00n5RQJ1g0Ay6JZW/syLGbHinWdhhNzBcw3Rkmc6z8WXUg2DNoZ1BGcMzzyTacdzEyMtz1kEYMRoDPNlGb8rGiqpqqB5hmMoZy68L2IszDc8ASPkE+eIEH8cy1x53oVwy3fEjxAsmDMMwtuO9rQpT6woby6IQBFysCJJt8vrL/bzDg+DP8/zrPdIhPsq7KtYPgreuTBBqCrmQRPJtekrhAWOhx9ejIgBG+Y50h6GXBfe6REKij5473DvsQghQjGynfctY6dWR6LtYvy4l1m0gKcn9wKCw835c//t+BAd8p4WjI+/XTieBRsHpspijK6pDkn1iFQJnaZoUYy82yQgAQlIoMEQULBoMJfaiUpAAhKQgARmjEAyvJfWQc4wn0rE/saIwd8YfIaQgaEGYw4V4z9iBCsLMYQQmgnDEdvYFyGcMBRh/OFnPCAIl4AowYpVRAvacx6+Y8jg/PSHESfOhRGEfvDowMiDAST6wKiGgYMx4qmBWEJhDBhsGBNji3BRGCk4lrFQ+M4+zhWrQMNgX++EivycCz9YVUr4Eww3GGFgZ5GABOoJAVanJ9GCZzzPNj4jpxAGYcL18fwjFA/PWJ6pCJfPpIrRmWcCRnDyDuA1x4p0BGae3Tw7Q8zlOwIxz3MM0Bw3swpCCe+VKBjEC0M2IZQQ7o9P5heeHhzH+4TnHO8H3icRGioSdjOHSKzNJ3ODDwb2EHRmdG6F+TVmtD/aM1euLeGoMMKHSBUvfvIW8T7MikghmCDsx7ue/E/ktygt3Bfv6CiIEMGLNlwbeFEI8cQ9xTlg+3iqnAeBib8FECs4ngUG3FMITNxvkWOr2kJBxWAzYj337R2p4nG5QarcK8yXe6NUL4tMew6D75hU906V8FD0A7ujUz071dGpVvscYi5+SkACEpCABGo7AQWL2n6FHJ8EJCABCUigjhDAkyCT5wKxAsMBRi6M+WHY4J/6MOojALACF4MRRgzaIAbEKt4wgmAkwsCEcQJjBe04hn4wbLEdAwbHRCJo2rIdAxoGMwQJxkAbjCQYkjCCRJgJRAzOzzgYAwYbvrOffZyTQnuMVZFEmzYR/mm6J0V986rIz336R8bwgtEFwxHXMQxcGlkKgfmzBOo+gezvNcbhnHE2FbzRMOoToihCB7GN5+hbqZLfBi+2XVJFzOB5zvE8j6evhE/fec7SbmaXrFjBubIJq+PcvLvi/2T2Z430zIsaIgZ5moIH4Yk2TpXnIe8YjkGA4X1S2TwWMzscVjHOvBMR7pk/q/6zhXcr79LCEFccg8GegoCN2M/1Lq1wT/BejlCCzJN3Ne9VPC14l9P+gVQRxEhOvU6q5H6IcI3ca9w73C8IFixYoG3cozXxDuJvgqdSRWhhDFxzxJ4yPSqLhHiakjwvrkzt2qdKeDV+r25IdcdUETRqYi7pNBYJSEACEpBA7SKgYFG7roejkYAEJCABCdRpAgWGegSMnPdFqmHMjhASGCsihAYhJCJsBoYL9mE4QVhgH3+v8B2jEdsxdmDQYPUlRgPCSGCsYGUmhiNKCBN8Il5gbGE1JEYxDCIYZOgzew6MSvTDGDA80I7+MK7RT+TkwKDAnKbnqKjvAkWeaWkfGKC4RjCGVRgyy2nmbglIoA4RiGd5rGDnWU5IJwy1PIcxLCM+Y3TFOI+oy4r8WHmO8ZlnLCJzhFbiWcszlmc6+yiI0jxLaiohd3neCqWNI0QMxs17BC6RA4M2vNMo9J/1GKmoEFGRcFhcAwrP31JdINM+rh3XKIQFPCk4vtDjg3Ej1BcLW8W1La/gSVNWQXCIvBSRt4Ix8a5FCEHswMuABQaIQtxf9Mk4e6YaSbf5u+DVVCP0GO/r4B33aXljrdL+jFjPdSQROdefe5YwZ7z/+BujsgXBhfwVx6c6MFWufe9UyRNDnxYJSEACEpBAgyOgYNHgLrkTloAEJCABCdQcgbwh//ekW0S4CE6eiy2dasSlxtiAISPCZ2CciNAbGLT4hx2xAKMPRg7ECowckUOB/jC0RBJUzoFBhp8jqXaLfBv2cS76wkhSkmok7Y6wVRgcMLbRNrwxYiVwGOvop6GEfWKufyuZlaK/pBWiGGwwzFXEyFa0PzdKQAK1nkCsHsdQznMZsQEhgmcmRleeqzx7ETEImcTzgOcqz1GETVbE0weG5vCkw9MCA3QkmsbwW1NiRUWAlyYw8I5gXggBvK/wtMC7Ag585/1DJZdDVkyozmckYyNZM8ZtzlNYeF/Cn/OHWMEx2bBM/BzhvsJDhuf5zCich/uFsfC+gB+fiF3sgyX3Ft4W3AfcG5ELhfuKCj8Yc8/RV3ZRwUwVK4oAIQTVs6mSkBymjLUqggVdw/yYVMkFw9zpb3Cq5LqIhRhFhuAmCUhAAhKQQP0koGBRP6+rs5KABCQgAQnUNgLZMAnT8zykQeIVEaGjwpOCsBIRixrjBKtxETXYz/EYtzBsYAxiRSYGjgjFQDtKnA8jTqz8J2wDx9IH7SNhagglGAxoT9sYEwahiN/+l9AMDdyrovD+4ppgXMIAZZGABOongXiuhsccn4Q84hk9KVU8Klghj5iBETryFEGDY8n3QJgbVs/z7MbwzDHhkcEzJDwtagNB5suYi3kc8C4hvFQ2xNRK6ecIDxWeG9n/twvFD0SPGRFnaDuoDFCIFRj5KbxLC88V+UKyY4zQXtXFn+seycwRKrg38KaABeMhTBgMuRdYRABv3iPcC4wfjlwHknHznsHLgnsN/oyf/ukrFkKUGZKpOiZVkMuCBRDwYw4ILYg+VX0PMvcbUyWvxcH5PldNCwLwvIBNrhQJK1Ud07IPCUhAAhKQQK0iUJbraK0aqIORgAQkIAEJSKDuEsjktiicBH+LRMWgEp4YGCvYHsYHfsboEfkwMFZwPMaVWHGJ0SBCZES+CgQL+kSM4JPtHBMhO+L4OBc/c84YS27FpuJE3b33HLkEJDBjBFLS7cLC85HnLavAI3wfz+aOqRLCBw8LYvBzHM/QCJUTnnEj0jY85SLx9ibpO0IFQkYkr45zIoawrTYXVtUjuvCOQiDAkI4BG8N85G+aUXGitPnzziovJNSsZIeAFd4H3AsIOvCJ8IxwIgQUP/fK84oQUdwTvJt5d2PIpy0LGkjIzTsccYD7A+aRS+ovc01J42d6SYIC5+Dah2j/R2VEhXz77Dj5Pbgk1R6p8rtzcaoXpRq5sxQtZvpV9QQSkIAEJDCrCehhMauvgOeXgAQkIAEJNAACyeBf2ixzgkBe0Mh6MIRogBGCxiFQZIUMwl2wIjHCS0VYC87FdwwIGD5oz7HRlp8xAkQOCtrzN1H8TPvwrKhzV6dx4yZNms0//wLffPUlqz1nqCzbYsWVv/7y889+mDYNo5BFAhKQQDwfecZGPp8ImYfRGeM0z09yBa2YKoZlRAyOR6TAyIxBNkQPQuAQDgrxAmG5Rb595FcoTazAG46wU5TIjTSzr85D6QQbphoiRJyPuYQXAfPH0I6hvmWq4Z0xI54UZc2rcCwzwgDPw2LeJFXpM+4JPGkiZxTvWsQJ+LCdewKvHAQH9pHAGu8E7iPeybzD+Jl7ie+8z9nHNvrHgE8tKlZUZdBVaZMXJ2K+le4i47ERbRFmTkr13FTbprp9qs+kOrbSndtAAhKQgAQkUEcJVGcMzTqKwGFLQAISkIAEJFBLCET8aT755z8bOgoDGEYpDGQYtsITg+8YrjB4sC8SafOdbeyLsFO04Tv76CsrSnCubEiJmR5WYmYwnz2Vq+54+Jnjz7pohteVduyyVvc7nhz92vIrtsSgVCdK245rrPnQi6+XNG3WLBumpU6M3UFKoI4RiDA88ZyO5ysGaYz2LDsnbwXhewj7MzrVt1PleIzi5LEg3M/qqeKRQf4LBI4IBVQWDp7PrNKPUp1G+7LOG+MrPCaEk9hOLoM1U8XrIgrvI0Ia/SW0YFknq8F9CNLUwtwWlR1ChJ+i3eOpcu3Dy4Z3LmLVyqm2SBXRatn8Nu4F7gnuDe4R7hXuGdpzD3EvMTburXj/c47cezt5UfyBJ0WxWtkJzKrjCzwyuEdeT3X/VBEq+Ltm/TyD3BCLeGXMqqF7XglIQAISkMBMIaCHxUzBaqcSkIAEJCABCVSGQCkeGNNFg7wHRggZWTEh4lcXO10YhuKTYxulc+V+ps/6Fuqp54abbIbRftRzIzAWVbksuPAizc+45Npbfv7ppx/fev1Vwm/UibLr/ocdM9vss82uR0iduFwOsu4T4JmKMTXC9mD0xnuNlfokI0Y4xBCNwRmjPuF8eH6PSrV7qqyWZ+U8HhZs5/jvU2XVfIRTirxDWVEAYzar8aujkIOAUFUVWchX3jkjyXWxcWFwn1FBoDrmW6yPYl4s5YXi4joVCsMsEMDrkeTq5PPgmsKE+4R7Aq8ZzsV1x+MEozxCFZ43z6faLVUSaSNETMx/px3nol+uVfbvgPg+s7jUaL8Fnhb8nULerZNT3TRVwkMheBEaK0TCGh2fJ5OABCQgAQnUJAEFi5qk7bkkIAEJSEACEqgSgQJhobIrVIseX9/ECsAO2nP/Q/lMjhYRnqTSvBOX2U4ectl1iy2x1NJPPXL/3X+kUulOZkGD5VZYqeW6G2y86dUXnXNaxBibBcPwlBKodwTKyAPwZ8pvEc8HnjmIC3hNsA3RAeM04aAQMUpS7Z0qq+zZ/1yqGLI5Bm8J8hEhbERyYdpjyCZ8UFas4BwYuaurYFyf0YJRPUJeZfsK74K6mDeyvOTniBWFAg3XnuvLtWPOcAkxhOuPYLV2qjAnyTbXGxEiONGWPvCwwAODe4f7gf64Z7Bd4GHB8bkFCOnerJPekKXdcEVEC8JDIVx0TpVsMq+kmltEgJdFZXJllHZOt0tAAhKQgARqI4GKrCSpjeN2TBKQgAQkIAEJSEACGQKrd+jclTBObCI0VFXh7Ljbvgf3WL9PP9qPfu7pJ6raT023227nPfdDqLh7+LAZDodV02P3fBKoqwQIx5PGHkbjyCvE6nhyOLCSnjA+5KbgOwIEBmpW1yNYUMMwjffBG6nSH8ZwRAqeYxF6KhAR/qnKz7eZxBkvEuZRLLcFHOpSicTOFRFZIs9IzA/hiWv4bqqICwhLhMVCtCCcFh4qhHxClGiRKqGzCHmEdwX3BPcG9wj3CvdMJOOGIfcUXhbcY5Q/8/deXWJblbEiWODtwu8DvxeDU61t939V5mUbCUhAAhKQQJkE9LDwBpGABCQgAQlIQAL1gMBOex5w2NTvp3yHR0RVBYvWbTt03v/oE08PHKOfH1EnBIt5mzZtttk2O+z8wojHH/5k8n9K6sHldAoSqGsEIgkyhm5WzxPGh/81MU5jbCYBNfkIqOumumeqhK5rkWqs1Oc7RllCCxH+ZplUixlnEUgwXhM2KltCFJkZ7DDk0z+eIJUpYWCvTJvKHounQjZfRmXbZ4/PJgd/M+3IhsHCu+G9VNsUuS6EBkOY4JrjKcF4uEYRJorrSjt+joTthI1aJVUSmXP/jEiVnEnMZ1yqJJwuyZ+TdiGO1Qmvv6pehMJ8FsmTAo+TS1NtkWrPVBHHEHT0sqgqZNtJQAISkECtJ6A6X+svkQOUgAQkIAEJSEACZRNYetnlV1h/480G3nfbTdf9khJPpIhQlQ4JNc+88zY94+Jrb546Zcp3X3z2yceffTL5ow/ff5fVsLW+bDJwux2bNptv/luuu/yiWj9YByiB+kcAASEqs8Nozep7DNwYvWNlPKvvP0z1xVQx/G+XKqvsMVY/lOqYVDF80z6XUDmPCgM1YaWi8HOxZxyr86u7sLqdgiG/tOcqYy6tFMsPUd1jrC6xIsYVXhaFOTsQn1jxXygY8DOCAqGKXkiV60gfhHPCa4JKYdvIVLnWtOHacw9wL3BPcG9wj4SnDvcO9xD3Uiy0zN1n9S0UVDk3BOIfLPA4IaxWh1S145QDzd0SkIAEJFC3Cfiiq9vXz9FLQAISkIAEJCCBRjvstu9BsyW3ituuv/ISclBUxcPiiJPOOp88EBecceLRzRdbYsnRz9edcFDb7LTbPv/54L13XnzmyUe9HSQggVlCAEMyRuioGJpJqI2Bm314J0TOCgzSr6ZK8myO539SjkUgxWhdkioGcAy1JGEemypG7kg2jOEcI3Ykc85OmNX5VS2RPyPbPis4lJbvYlIZJ2xeicFkhYCsQFOJLqrl0KyXRWGH5CHJRmngOrHan+tJ6Ca+41HDNeNaRP4JPDPYj4cN1zrCfXEP0JZ7AtZcU+4V7hnuHY7lXpp+bzUwsQL+zJ1wW6uniqfKWqlWR+6VarlZ7EQCEpCABCQwMwgYEmpmULVPCUhAAhKQgAQkUEME5l9gwYU233bQYIz1eERUJeH0+ptsvuWA7Xba9f7bhw+b8t9vv0HwGP1c3QgHRd6Olqu2aXvWCUccWJW519Bl8jQSaAgEwsuCxNiRHBmD84+pEr4JYzaiAN9JqEyug4dTJfQToYHYRqLmO1PFoI1hFnGC/1l7pBpGbViSLwKD9qhUl0+V8EFRMIKvUEHghNtBKCFcUacKtik8rHUZ7cpLXp1tml1MWJl2VRz235px/SqSuwJRCc8TjkWwQOBAmCHUFwmi8bQgpBMhnxCd8LjgGu6U6rap0v71VAkdhtfKyqkiWiBOLZJvw3fymnAO7iXuqYbmWZG9QHAmLFSvVAm5Rb6qu1Ot1+GxsgD8LgEJSEACDYuAHhYN63o7WwlIQAISkIAE6hmBLXccvCc5HG66+pLzmRpG+8oY7hdbYqmljzvzgis+/ujDD848/rD9u6y9LitoG415/pkn6wKqrQbtute0qVO/JxxWXRivY5RAPScQnhZ4Q2DUxthMyCJWzscqfMIGvZzZzj4M9BhlOR4DNmFvMIKzSp9V+eS0QPwgNE4k+cZwy4pzCoZxCoZtQlBVpDDGNVMdlGqhWPFxRTrIH1OWR0Iluil6aITLqmg/ZYWnKq0PuFPKEyvwloAzjIenSsJsRAWSjiNIIERwXREj4MfxJNvulWq7VBGuOFd4UjA37g3acE/ggcE9Etu5F7iHuE7Z5O7/G23DK9zXiHr8rnDfzwpRq+FRd8YSkIAEJDBLCOhhMUuwe1IJSEACEpCABCQw4wTmmqtx438M3uuAkvfeeSvCIVVGrMCT4pTzr7hhvvnmX+DAXbbZFMN/l3XWXe/9d96c9PVXX2AgrNVlgYUWXmSDfptvdffNw66aljKO1+rBOjgJNAwCISZE+CZEBbwh2M5nt/wnCbcxYhPqBqN0i1TxrkCsWD9VEgtTyH9AX8TuZz8r8JdOFaM5fePdgKG9JFUW4+EpUdFV52X9L1zpPED58VbmA8M854mwWNm2kUib0FB4IlS0wKSyZYFSGjAuwjPBnHB7fM+GIoI348RwTv4QrgnzwWOGT/avkf9EbMK7Bm8WBI6SVAmltWSqiBQIVLQnlBSiC/cK15VtXP+G7F2Rpp8reBghBnGN8WSBXQh1cYyfEpCABCQggXpBQMGiXlxGJyEBCUhAAhKQQEMksPGArf9Bvokrzz/7lBAqKuNh8c+9Djwcj4rLhpx+4itjR49cuPmii620Sus2tw674uK6wHPrHXfdq3HjJk1uG3bVJXVhvI5RAg2EQIgWGJvD6M1qeYQGDNKxOhyD9WupEtoJ4yshhPBWwEiPcZzvGLfZhwGcT4zrfMeYjcEfYQODNkZuzkHhnIR6wnuiqoVE0FEYT6xmj7BJIcjE/9PMFSN7YWEsjCubCwPD862pYvzfJFWM+SSgpuCVQH4O+kIMoP3Aqk6iCu04H9dkqVSZU3g4EMYLIYL5wgDhiSTQXLtY9U9YLzwmYMO1oy+8Krg2MGQb15jQYM+mSoJt8jJwHTknxneOC+8MOOUSrzfAvBVMO1c6Ljt/owkf5fR4uCPu7JcqIhJiHmHVKirQTe/TLxKQgAQkIIHaTkDBorZfIccnAQlIQAISkIAESiGw014HHDblu/9+e/8dNw2LQ/78488KGS9at23faZ/D//XvCS+9+PyVF5x1Cu3XWKtHLz5fGvnciNoOHe+SbXfefd+xLz73NB4htX28jk8CDYxANh8ChmcM8awMx0sCIza5KVqmGomEMVZjEA8Bgv9TMXzzc4tUCYdDXgMM5/TDPraxip++2B5JuNlGX5yHkEX0TZuqhm4qFnqH8RHeKLwTMLQzBkp2+wPpZ4z/EbqqVf6YTdMnwgSc6D/CMYVgEfkbOKZYgSliAnNF3Ij+ObaiuSg4FkacM8aONwdeLvClIrQgHjEO5so22pA3hDFwbtoyXrwsECO4phjUS1LlmnAM+2CGyMH1oA3HIdbgLYCoQx8cj3U+RK8GLVYkDoUFXhTBFZhYAAAgAElEQVSuBYJSeWG8inThJglIQAISkEDtJ6BgUfuvkSOUgAQkIAEJSEACfyOwdq8N+uINce0lQ8/88YcfMJblStIryhUs5p5nnnlPu/Ca4bQ79oDddvzj999zq1jXWKt7Lzw0xo16ntjktbr0HbDV9niXnHPi0QfX6oE6OAnUcwJp9Xtp5c+fd5u++pv/O3lOYVjH2IoBGzGCsFCswH8qVYzhEZ+fnzFkY8QmWTMr9zGUY7DFUI53Aob2yG9AuCHC2BFiClEgG7ooa8yf0auRNRBnQymFwZ/+s9vxoGCcWdED438IERjmEQla5OeK+BKlNLGC/TBgLMyt0LMDTrwHsl4dpc0bvuFJgZDAOGlL/7DkmiH24PVAjgm+My6SmnN8nJ+QXQhIvEtggchxb74fhKleqSLkTEwV7wo8LegLjwG2czycOF94z/zRkD0rEofpJeNlASPezwhGIXYZDjELy+8SkIAEJFAvCChY1IvL6CQkIAEJSEACEmhoBP655wGH/fbbr7/ecu3lF2bnjvjwZ0q9XRaPw044Y2iLlVq2Onyvnbb+dPJHJErNlc7duvd8983XJ/73m68J81Gry6Dd9zvku2+/+fqpR+6/u1YP1MFJoAETSAbnP5JowfMoGyYKIhipER8wjuOBwMp8DNwYvDF8T0gVUWOjVAkLRRgowiYhSrBKnxX8GLzJiUBIIgzsJOnG4wCDN4Zd2mCMxwjOvooUzp0VHyrSpqxj+H+7rP+5GSuJqcP7Iys+IMZg4GeuzDEKc0LkiWTXhedHhEBgQLDAcyErghQbK+ekP64Fn7BDrOAacW7GBleEihAz4M34YlwID4gX/Bwhrcgn8liqhC3i+sIVjxP6p1+u44v5MUY4L65/hBIr8z1WbCINYBtMyGPB7wKi0QopXBTs/0TUsEhAAhKQgATqCwH+8LBIQAISkIAEJCABCdQhAq3atOvQtXuv9R+7/+7bvvjsEwxT08sfqSQni1K9LHr36T9gyx122ePOm6694okH77kjGi60SPNFV2y56mpjXniWlc21uqzZo/cGLVuv3u6hu2+76ddff8HAZpGABGovgRAseC5RMdKzOp9n15hUWTFOPH4M2mx/IVVE076prpUqBn/CQb2XauRN+CB9xwiOMZ0wUwgXGNEjlBTHkxcB4zg1yl+el0WQVUSsKNeLrZxLgSiSLYWhqgj1hCEf4z1jJ+9HtkQIKESFYgVG8VwsS6xAGIAdTBhTCARsgyPnfyvVl1OFNWOhDbknGCMJz7leeF7wiZjEd9jTnmvHNeRack0jFBTXmmvOtefcbOeeiPsjK3ClzRYIZAQJeIVYlc21IigJSEACEpBAvSGgYFFvLqUTkYAEJCABCUigoRAYtMf+hzLXG6648NzCOec8LFIpxoIQSiecfdFV7739xutnn3jUQdlj8K7g55dGPltm/opFmi+2+D6HHXvytXc99vztT4yauP+RJ5w2WyrFztetR+8Njz39vMtmTyX2M4bDTzzzvFPOv/KGpZZZrkV516zH+n36nXXpsNtueeT5CZffcv+ThMHCu4J2d99y/dXltXe/BCRQKwjwTGJFPp94RhB6iNBJGN8xkGMcJ6k2BnFW22PER5RgNTkryElSzRJyEnezuhyx9elU8dLAeE6fz+WPj9wL9I2XAaGn6JdC+xktM/o/dKEo8mZ+QIRFwujPmJk/8+iaarHnK2Gf4DPdQy4zqXj+wxE22YK3CYICn/RRkipCBIIF50foiATm/Mx+vFPoC2+JELnjeISH21IlZwiVa8q14ppx7Rgjc6E914BrHLlGuD4cz73A9cveI+lHSykEECy472HPtZzR+1HQEpCABCQggVpHwJBQte6SOCAJSEACEpCABCRQOoHFl1x6mT6bDdyWZNNvvvYKYVP+Un5PikWx1ogGp55/xQ3krzhqn122+/mnHzFWTS8IFnhnjB/9AvHFi5b+W22/09GnDLl4jjlmn2PihLGjm803/wKD9zv06LcmTXz5sfvvwmg1vTRu3KTJKRdcecO88zZrdvYJRx74yy8//9ymfacuF1x3+wMLN18UA2IjPEGOO3jPfxY7GcLGyUMvu67L2j16vzDiiUc+/ujDD9bru+kWZ1027LYVVm7V+pWxo0e+88ZrGMUsEpBA7ScQq+YxhmOIJ1wTIYRYVR8ixfj0nZwWGOgJJ7RqqsTnZ4U/x5KnghXlGLn7p4pAgbE9ElB3Tt8RJGhPn/yvyycG3fBi4Ny14X/g4WkcCBUYn9dOlVBKjJEwWJROqeLJwFzJV8CzDjZRCNdEoQ0iByJOFLbBtdC7gmuACBFhp8JTBPGCMFJ84vEAP5jBGlbkAyFsVZdU8XJBhOA9A0v62jx/LsaEJwbXivcIbbiGeHzwrsKzgnmEeEHf4W1Df+Fhkb5ayiDA7xCeL/wOka8F0WpaCg2V9cIQoAQkIAEJSKBOE1CNr9OXz8FLQAISkIAEJNDQCGw/eK8D5pxzrrmKeVfAAtGhGJNd9zvsGMJI4Vnx7luTCJXyl9K52zq5/BXfT/muMFxJ7rh/7nXg4f8eevmwZ594+P6Nu7VZfvdt+vXeecCGGNoatW7bAUPhX8qG/QdsjTfGHTdefRliRctV27S9dPi9jyWRZfyhu+8wEC+Q5osvwWrbvxUEieEPPTM2NV9yy/W6tjlo8Lab0ebBu269kbBVeHTcfM1lFzS0a+98JVAPCIRRGmM3oilhjfCwIMTNsqliNMfQjTcFhnhCCeGRwDMGQzer8SMxNEZ2jsXozUpzDOP0xerzSali1CUcEUIH58JgjsGeEh4XfOecGH3xRoj9GPc5f5TqyqeAQR+xgvOvnurBqW6dKuIC40CEicJ4mAMeFxipETBeye8kf0HbVDFa02eMm938j58ThQsK4g+M6JP5lqSK4MO5aYPwMypVkp0jIHAsYZtgiRjB+GDJdkSRVVLlGkTyZ64L14hrxTXj2sGQa8l1oj3XmGvNdeLac10icfqMhtpKXTWYwr3RLdUWqVYkuXqDAeNEJSABCUigfhCoDatL6gdJZyEBCUhAAhKQgARmMoGmzZrNR/6JD955643nnnz0wWKnIyRUYYimjl3W6r7XIUef+PgDd99O7orCdgssuNDCK7dabfVbr7viomJ9cs6Djv33WZcNOf3Ey4eeflIc8/PPP2HgakTy78J22+y0+z5Tk/px9YXnnEZ+jPOuvfU+wk2R6JvxMc7PPpmMkfEvZYmllln2ilvvfzLpJt/uvvUmvdIHhq1cIZQVn7R74uF775zJuO1eAhKYOQTC+I8RPjzCMLojYGIAJwk3n4+kyv+rfKewH+M2xnba4ZVAOwz5GL/xMsCQThuM4qzqx/OrfaoY8DHKR2biyJnANoz+GH1zz7N8YX/Wa6Fo2Lt0DIJIRRN60zXj+kfmPHzl+YmnAs9Dwi4hRGDwhwNiwuRU8bxAXMDbIQrbEBBapJpdiIhgQ1v4Ml+M24gVcKePCMNEP7BCjMDTg+94qCB+kIsC8QKhAU8L+qE9fXI8ojdeMHh/0D/CAwxJpo0gUpIqYgUeG2ukipiB0MFxXLNgDXtzViQIFSnkscCTIhXEN+4LCh4tWXGtIl15jAQkIAEJSKBWE1CwqNWXx8FJQAISkIAEJCCB/ycwYLuddiUM05B/H3tYaXkqkoPF740yOSUWWGjhRU6/+JqbP/1k8n9OPmL/3Yvx7Nh17R6ICOOKhIPquk7P9Y45beilt1x7+YVZsYJ+yCfB50cfvP9utl+8Kdp17rrWFeedcTLCw2XD73386y8+/+zo/Xb9B0IFAsocc84552sprFS2XeMmc8899Oqb75236Xzz4cGRFSs4rsVKLQl/0Wj4VZec9/tvv2G4tEhAAnWPAAZqBABEh/ge+RQwbGMUZ7U9q/URDcalSlgoPLowzGKx3SJVDPt4AGDkx7CPoPF0qggY5FNAvOCZgcGdvjCmc94Ip8S5EQbmTpX/i/EuKxpSL20vrUR4pdiPgb6sPBnkasgWjP0IM1ulShgonqWIEIyDz8jrwZgRDWATHikwi++Mg2PoH0EAIQBxBCECAYJ588yMXBGcl8p52LdSqiEisK1l/nzwRri4N1We97TBUI4XBqIIOTYmpnp3/niu18h8v1wD2iPE/Cc/rsidkX7MXfvgXV0eLPTbEArXOgT/0sS0hsDBOUpAAhKQQD0loGBRTy+s05KABCQgAQlIoH4RmH2OOebYfvDeB3z91RefP3jnLTeUNrukB/yeUkxgrEK3mO20C666cZFFF1t8ly026o7HQ7F2nbqtsy7bC/NX4NFx4jmXXPP6y+PGnHPy0blE19mC8JBrN2ZkNoxJo4HJI4McGcNT2Kad9z7oiJVatW6zXd8enX7Je2Rs0G/AVgguL4x4/OFsf/sdcdwpq67evuNR+w7evuS9d1ilO73MNVfjxj3W69OPOdx183VX1q+r62wk0OAIIEhgaA3BAkEh8h9EXgaM2azwb50qx+NdgOE7knRzPHkvMMSzypznHgZ6nnN4PYShHu+Kt1NFIEX0WC9VRAo8NzgvRnS8twhXhBE+WxAFOIaCR0NhSGW8FaLgbYF3A+dDQGCszJF+Syt4JfTM7ETs4Jzh3RHhnfAgQVxhTsyX76yyp3K+SGTN+ZgXPyPA8P9+iBIIEvBG4CGkFCGdGD+86JMQTjzLEU7gjUdEhHSCK2JFJMrmO+zxcolzc924Riunyrjpg/ZwQSiBDf0Ez5xI0eSq3JgslSMQXo1cP+5fiwQkIAEJSKBeEVCwqFeX08lIQAISkIAEJFBfCfTu03/A0ssuv8IlZ59yHDkhSpsnHgwk2Gb/HgcddfzavTboe96pxx3xWhIdSmvTKXlYIBB889WXGJSml0OOO+3cRRZddPF9dhzQp5hHw3obb7rFh++/+/bkDz8gEWuuNElZvfsN3HZH8k2QIJxQVPvsOLDvV198hsGtEZ4VfTffavtxo55/JhsSarV2HdfYYbd9D37+qcceevS+O24pHOsG/TbfitBS11485IxpU6di9LJIQAJ1gEAySJdWcobqn3fL7cZzgN9rnm14FmB4xxiOMRajPgZ8DN0ICnhNYBznOTE2Vbwr8LaI4xAI8NRA9KQfnj2EMOKTczyTKgZ3hNoIIYVQgPEXIYOCFwffEUF4nkay6ggplT9s+gdzoX2Eh4qQVYXHFfuZMSC+4AlCYm1YYOBvkTmYvvnfPUQTOCFMwIhxcj44sJ3+ED0YE/MoSRWxAvEHwSGSaNM9gsL9+W0IHAggeE8EQ7ggGJFvg/45Htas7n8+32+f9Nkr1RAjuFa8S7h2nBfhJpt0fXoIQcUKLkGVCmIQQhPXE54h/lWpMxtJQAISkIAEahsBBYvadkUcjwQkIAEJSEACEihCYIfd9jkoOS38cNv1V15SFiCSbiMarN1z/T57HHTk8S8++9Rj119+wTmltZm3adNmq7Zp1/He2268NnvMKqu1bb/F9v/c7fKhZ5xU6O3Aca3btu9Esu0LTj/hqGy7jTbdYpsUtWrBO2685vKTh1x63dUXDTkdcSKO6d57o00Wbr7oYuefdvyR2Xb7HXnCqb8nVeSck44iCe3fyqA99j/k119/+QWvDW8QCUigXhHAmB2Jl8P4itEdg2xJqhjjEQoQLPAKWC1Vwh1hPCfBMx4BGNUJTYTYQWUbK/0RNBBUETDWTxWD/rOpYtAnTwP5FQhdhMEXwYOQTAgUiAYRKgmRgPMXelcwZiqGekQDvDyyIa7Sj7k+MS4XtmUfY8HgzDzwVuibHyfHRj/0TXv6jlwe8EAMYDvbGCs/046f+c646AMW5PzgZ+YQ+UE4J0IC4baYM+PEY27TVPGseDF/fJf8PjxUCKlFn3ipwIQx008kTH86fUfEQNhAKEHs4RpyTZkrbSPpul4VCUY1FFjDWcGiGmDahQQkIAEJ1B4CCha151o4EglIQAISkIAEJFCUAMIA4ZduHXbFxYV5HQob/PHnH380X2yxJU678Oqbvk0uE8cduMdOpeW7oG37zmuujddDYTioPQ8+6oRvv/7qyxuuuODcYoPaZZ9DjiLs0z233nBNdj8ix8TxL41KwsTG06ZN/f6qC88+Nbt/82133CVtnvLYA3eRDDdX2nZcY8211l1vo1tS0m88NgrPh/gCA0SV8NTwVpGABOoNgcKkyxjeMbATSigSYmP0jvBCeFhgqEVswBMArwba8J3wSBjJ2Y/RfVKqCBYtUsV7gVBIiBl4MCBaYPzHYB+eFhj/6QsjPMZ/PAQ4N/tDREhfc+GW2B4GY8aLFwaGefqmX8QGhAC24UGBWEDfkffig/x4yBcRDPBMYAycm3ngrYAYEgIDniEwCU8QhAPGhmcE5+VcCBGMDYGB/hgrnhKMlePwNMFDgnGQIwOxB7sAXhwlqb6ZKiIHgk8IPTBjP/0Fa8ZIP4Took9yVzA+xoxgwXeuYYgnIVbwaakigUzi7chfwrWOEFxV7NVmEpCABCQggdpFQMGidl0PRyMBCUhAAhKQgAT+RmCHXfc5EM+JG6+4aEh5eJJe8ceiiy+5FCLFPjsM6EPOi7LadFxz7R7snzDmRVbG5spSyyzXotdG/Ta/bMjpJ/6QVIfC9nhXkIdi2GXnn42oEftbrLzKqggrN1558dDtB+91wA79e3YhRFXsJ6RTj/X79Lv75mFX4S0S2wf+Y+fdmd9NV140tPBc5OE44OiTzmD7TSnZdnnzd78EJFBnCWQN2RjeMcRiIGc7zxEqggShnjDQIjhgJEeEQGDgWcTzDMM6Bne8B/h/d/lUEQTwHCB5N14DHIPHAdt5RtJHhFlCKIhQVMBEeKByDgQMjuO5yLgw+iMwYNhHOKAd2+ibc0doJs6H4T77/3d4ZHAORAhEDfriWIQO5hvngwPGf/YjViA+wCCSakeeCESEEE2y+Q1YgR8iDdtJTI5QEsfTz9Opwpd+4cE8YIigAUOuB6G1CCmFsRzBBbGIT65JiEUIN3BgTMw/8pWEYJE2WaqBANeA8F3cIybergagdiEBCUhAArWHgIJF7bkWjkQCEpCABCQgAQn8jcAizRdbfKPNBm474pH77578nxJCmJRZwpuCMFCjnhvxeHnHd+7WveeXn3/6ySep8zi238DtdmyUOkJYKGxPfoyjTx16yZTk6nHdJUPPzO4fmLwrfvvt11+7995w46Gn/uvwTyd/hNFweuk/cLtBc84511y333DNZbGxcZO5596w/xZbj3j0gXuKzW/bf+6+b6s27Tq8/NKoF95547VXy5uP+yUggTpNAKN2hAviE2MsYY0wlmNw52e8sCJfAsJnJKLGUI8IQMWQi6fBtvl2tKE9hn4MveE9gIhBAmsEA/rC8IuAwbNrpVTxYMBbAEGC/j9ONYQHPBgYB4b9CMOE2MEcOJ7zYfynz6j8zBw4H3PCqI8AQRvGRl8cG/kf6J9jEWM4HtGE4xhDrKrnnAgDiCiEt0JEgBmeFYwZIQFhgnPQF/vxUqE/cmAwbzwlWuTPz7GE3kIcuTVVnrv0z1gQiMIbhXPAj/HgYcHxXDPOCzPmieiSvZ7pR0s1EYA31wVxy7xO1QTVbiQgAQlIoHYQULCoHdfBUUhAAhKQgAQkIIGiBAbusMsec83VuPGwMvJQZBv+mhI9vDJ29MiLzjz52PKQNm7cpMnqHTp3feaxh+7LHtu7b/8BEyeMHV0s/BLjIYTT8YfstXM2PBVCRP8tt9+Jzw8/ePft+28fPqzw/JulcFCvjhvzYlZ46NR1rR5Nm803/yP33nFz4fHLLL/CSgccfXLOu+KOm665vLz5uF8CEqgXBLL5DTCqh6cB/7vyHaEAgz5GcYQFvAEIB0V4I0RdVvtjhGc/4gOhoxAa8A6gbwz27Me4j6EXQ3+ERMLIjjiAiIEoQHik0alGiCiOw8jP+UJ0YCyR8wJPCMYYIZsQLbKhrdiPIEAlBwSfjIdxIHKEaMJ2+qcyDgzT1PCAYMzMBdECAYH5Rbgn9jHunvm+w6BNX7RnDIgizAmWCA+IOIyT7STYJqwT+T9g+EKqE1JF5KBNhJTCswLPC7xJGBv9MIbI7ZETn0ysnShUcyEsVL5MmfDRlPD2qeaz2J0EJCABCUhg1hFQsJh17D2zBCQgAQlIQAISKJMAuSW22nGXPfEuIC9ERXCdfMR+u3/79ddf4ulQ3vGrte+4BqLFy2NHYZDKFcSD5NHQ8ZqLzz29sP1Kq7Ruc/Cxp5w98pknHy0UJHputMlmhHxK6Sm+O/Xog/cubLtau45rrNxqtdVPPmL/3bP7unbvtT5jffGZJx7NbicZ+JCrht89z7zzNv3vN19/9fgD99xe3nzcLwEJ1D0CyaBdWvnz591yuxAAMH5HngiebYQlwrMghAkM/mzHsE7OCv7P7ZYqhv/XU8VY3yvfDx4AEdYIDwGM8hjiS1LF8I7xH/GA4yKfBZ+ID5H8OkIdMSYMxmxHpKAf9hHeiTGwjbEhBITgws+IA3g1IHQgGiC20JbzRAJtjmc/XhL0Q2UbLBgzfXJejmFszDFyYSAkMHf4wIU5YeXGG4ISP9MeFuS4aJM/Px4rMKM9YaN49zBPxstYEXU4P31zDRgzQgUc2DfdS6auixVN5p5nnngH5blV+WOFlVu1/vijDz/45eefYFRtJYkX5gSpNpp2JAEJSEACtYUAf1xYJCABCUhAAhKQgARqIYHeffoPWGyJpZYmV0RFh/fZx5P/QzLsihzfLrk3cByCSBy/5NLLLkfYp08++v8QUeybb/4FFhx69c33TJs6ZcpxB+2xU2H/A7YdNJhtF55x0jGEmPrb/u0GDWZcj93//8m2OYZwT4SOmjZ16vSQFrPPMcccp114zfBll1+RkCyNHrnvzluq28hTET4eIwEJzFoCGLzzRu8wxGOcxzAeHgUY8THWYzAvSRWDfHhAsA+viodSfTBVBAiM/ISKQjAgTBRiCIZ8jP2EY5qcKu0w1rM/2rRI30naHR4OHB95NSL8U+SbQHDgeYYxH7EADwfOy3ORcbIdj4bOqa6dKoZ/jM5sY56EoeL8tOX8zDkSbXNO/odHaMCzgn6ZMx4hiAsdUm2Rb8848DgJMQVmzJG+mDN9MUdYwIS+OB+sYAY7WOBNAlPOU5JqJPhmH9/pl2sSIaHiWmU9ZdLuulcuHHb7g+deceOdMzrylqu2aXvrYy+83GGNNbneFglIQAISkIAEyiGgh4W3iAQkIAEJSEACEqilBLYetOveH77/7tvPPP7XkE3VNdx2nbp0I/n1W5Mmkog2V/Dq4LP5Ykuw4jdXklax0EXX3/kQHhS7bb1Jr2+++pKQItMLosraPdfv88bEV8bfcePV0/NTxAHkqei7+dbbj3ru6SemJReMbFtWry6w0MKLcN7ff/vtNzw+Th566XXrbtC3/8inn3hknZQP4/EH7ta7orouuv1IoA4SQLRI3hYY9TGKR4goVv0jFvBMCeECUQBDOc8vnlMkmMbQjuEer4fIcYExnrBJ7F8tVQzueBoQJorCfgz3bFsiVYz8hDxiO+GSuqaKMIyBPxJX03/7/FgYZ3hIRPJwzoGHQuR1QFDAewLPCgrzQThgToSJoiCCIFAwP9oTnmqpVBEeOD/CA3NiO/NtmyoCCHN7Or+tf/oknBMFkQORgX4npYp4smq+D/gyB+a5YqqMm/2Ro4LxwoHzRqJnxh/zCU+YOi9UACo5Gy5Ajic8AAnLmKItck2rVA485uQz6ePHH6bB0CIBCUhAAhKQQDkEFCy8RSQgAQlIQAISkEAtJLD8iiuv0nWdnuudeszBe0ci7eoeZpuUv2LSq+PHIhRE3yn9xJsYaP4xeK8DPip5791kY2m858FHnzD33HPPs8e2/dd/6/VXp4sb0abfltsNYoynHHXAnn+kUjhOPEXw0Hj+qUcxAP6llKTzdeyyVvdTzrviejw9ttxh5z1atl693QVnnHj0CiutgiGtUcl7b2N8s0hAAg2YQF60CK8GSOARgOE88kdE3ge8DchtEYmseb6FFwbGfhJuRx4HvBow9iNEdMq3QbQg9wWGewQGxAEED7wrCJeEUZ+CWIBYghjA/9WIAYyF89IWzwq+R/gnjmGMjIXzMi720z+VtoRdYo54NCBaIA6EqBG5MRANmHt4NiBkEMIp5sjc6I++GS8/8yzFe4T8E+TOwHCOIMGYqDBBnAjvCYQTtiN+RJ4MxBnGwJgQJeifyvii1Auxgsm0T94QeBsioq/atn2nioZlzLDIfe3Qpds6CO98n/r9XwX7wmP9WQISkIAEJCCB/xFQsPBOkIAEJCABCUhAArWQACLAF5998nGx5NXVMVxyRCyx1DLL3nfbjddm+yP00g1XXDRkl30OPvL0i64ZjgDx+AN33XbWCUceWOhZEe06dV27xxnHH77/pFcnkKT1b6V3334D8Kx4+J7b/5ZY++6bh13Vb+C2O/bdfKvtqcz5uIP3/OcDd9x8/bGnn3cZq1qzyb2rY+72IQEJ1E0C2ZwI+fwWIbZiwOc7gkCIGHzHgI6ogNcCRn0M+HgkcHx4MSAssC08KOgnVtNH+CSAYazvnioCQAgLhH6KkEx4QURuCdohAFDDoI8YEOIE40IAoSBoICZwXsZASCj6YR4chxDCefjOWBkb4gEiCx4inCvCVSFIZPNd0P87qSLg8L8/CbVJUh7JxtkPF/piGx4qCBkIGoyDNiFQMI/I3RHCRL1Nqo2QDhwK3ohVFSz2O+L4U6OfH9KLML77KQEJSEACEpBA6QT4Q80iAQlIQAISkIAEJFDLCBDzemrKF0F+h5k1tB7r9+n3wojHHy7mFbHKam3bp6hQS7/75qSJn30yGeNclcuCCy/SnFWqiBHFOiGkVKs2bTt8+flnn7z/9puTfvnl55yBr20yEqWmiz7z+MP3V/nkNpSABOo1gSRcZP+njRwNzBnBIhJdIyV5JGcAACAASURBVFggLCAKRFg6vA7wEMAIj2DRIlXEAJJ2h7cB4aIQBfA0IMwU+Rx4jkWYJ5Jbr5Jvx/nwRuA8eGkgOCCQhDdF5KbAaM35OC9jj8TcjDHaMA9CReEtwn4EDcaAUEA7vCneSpX3AyGqOJ7E2TyrES0YA3Mg7BNhrZgDOYFoV5IqY4jxhgcbHiPhVRHhn+AVOZEQbJh3FMSKeluuvvORZ5drseLKhER8+rGH7jtyn523rexk11p3vY0uuemeR6Nd99ZLL1AYFrGyfXq8BCQgAQlIoCEQULBoCFfZOUpAAhKQgAQkIAEJSEACEqiHBPKeFsyM/22jYtiP0El8x1AfSaox7vOdz/CmQCjA8wAjPwIBIgMVkQFPCMQDRIhs8m/CRJHkmrwRCAoUwkVx3t6p4jmBxwRCAAXhgPZ4R9An5+JnRAmO5TjGjycGhf14gVBHpIpgQD4NCmOZmCoh+sg3wfxi7oyFseMJgmDC2KnMEeHig1Qj5wcCBSIEIjGfjIfvEWaLnzkvff8tmXZ9FSwQ2J97Y/J3zz/12EOLLr7kUosm9X7jbqshTlWqXH/vky+2ad+py3vvvDlp5Varrd55+QXnmFkhHis1MA+WgAQkIAEJ1HIChoSq5RfI4UlAAhKQgAQkIAEJSEACEpBAuQTCoB6L8hAj4jtGeGqEWMJgn83hwP/FeB3gfcF2RAc8EPA0wLMBMaEkVfJFICCwnZ8RCugTrwbEDc6JBwaeGJyPPiNfBCIAP3MuBAXOQYmcGPRByCd+pt9IMI7A8W6qeFAQsim8Nt7IjwHxBe8MRA/aUxgz5428HpwXTwk8QEKk4GfGi3CDmMF4g1fkIpoe+intqzf5KfKMSv1AZEC0eP2V8S8hVmy3y577I1x8+fmn8K9QIW8FXoIP3X3bTc1TJz8u+8M0xYoKofMgCUhAAhKQgDksvAckIAEJSEACEpCABCQgAQlIoG4SKLLKP2tYz31PXhjZbVnxAgM+wgGfkfsCzwaM+Gyj4PEQ+xAzwvsAoYDtJKjGk4KCcIBQ8GKqJM5GMAhPjpL0nb7xdkCEQKBAIMDbArEDEQNvi2wbRAj6p89Ioo2gwTg4N2NAZKFf+uNciB2RKwHvCAQOjo8k5XynL/bxWShSpE3/41VfPSiYW1mlU7d11mX/axPGjl508SVSovY9G63eoXPXEY8+cE95bWP/ngcffQICxTUXnXv68WddeOW0FOKxom09TgISkIAEJNDQCehh0dDvAOcvAQlIQAISkIAEJCABCUigHhMoSNad8x7Ib/sjiRkR8igM+ZHAG6M9ogU/47FAQdxglX2IGRihEUDwVCD3BYIBnguIDwgF7F8kVcJB8TN9IjRQ+F88RATEBvYTxgnxApEkwkkhWnAsHhWRQyJEFz5py5zoFw8QSnibZAUJtjFOtk1Plp3JAdJgPCjyjEr96NR17R7kdnr9lXEvLdx8MXKENMLroqKCRff1Ntqkbcc11nzyoXvvfO/tN16fZ955m06basLt8ri7XwISkIAEJBAEFCy8FyQgAQlIQAISkIAEJCABCUigQRDIihf5CRfmZpgeBikdG6GR8NJAXIjE05EjA5EA8YLjqPx/jWhByCnEBzwpEB7IK4GQwXb2I4BEzgg8IkiSHV4TeFjEfvqnX4QIRAwEB84X56RNNsfEHwXiDFPM5q38vXD+RXg0iPugtEnOPsccc7Rfo9s677016TVEBup3337zNR4WFQUT3hVXnH/Wv2kzz7xNm34/ZQpeMBYJSEACEpCABCpAQMGiApA8RAISkIAEJCABCUhAAhKQgATqH4FM2KOiHgZ5oSLrsRDHhXiRS0iN4T8diwcGNYSMCCHFzxzPJ/sRHviZgpcEYgbCBNv5HiIEgkdsR2z4PT+e7DnjouS25ZOQx3726TlRids25cZu37RZs/leGTeGsF658trL48a069x1rdlSKS8PBd4ViBt4V7w9aeIrtJ97nnnm/aIS+S8qMVwPlYAEJCABCdRLAgoW9fKyOikJSEACEpCABCQgAQlIQAISmFECBR4IhcZ/BILIk8GpIi9EhG7KCQepIkTwyfYIM8VnbCMvRvQdx9KW7bkS48h/Th9HKYKLIkUVL3ynNf+Xv+KVcaNHRheIFyTRXm6FlVp++P67b5fVNd4VhJO6bMjpJ8Zxc6eYUD/98AN5SCwSkIAEJCABCVSAgIJFBSB5iAQkIAEJSEACEpCABCQgAQlIoJBAeUm/8x4PWQEhvCcQJighakTX2ZBUAq9hAh1T/gpO+fJLo16IU08cP2YU38ljUZZggaiBd8Wj999567sppFS0x8Pixx+mKVjU8LX0dBKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCCBOkvgqZff/+KJCe9+lp1A02bzzT/uw//+fsRJZ51f1sSuv++pUeNKvv2txUotW8Vxs6cy4aMpf/576OXD6iwUBy4BCUhAAhKoYQK4oVokIAEJSEACEpCABCQgAQlIQAISkECDJbDCyq1aL7RI80Wz3hXAmDb1+ynvv/PmpLISb+Nd0bbjGms+cNctN5S8985bAbHJ3HOTRL3RTz/+QCL1ai9zzDnnnE2SC0dFO+ZY5rHSKq3bVLSNx0lAAhKQgARqmoCCRU0T93wSkIAEJCABCUhAAhKQgAQkIAEJ1CoCndaMcFAvPl84sFdTHotWbdp2QCAoNmhyV/z226+/Xj7k9JOy+0NM+DHFhKroZFdOmb/xyLjq9oee3qDfgK3KanfcmRdcceVtD46IYxAizrp02G23PvrCyyecfdFVeIfEvrXWXW+jR196c/IN948YfceTo1+77fEXXyUvR0XH5XESkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQnUAIFTzr/yBsI3kaui8HSbb7PjLuxr3bZ9p8J9Pdbv0499x5w25JLCfYsvufQy7NvnsGNPrsgUthq0615j3v/qZ9pQn5zw3udltUN0IBQVx/TccJPNRr/35U+j3vn8hwdGTnx//H+++wOvD/aRR+OJ8e98Sn97HXL0iUOuGn43/V9y0z2PVmRcHiMBCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkEANEXjoxddLRr712dRiXhTkpcDAv/Wg3fbODme2VPBmQCRovtgSSxYOFQ8G2u26/2HHlDeNXfY95CiOvf+FV9/rvt5Gm2y06cBt+PnUC666EcGhsP0CCy28CLk19j/yhNPadurS7aUPvv5l+EPPjVtqmeVacCzhraLNen033YK+Nh6w9T9iGyLK7gceeVx543K/BCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACNUQgPCEuG37v48VOiTDx9MQPvy5Mnt138622Rwg46Nh/n1WsXcvWq7dj/6A99j+0rKlEP3hLLLDgQgtz7Jo9em9AWzwlFlx4keaF7QkXxX7EjQdffO2Dmx585qWmzZrNV+w8g3bf7xCO7dhlre41hNTTSEACEpCABKpMoGj8xSr3ZkMJSEACEpCABCQgAQlIQAISkIAEJFCHCHTIG/LHjR75bLFh/5nKxPEvjcKTIfbjibH3oceeRFLuay8eckaxdk2aNJmb7b/8/PNPpeFo3bZD5xPPufjqd9+a9Nq+O27R9/sp3/2XYzfdcvud+Jz06oSx//3m668K23fu1r3nTyk5xto9N+jTNCWrGDywT49pU6d+X+w83/3322/YvsTSyyzX6KU6dGEcqgQkIAEJNEgCJt1ukJfdSUtAAhKQgAQkIAEJSEACEpCABCQAgQ5duq3D54QxI58rjQiJt5dfceVVCMXEMVvtMHhPQj5df/mF54YgUNi2cZO5c4JF0iuKChbzJ3eKoVfffM8vv/zy8wE7b90/xIoU1WlFvC5oO+b5p58sNibyU0z9/rvvttlpt32GnvKvwz//9OPJpY19zAvPPIno0mP9vv284hKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCdRSAjc//Nx4kl03SckiShti13V6rkdYpXU36Nu/2XzzLzDilQ++fPrVkq9KC8NEP2utu95GtNlki212KNYvibrZv2H/LbbO7j9pyKXXRuLtXhv127yw7eypkDeDY0i8Tciq8tCSYJs22dwW5bVxvwQkIAEJSGBWENDDYlZQ95wSkIAEJCABCUhAAhKQgAQkIAEJzHIC88w7b9NVUq6JSa9MGPtzirFU2oBee3nsmD9SIXwUSbTJK3HtJUPPLC0ME/38v4fF30NCEQpqy+Sl8cAdN1//+AN33x7nXbnVaqv3H7jdIMI9se3N114ZXzimZVusuHKIK9dcdO7peE+UB/K6S887izb/2HXvA8s71v0SkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQnUMIEua6/bG0+FA4468fTyTo03w73PTnh79Htf/vT4uLc/Kcsjg7422nTgNuGVke0bj4gb7h8x+sW3P5/WfLEllszuu3T4vY/hCUGoqOcmTc7lsygs62+82UD6fWLCu5+RS6O8ccf+q+94+JlnX//o23lT0ouKtvE4CUhAAhKQQE0T0MOipol7PglIQAISkIAEJCABCUhAAhKQgARqBYFIpD1u9AtFE25nB0keC/JWNG7cpMnVF55zWlkeGbRLh+VyWPz266+/ZvvpsX6ffqt36Nz1xqsuGvrVF599Gvt69+k/oFuP3hvecOVFQxAyPnjnrTeKQVp51TZt2f7QXbfe+Ptvv/1WUZCMOUWzWnDzbQcNrmgbj5OABCQgAQnUNAEFi5om7vkkIAEJSEACEpCABCQgAQlIQAISqBUE2nXq0o1QT6+MHT2yvAG9NmHsaI757JPJH901fNiV5R2PsMExSVP4i2AxaI/9DyXk0/WXXXBO9EGIqWPPOO+yyf8peX/Ypeef3XLV1dp+/NGHHxQ7R6s2bTuw/dH77ry1vDFk94985slH33/nzUkDFCwqg81jJSABCUighgkoWNQwcE8nAQlIQAISkIAEJCABCUhAAhKQQO0ggKfD25MmvjL1+ynflTeiCS+9+DzHXHrOqcf/8svPP5d3/FxzNW7MMUmwmO4FseQyyy7fuVv3no89cNdt6ZTTQz7964zzL19gwYUWPnrfXbZvvtjiSxBu6pOPPiwpdo5V27Tv+PmnH09+/ZXxL5U3hsL95MxYZbW27RdfcullKtvW4yUgAQlIQAI1QUDBoiYoew4JSEACEpCABCQgAQlIQAISkIAEahUBjPaLLLr4EuNHjyw3HBQD//D9d9/eolfnVe+7/abrKjKROeacI5df4vcUtymO7967zybksBjxyAP3xLbdDzzyOPJSXHTmyce+9vK4MYSdYt9nn3z8UeF5UkSnhRA9Rj79xCMVGUPhMS+/NOoFtq2cPDiq0t42EpCABCQggZlNQMFiZhO2fwlIQAISkIAEJCABCUhAAhKQgARqHYE27Tt1YVDjx4x8rqKDK3nvnbcqeuwcKSM2x2ZzWKzWvuMabJuYDy+18YCt/7H3ocec9OTD9911/eX/CxG1eFIk+Jz6/Xd/8/po1aZdLhzUSyOfHVHeOAhJhQdJ9rjZZp89ZwcqDFNVXl/ul4AEJCABCdQUAQWLmiLteSQgAQlIQAISkIAEJCABCUhAAhKoNQRat+vQmcFMqIRgUZnB40nB8b8nF4tot1DKVcH3/3779Vf9t9p+p1POu+L6N197Zfy/Dtx90J+psK9xk8a53Bc/TJv6feH5WrZu045tb0x8eVx5Y9lyx132vP6+p0Z1Xafnerl+k4AxeN9Djvrxhx+mpXwcY8pr734JSEACEpDArCCQU/stEpCABCQgAQlIQAISkIAEJCABCUigIRFotVq7DnhMfPPVl1/MzHknweL36P/Lzz79hO93PjnmdUI/fVTy/rv777RVP5JwxzGvjn9pFN8P/tep57z39puTJn/4wXuxj/wT3337zdeEpypvzM8/9dhDhx532rlnXnLdrXhkrNa+0xpLL7v8CmefeORBSQuZUl5790tAAhKQgARmBQE9LGYFdc8pAQlIQAISkIAEJCABCUhAAhKQwCwlsELLVq1HPTfi8Zk1CDwZ/kglGxLqxqsuHvr+O29Oar7YEks++dC9dw7esu+6X3/1xefZMUxMgsXVF55z2tLLLb/CSqu0bpPd13LVNm2fSO3CG6OssSOGnHj4vruSwHvD/lts/cPU778/fK+dth5+9aXnz6w5268EJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAKVJNBpzXXWbdpsvvkr2azCh6euF1hjrR69Ktyg4MCUAuNvUTE22WKbHUi8XZk+55qrceMFUiyqyrTxWAlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABIy7K2AAAAI9JREFUCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhAAhKQgAQkIAEJSEACEpCABCQgAQlIQAISkIAEJCABCUhgVhH4PwbQv9cuSoUuAAAAAElFTkSuQmCC"}],"notes":"","preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nO2deXwc1ZXvv1XV+95q7bI2S7K8G68YYzaDCVsgEAiQCeRlJpm8mSxAVjJbkmHyknl5WYaEEMgykwUSJgEenyQME8hCIMYGY7zgVba1WUtr6ZbUrd676v1xu1syeGmwNvvd7+dTH0nVt27faql+Oufcc+5VTCbTLsMwWpBIJJKToCjKYUXTtFg2m7XP9mAkEsncRdO0uDrbg5BIJGcHUiwkEklRSLGQSCRFIcVCIpEUhRQLiURSFFIsJBJJUUixkEgkRSHFQiKRFIUUC4lEUhRSLCQSSVFIsZBIJEUhxUIikRSFFAuJRFIUUiwkEklRSLGQSCRFIcVCIpEUhRQLiURSFFIsJBJJUUixkEgkRSHFQiKRFIUUi7MKhZZFS2Z7EJL/TzHN9gAkk1GY19jC0vNW09jcTFl5BVarjWwmzWh4GJu3nKZKJ3/9/jvIZPXZHmwBs93FrXd+kL3bfs9rO3fP9nAk04TcCmAOUFZdzw233cmmK69mdLCHXTte4WjbQQaDQeLxGIYBl7zzvaxfuYCuvhCtrS089dOH+M9HH0U3Znv0cMc99+FTRli36To+8p53MBZLzfaQJFOMpmlxNE2LAYY8Zv7wlVUbn/7yA8Yjv3rWuPn29xoej+uE7SwOn/HIMy8alWV+AzDsbp9x1xfvN+778pcMZQ7cx0OPP2c4zKrxkS98y9iwdvmsj0ceU39omhaTMYtZ4pLrbuO7P3mMA1uf4Y4bruSXP3uUsbHoCdtef8ff8Mdffp/+wTAA8cgI//b5uzBKWll93sKZHPabUK1ebEaEWFpnLDSCz++f1fFIpg8Zs5hxFN5/zxdYt6yBj9x+HcPh0VO3Ntm4/p1X8pFb3vGGVwy2vvgnWhcuY/vOA9M33NPgLiknGh4AwGy3kk6lZ20skulFWhYzzJ33/DML5zm5+68/cFqhAFi76Xp2P/8rIvE3xwEqKqsIhQenY5hF4/T6iYyI+ygrL2doaGBWxyOZPqRYzCAXXns75y+t4Z8+8xnSmeJmM6664SZ+88RjbzpfVtvCFZes48UXtkz1MN8STqedWFy4T/UNtXS0d83qeCTTh3RDZghXSTV/+5EPc9dfvJN0kdOeZoefBTVu9h/pKZyzOT1svv493HL7bXzl3o8QmeWZB6vFTjqZwOIqxamPER6XMyHnKlIsZoj3/s0neeJ7X2UoHCmqfaCmiS989X6q65r44RP/ja5nAY2WxUtp2/ki97z/3UW5MdONyWRFz2RZfdFmtr/w29kejmQakWIxA6hmJ5deuIoP/Ouni75mbLif0ooqHv76lxgOjxEaDDIyOsb8hcu4cNM7+N7jz/CDr9/Hb3799DSO/HiqGhexpLma5579XeGcZjaRSWW4+oYb+cmX7wLghjv+lt79W3hl+84ZG5tk+pFiMQM0Ll3DkZ1/JllknAKgdeVG+vdv4ec//clx548c3MezTz1GRW0T//S1B/F6nDz66C+Oa6OqGiaTRio14RI4PAGuuHIzTz/5GJmscdL3tTscxGOxE762ZPVGrrlo8XFioZo0fDUL8GljtHX2Ud6wlBtuuomBw/WnFAun2wt6hvHx8Te9pqoa/pIA4eFBdGNirC5vgIoyP0cOHz5pv5LpQwY4Z4Cqqlp6u9qLbm+yubj7s/fyna995aRtgt1H+PSH/oIbPnA3DovQ/NbzLuDjn/4s//LQY/z4qd/SUFuZa61w7/9+kJve9yHWr10BisYnvvQdfvnsizQ31BT69JTV8dAjj6EAvuoWPvO5e497T0VVqWloQpl0TtVUNl13I48+fD8ATrcLj6+EdZtv4ok/bOf22245/t6sDj731e9x/w8f4cHHfsOtt9503OurLr6aH/3q93zxG9/lP554Go/DDEB5XSvfffRx7v7iN3jPzTcU/VlKpg4pFjPAeCyCw+0urrGi8on7/o0XnniYtvZjp2waGx3kcFeIylIP3vI6/v4LX+CJn/2M+go/3//+T7jq2usAaFlzCV5jiD++8BJWm5Ub/+oTmCPt/OiRx1m5ek2hv6tuvoPf/9+fYwDlNbW4XM5J76Zy7Q3vIpzQ2HTJ+omzmsq+rb/lpVdETUj7nq1859sP8MuHv8on7/oES1ecd9yYP3zvv9Kz63f81S3X8cGbr+HZZ/9YeK2iYRH3fOIu7rnjej56x7v57Mc+TCQm8jZuvOPDPPbAv/Dgtx9g0TLRp2ZxcNGmTcV9rpIzRorFDHDgta2cd+FmzJpyynaqZuauL96PafQIP/7xz07br8nqoqHGR3B4jIvecSO//cUPOHasi92HurjogtV4fV7c/nLu/vTn+PF3v43bF0C1Bbjx2sv45te+jtPpJBYXAVez3cPtd97Jjm1iKrasvJrxyEjhvRauuwwl0snnP/tZbvvgRwvnz19/Mdu3TkzfqiYbt77vL/jvp39N1bx59PdOCF794nVct3kNjzzycwA+/+1HKfWYC69/8BP/wG9+9hBDoVGaVl7MXR//CAbg9FfyrpvfzcBgiPd/6MM891+/AuDKmz/AquWLT/s5SaYGKRYzQHw0yDO/f4VPfe5zmLQTf+Q18xfxtf94HD10iK986X9hsdlO2afd5ePv/s+DPPfYw4wnM4CBqggx+ubn76a8cTEXXvNevvnQD3ji4S/z6q59lJaWcdMdH+In93+JZDqLxWzFyGYBhb/5uy/jsiq5WReFy6++jpr6JgCsTi/3fPZeHvzaVwh27MVTXg/AorWX8Y6rL8cgH1dQ+KtP38fePz7OkY5e7E4nsXgcAIvdzb3//BXio2GyBpRUN7F+/TqaFiwC4PzNN3PlFZcwPjYGKNx4+x1kM1kAPvjJz9PXfoB/+ub32fbr/+DPW3cQqJ7P7be9ix/94Idv+/cieWvIqtMZQlE17vz4P3DZxefzu988xaGDB8hkdKrr53PBpZupDLh56Gv3sW3bdkDhi995lAqvme0vvciRtkOMhMOoqkagopqlq9axYsVynvjRAzz15FMAeMpqeeDff8wTP/keNm8lGzes5J4Pvp/UpKDq13/+HJWWCO+76UZ0YPnGa7jnrg/TNzxOcqCNZ7fs5S//x20EQzEiPfupXnYxPfu307x8Hb/71S+49qZbONTWgcc0ztPPvcRtt9/Kfz/7B0qtcb7//R/z15/9Eo2lJv7+U58kk9UprW3lWw89yOOP/pQrrr+V3/3nd1m2+b2khztpWrKSJx/5d95z51+y49UdLF7YxLe+8U3u/cK/MDQcRlEMBo7s5MlntvKx//k+7vnY3Xzz33/OS799kkhC550338q//ePH2L5DlsTPBJqmxaVYzDAlFTVctOlK5jc3Y9JU+o518uqWP3Fg/z6MN0xSlFXXsXLtehrmN+P1+dCzaYK93ezbuZ3dr+1405oW/vIaLrvyKuJjQ/z+madJvqFOo655McmxQYIDEynircvXYFHS7Nm1C4D5C5fjsirs2bULi8PNqnXr6Ty0h97efs7bcDk3vuc23C4He1/dwmM/+gGrr7yVazdvwFvRyM7nn+LhB75DdlLdfEPrcs6/YD27tz3P/v0HMVlsrFy7nq7DewkGB6msa6KhroYd27aQSmdweUtwOaz465fw/vfeRN2CFXzug++m81g/dpePTVddh82i8uJzTxMcGJri347kZMgSdXmc8XHpje83Xj4SNC6+cO2U9rtkw5XG1sP9xjVXXT7r9ygPWaIumQoUheef+y8+cNe9mNRTB3DfChdeeiUv/PpRnn7md6dvLJkRpFhIzggFOLD9j+w40M/VV18xJX0uWX8l77rhGsKh4SnpTzI1SLGQnBEGgGHw8x8+yDvfc8eZd6ia+OinPsOD3/hXVFU78/4kU4YUC8kZYRgGiqIw2PE6qq8ej/3MKghWbLyK8JFXaGvvOX1jyYwixUJyRmSzWZScBXC0/Rj1ddVn1N87b3kvT/7sx5hNJrIZWe4+l5BiITkjkvEkDpuYeY+Nj+Jwe952X6rFyZKWal7bvR+Hy0s8Wlw5v2RmkGIhOSOGBvoor6oCIFBaycjw2w9KVs1fQvDwbjI6lFVUMtDfP1XDlEwBUiwkZ0T3oT3UL13PgqWraKxycqSz7233FaiopL9HxCoWLl1O24G9UzVMyRQgxUJyRmTio3zvoe/z4Y/fzVf/4R7ewpIdb2IsHKKiuoZAdSMrF9exa8/BqRuo5IyR6d6SuYOq8akvfYulrY088OW/45VXXpvtEUlyyNoQiURSFJqmxaUbIpFIikKKhUQiKQopFhKJpCikWEgkkqKQYiGRSIpCioVEIikKKRYSiaQoVMMwpGBIJJJTYhiGphqGMXVroZ2DVNfWsWDxstkehkQyqxiGoUir4jQMDwzQe6yL1iUzLxiKInVcMneQYnESGptbURSFRcvOIzo2it3uPP1FOdweLzW19Sd9vX5+CxbryTcRam5dfNzXYvGVBCivPH7xmZaFS7Ce4r2A01pOl18zsbfo5utuLGosi5evLKqd5OxBisVJMJnNqJqGZhLLxKVSSfyBspO2n/xa1bxahgaCACdcR9IfCJBKJk7Yj6qq5Hf4UjUNq82G3VGcUFXV1DI8OFD4ubl1MQPBPswWCw6n66TXWSyWU/ZbUlqGw+nCHyjF6y8paiyScw9NUZR/BOTKqG/AZrORTiVZd+El7Nv9GuWVNaRTSUxmM15fCeO5VZwqa+bhcLmwmMUDV1ZZhcvtwWazYRgGF13+Do62TZRaz6tvpKKqhtDQIOVV1WgmE5XVNYyEQwA0tS6mel4tLreHxuZWfP4APV3tVFTXUFFVg68kQDKRoKKymrKKShwuN5l0mpraeqw2G8E+sR6Ew+li1foLOdbRjsfnx2KxYjZbqJpXy0h+1WxFoXnhErz+EtLpFFabDZvdQUlpGZGxUYDCaza7nZraBgb6ehkM9tOyaCmpZJKyiipi0QjLVq5loL+XhUtXkE6lKC2vIBYbx+X24nS5sVptlJZXMDY6sX+q5OxBURRdisVJ0A2DqppanC43/b3HcHu9mC1mGua3kMmkCQ2JXb2aWhfRcfgQVfNqqWtswjAM5rcsRFFVRsNhQkODRHIPSE1dA4Zh4PX5CZSVoygKK9dt4LWXXyKbzbJ4+Uo8Xh/bXvwjg8EgJrOJRDxGNpNh1fqNlARKyWazuDxe/KWl1DU0kc1mqKqpRdM0dF1naECsLpVOpzCbzYxHI2iqxqJl51E/v5lDe/eQzFk1S1euIR4bR9d16hqbxPus20AmnS6IzoLFS9m/ZydLlq+kr6cbVVWpqKrB6XJRWT2PsopKxkZHcbndeP0lBPt6mL9gEdlshkCgjJq6BjLpNKvWb8AwDPqOdc3Cb1NypiiKoks35CSkkgmWrFjF0bYDLFu5hsFgH9FIBBQ4fHB/oV2wt4f6+S3EYzFsdgdt+18n2NdDIh7DVxJgsL+30LaktAx/oJTe7k5cbg8H9+6mu+MoqVQSgH27X2NsdARd1/H4fIyNhMlkMjS2LKC97SAdR9rIZjPMq2sglUyyb/drjEcjuL0+9r++67jxq6pKJpOmJFBGoLyCgWAfA/29x/1nV1BoWrCIRDzG8ECQZCLB4YP7MCbto6igkEmnCQ0P0XH4EAC+khL27NiOryTA0ECQyGgYRVVxezxERkcwWywc6zhKMpkgmYgzEg7R291FJnP8doqSswtpWZwEQ9dJJZN0tx9FUVTi8RjJRAKHw8HYyEjhD7+xpZWBvl7S6RSqqpJKJQkNDZKIx4iPj+P2+ojmTHoMA78/QMeRQ5jMZtJpYaEkE/HC+5pMJsajEcxmM2OjIzgcTsKhENHRUYYGg4xHI4SHBhkdCZNIxBns78/1lcLj9TEYFJZFRfU8YtEo0cgYChAeHmIkFCIeGy+8l93hwDAMjrYdpLyymvDwID1dHRiGXnCzMpkM8dg4AznRMwydeGwck8nMsa4OEvEYNrudbDZLIh7H6fYw0N+LruuEhgbx+v2MjYbpaj9CJp0mNh6dgd+eZKpRFEVXFEVJGoZx6giX5Kxj5boL2PXqy+jZ7GwPRXIOoChK+sx2hJHMORqbW3F7vUTHxqRQSKYUaVlIJJLToihKWgY4JRJJUUixkEgkRSHF4m2gKMqbMjNPld6dp7G5FVtuq7/qeXW4TrHVX/W8usL3mslEWUXV2xytwGR6c3iqorrmtNctXrGq8H3rkuVnNIbyymoWLl1B/fzmM+pHMjtIsXiLaJrG+os34Q+UHnc+UFZx2msra+ZR19gEwMWbry6kkp+I8qqJGo/yiioM4+3v3lPX2MTiFaswmcyFcy63B6fTfcrrFEVh1boNgKg7OW/N+W97DAAWq5UDr+/C5fEW1d6kKqxpKKXa5zij95VMDVIsToPJLB6wfAXogsXL2LtrB8ODwUIbm92BYehYrNZCPYnNbsdqO76AK51KYbZaqZpXR7Cvl2QijsVizVkqKpomxMPpcpNOTSQw+QNlREZHsVitOF0uNE1DURQCZeU0naDYzGQ2F8abt0r27ny1kBuiqCqtS5ZxrKsdu8OJppkwmy2YzWYsFmuhn8rqeRw5tB+H00XLwiWFZLT8Z2IymzFbLLhP8PBPHgOA2+vjWGc7Lo+HaGSsqM9+06JqWiu9rG0oRVNlBe5sI5OyTkF5ZRXX3Xw7I6FhHA4ny1auwe31EhoaKiQXtSxawpLlqxgM9rNg0TJsdgcXXrqZ81afj8fnp/NoGyD+q/pLSslmMpSWVzDQ30cykaB1yXI8Pj+r119IZU0tDqeTRUtX0Hm0rZAYtWzVWhqbF9Df083q9RdRUlpOaUUlmXQah8NZSPEGWL56HedvvIxMOo3H58MfKKWqeh493Z1kMhkA1l5wEZXVtcRj4yxZsQqHy0VDUwvnb7wMi9VaSMluWbSUPa9tZ8Wa8xkK9mOxWEilUrzz5tsZGghy+TU3MDjQz8p1G+g82lbI/Fy2cg0bL7uSVCqJ2WyhuraOloVL6eo4Sn1jM0cPHTjl525SFdw2M6FokiXVPn5/oJd01kA38iV2kplGpnufhtrGJjRVw+X24Pb6iI2PE+zrOe7hdLrcpFJJdF0nnU4xNNBPZHSEQ/tfLxRjgYhBdLUfwe5w0N1xFFVVmVfXQPvhg2iaRjKRIDw8hMVqJZ1OMRic2GB4JDRM37FuPF4f7YcPEY+No6oaC5esOM7CKauowmy2FAreVq7bQH9PN20H9pKIxwvjDQ0NMDoSoqa2gYP7dlNTW08iEWfbi38gHBoq9Keqikhb9wc42naAbDZDY/MCTGYL4+NROo+2MdDXW8jYBCgpLcdmd5CIx7BYrJy/8VKOHjrAaDiEoeukc6ntpyKjG9SWOFlZH8DnsHBebYAanwOTJv9cZxOZlHUSVFXF5w/wyksvkIjHcLk9DA704y8JvKmd0+kmMjaC1+enpLSc3TtexmK14ZhUWq7rOiPhYXZs2wIIS0NVNRqbF9DT1UFPVyflVVV4vH7sdmfh4QPhAsViURpbWkmlUhw5uA+P14fd4cDhdANCWLw+P4l4jKNtB3F7vBxtO4C/pJRwvsoUyGYy1DY2MRIaJp1KoygqxzrbyaTF913tRwpt82X2zzz1CwAiY2M0LajmtZe34HS52b9nF4GyclR14iF2ezzEY+Mc3Pc6breHY10dhfJ9q81WsG5Ox96eEVRFodbv4IVD/cTSMsFstpFJWW8Bm93B/JZW9u0+ezbsPW/tena+snW2h3FKTArYNNBUCFih1AbLKmyUOMyMxJLEsyq7gwkG4xDLQioLySycwYbtkreITPcukpJAGaUVlVRU1bD1T7+b7eEURdOCRZgtFuayk+80QY0TlpfAYj9YVHCawWeBgC0BJFBLwKpBdznsC4PDBIMJeHUQuschlICkVI0ZQVoWRWKx2kglk8zpp28SiqJgtlhyY55baAos8MLVtXBBBYSSsMgHFk1YGQZgVmEsBXYTuM2gG9Afh+4o9MZgPC2skQMj8MwxGDrxwmOSKUJRlLQUi1nEbTNT63dyKDhKRj87ROhM0RRYEYDbmmBdmXAlUlkotYPfIgQAIJIWrkY8KyyNEiukdRhLQzwDXVEYz0DWgJcH4LEjwuKQTA/SDZlFFOB965sIx1KoKrzec+4vN6cCLV4hFBsrhQAMJ0FVhEti1cBlBpMKbos4rxvCPdENIQwO84TFYVEhmgG/FUZT8Ey3FIzpRIrFLGA1qWR0gyODEUqcVjqHoiicLQ7O26fBLYTismohlolsPj4BHrOwMjQFDENYEQ6TcEvyaKr4g01rwjXJ6EJgAD7QKr4+1SGsD8nUI5OyZgG7WWNjSyWVHjsmTcVtMzOezBBPZ85ZwSixwqeWwwWVUO0QgcwyuzjvMgsrQgUURQiJbojDlJuV1Zn43qwK98SiCgvDYwGXCZYHhFDsDwsrRDJ1yAV7Z4lUVqc7FKU+4GIsnuK5/b2MJ89dobBrcFUtbK6BJq94sD25+IR2kizujCFiFmZVPPiRtLBEbJoQFJMqAqIY4rzDJASn2QtHRqFTrt43pUixmGEURcHpdOL3+9m0eB4HhhJ43C6SmEDVSKfTxy2Wey6gKXBhJXxyucif8FjEYVLFQz8ZA2FVgHA5zGruXM7aSOXEQidX1KRMxDWiabCZoMQGjW54sV/EMSRTg6IouoxZzAAmk4mKigpqampoamqirKwUj9PJtY3z6exoZ2k0QldPH8eOHaO/v59gMEgicW5E6po8IpiZ0aHSIWITmiIsBxMTAhHPCJeiICDG8VZHVhECAkIgDGNCPArX5YKg1Q64pg5+2iYsEsnUIMVimvF4PKxfv57Vq1dTX19PdXU1LpcLv9+P1+slGo1it9sJhULs3buXHTt20N/fz/PPP8/g4OBsD/+McJlgfTmsKYXa3IZoeYtCQ1gE+WJSyxtsWwMhCHnLYTyTmwXRRFBTyVkVebGx5mZM4mkot8N1dbBzCLYOnPuB45lCuiHTiMViYcOGDWzYsIFLL72U+vp6qqqqCAQClJaW4nK5cLvd2Gw2HA4H8+fPp7KyEsMwxIY8fX2kUmevLd3qg48uEdOgbrNI5TZpQgRAPMSFynNlwgXJo+QsiHgWUroIiFq0Sa6KAll9Qjj0XNtkVoiS0wR/7hfXSs4MGbOYRhRFYfXq1WzatImLLroIv9+PoijYbDasVivptLCPw+EwsVgMq9VKKpXC6XRSV1dHNBpF13W6u7uPKyo7W1AVYVWsKhNTo4ksVDvFg64gRGA8I7I3nTk3IqOL19I5F0MhZ4UoIn6Rtz7y1oSiiCOVEwdNhWA8N5uCcEG2D0F47iWxnnXImMU0UlZWxiWXXMKiRYvweDxks1nsdjsmk4l4PI6iKFitVhwOB+l0mnQ6TSqVIhKJkEqlWLt2LWazmfb2dg4fPjzbt/OWMeVSuq2aeNC9lgmLQEc85E6TcCsMxAOf0UX8wayKnwfjIiiKIvrL5KyItC4CnBZNxCjyhwbMc4r4hzkjXJN6Fxwpbq0dyWmQYjENKIrC2rVrWb16NU1NTSQSCaxWK2azmWQyyejoKCaTiWQyidVqZWhoiNraWkpKSkgmk8TjcRoaGgC44oor6OjoKLq0e66gIIKblXaRR+G1iAc9H6fIWximXKzBqk0kZKFMZHHmg5pGLudCAbRJrohJgczkxC0FesZFgVq9W+RxSKYGuZrINGC1Wtm4cSMtLS243W6sVivxeBzDMAiFQvT39xMKhTh06BA9PT3E43EikQi6rhOPxwkGg4yMjNDU1MTatWsJBAKnf9M5ht0EdS4R2HSbhbWgG8fHJdK6sBbyqdxqbsbDyM2E2LQJYUGZSLTK95HIiunRWEbEJfKxiyqnmEZtcAtLQy7INzVIsZgG3G43jY2NBAIBbDYbFosFXdeJRqPYbDZKS0vJZDIMDw+TyWSoq6vD5XIxOjqKw+GgqakJl8uFx+Ohrq6O8vLy2b6lt4xJERaFlrMSVGUimKnnBAKEAKRzsYqMLoKTyqRrjFwORSw9ERjNT6+achmcBXcmLzq5vjRF5HRIsZgapBsyDZjNZsJhsQO6pmmkUimy2SzpdJqysjLcbjcmk4mqqio6Ozux2Wz4fD4URUHXdbLZLKqqEo1GCYfDmM3m07/pHCP/wIOwKvIuhs6EaJhUMZuRNSbcDN2YEAUQa1UouQBn3o3RJn1VAVUVeRuFNPFJY9AKEdWZuvNzFykW04Cu67nVurVCnKK/v5958+bh9/sBkaiVSCRYunQpVqsVXdcZGxtD13UMwyCdTmOxWNA07aycDcnqMJISz2jWADM5N8EQLkP+4Z9sdeRzK/Jl68msOO8wTWRx5q2NQg0J4rr8OhgwUXymG8JNOceSYmcN6YZMA5lMBrfbjaIoYhEasxmXy4XP58MwDEwmEzabDZfLRSAQwGKxMDo6SllZGR6PpyAeqqricDiOC27aHU4s1rkftYtnxSpWwbh4WAtCYMBQ/PjpT4MJt0RTJwKfidyUqFkVAjB5N4D896oiRCWRnfjZQPw8GBcl61IrpgYpFtNAJBKhra2NYDBIJpPBZDIVhCORSGAYRiHnwmw2k8lksFgsqKqKzWZD13UymQxDQ0N0dnYSDAapa2xi6co12B3OObn61RvJGnBwFDoiwsKYHKNQFCEkhjFhJeRtp4w+YQnkYx4wYUnkvy9cl4t5aDmRyOgir6I7CrtDMBCfwZs+x5FuyDSQTCbZsmULjY2NJHMPdm1tLYODg2KV75ERrFZrYToVxCrheeHo6+uju7sbTdN4+eWXiUSibL7+Fva89gojk5bqn8voBhwcgUurxH/5lC6CkGYVKuzi57x1oRsTrkNKn4hHOE0TFkTeOpkcrMwLg9N0fF9DCZGQpSpiRS3J1CAzOKeJcDhcmPXwer3EYjE8Hg9DQ0OF6lOXy4WqqsRze3rE43H6+vpoa2ujv7+fgYEBnnzySYaHh7FYLRzr7FxDVnUAAAeRSURBVGD5qrVERkdIzvFCMx0hDusrcjEHhKWQdz3SOeshn6Y9uQYkq4vpVjUfnGRiajWPogihMOdmRPI5GEkdIimxrkV3FH7dOeGiiOvk3MjbQaZ7TyOJRIJEIoHX60XXdRwOB+Pj4yiKUkjAcjgcqKqKyWQinU4zPDxMKBRiaGiI3t5etmzZwr59+9B1HbPFSjQyRlf7ES649Aq62o9gzPHAZzwDZTZRBVpmFw/15JkQbVJyVj7IqSpg1iYCoG90PQol68pEFmc+zgFCKMJJYVn84ii8HgKn20NDUwtefwmGrpNISN/krSLFYpoZHh4u7GOazWbRdR2v11uY6RgfH8cwDLq6uujr66O9vZ3Ozk7a2trYs2cP27ZtK7gxo+EQ6VSSbDZL37FumhYsLGwCNFdJZkWlaKldZHAGbEIE4Hh3QpkUOdPUCSshLxCZN8Q78kVnkwvR0oZIzhpLQ2cEfnsMnu4Sgdbq2npq6hoYGw3T13Ns2u/7XESKxTSj6zqhUAhN0zAMg3A4TH9/P0NDQ8TjcaLRKB0dHRw+fJjXX3+do0ePcvToUXp6eti6dSuRSOSE/WYyacwWK6lEgmx2bu/UNZoSbsiqUjEd6rEIywEmHvz8OhT5TM7BeM4KYWImQzeEe2LWxPlsTkQMYyKPIx+r6IyKtSy6x8W1kcgo8+oa0XWdy666jqFgf2EfWUlxKIqiy60AZgBVVSkpKaGyspLy8nLMZjNjY2M0NTURDocLFajBYJCBgQEGBwdPWwuiqiq+kgChobm/5oXfArc3iwVpWjyi+jTvZkDOetARKd06HBsX7osn91eZyWVlFqwIXRwWTbS3aMKK2RsSRWOPHoZne45fh/OCSy7nlS1/QlVU3nX7nezY+mcOH9w3kx/DWY3cN2QWsFgsOByOQrKWzWYjlUqRTCYL06onwuX2EI2MHfe9qqonTNiyOxzEY7FpvY+3Sr0L7lsj6jXq3WKBmvziNnl3A8QDnspOLKuXF4jMpOnRfI1JPigay4iNhwbi8Jsu+N5+sUXAZDRNQ9U00qkUiqJw+TU38OrWFwkPnx2zS7ONoihpmWcxw6RSKUZGRhgcHGRsbIyBgQFGRkYKhWYnQjOZuPpdtwBiF/Qrrn0XwAmForyyGrfHO3038DbpisL9r8P2QeFmDCdyrkfu9XxcQlVyQUtlIlszX1iWf13LCUxKh8Nj0DYK/TERo/jZ4TcLBSDS7XMLCRmGwR+e+RULlyyf/hs/h5B5FmcBCxYtpfOoWNNiyXmradv/+knbVlbPY/eOl2dqaEVjADuHRTWo2wLzU6KE3aSKwGc+PpG3GNI6ZDLCwsjqE2nhGBP5FYdGRd/xLLzQB4+3i4zRYshmswwE+7HabHN+GnquIMXiLMDucBKNRli4dAXhoUFCw0MsWbGK8WgUu8OB2+Ol7cBeFi5dwdjo3N3ZLGPAtqCwDG6ZP7GEv2GIVbknWxAWVaRqq4h2rlyZe0qH3nERmzBy7V4eEBZF9/hbS+0e6OvF7fZKsSgSORsyx5nfspCe7k6aWloZ6O/F5fFidzgYGgxSWlaBx+cnHo9REigDYPeOV+b0dgI64r//cEJYC2kdtgRF7CG/90c6V4nqMInydAORrNUTgz0hEcg8Ng6xrLBWnuwQbs5bvet0KoXJbJZiUQRyWb2zALvDwWg4xI5tW4iMjeLzB/B4fVgsVmx2O+1tB/H4/JRVVGI2W9Dn+FQqCEvhpaCIN9S5oNUrrIZdwyIfo94tMjgj6YnFcaIZaBsBn1Xspr5zGLoiQkBGTrOmcXPr4sLMR2NLK+1tBwEwDJ2xkfB03+45gxSLOc7BfXsAiIwJB/3A3l04HE7GRkdQVBVNVenv7SHY10MsevYUQuQtjKEE7AvD833ifI1T7C9S5RAuhoGwLrqj0BfLLYSTEfkb+fqS07Fu46UcPrQfm83GJZuvKYiF5K0hxWKOk0kfv0tOOpViNB/Vz2YLlsRIaHjGxzYVZHP1IOO5GYzu8dw6m5NSvXVyi+K8jf69Pj89XR14fX6aWxezd+erACiKimHoKIqKoiiYTCZSqblfzTubyJiFZE6iTzrOJALT3LqEfXteo7l1MYl4nGwmy3g0wjuufzepZIINl1xOIhFn5fkbONZx9KxcaGgmUBRFl3kWknMau9PBeCRCXWMzB17fhWHoLFi8DM1kIjo2xtjICF3tRxjo6y1k0kpOjBQLyTlNeEhkaD712E/RdZ1kMklFVTUdhw9htlrZt+c1vP4S7E7nLI907iPTvSUSyWmR6d4SiaRopFhIJJKikGIhkUiKQoqFRCIpCikWEomkKKRYSCSSopBiIZFIikKKhUQiKQopFhKJpCikWEgkkqKQYiGRSIpCioVEIikKKRYSiaQopFhIJJKikGIhkUiKQoqFRCIpClVRlLm7yYREIpkTKIqiq4qiyBVKJRLJKZEL9kokkqKRYiGRSIpCioVEIikKKRYSiaQopFhIJJKikGIhkUiKQoqFRCIpCikWEomkKKRYSCSSopBiIZFIikKKhUQiKQopFhKJpCikWEgkkqIwKYpyWNO05tkeiEQimbsoinLk/wF54xEX2izE6wAAAABJRU5ErkJggg=="},{"background-color":"linear-gradient(to right, #f46b45 0%, #eea849 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/45-degree-fabric-dark.png" , "items": [{"x": -622,"y": 444,"w": 2791,"h": 472,"type":"text","text": "","text-data": "RGFua2UgZsO8ciBkaWUgQXVmbWVya3NhbWtlaXQh","font": "sacramento","color": "rgb(207, 227, 242)","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -615,"y": 771,"w": 2768,"h": 315,"type":"text","text": "","text-data": "IA==","font": "raleway","color": "#505050","font-size": 28, "font-style":"regular", "justification": 1, "align": 1 }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nGS9WbCt21Ue9o05/3+tfa6urnTVXHWAaEQnZNNHQDBgBygDiROcxrFjuxKTqjSOH0LsSuOXxE5VKg9UEle6Iq5UhQcSUsSJQX6QA8aQADEQwASEjSUwkpBkJIO6c/bea/1zjjyM7xtjrsupku45e6/1/3PO0X+jmfZXvuNr/vpLT/ZvBmCA+wDQDTAYHDAH4HCMCbQGB4AGYALoZhjucABm8fMBYDPD4W7dLL7A34/pDgO6mfHHmHBszdDMcEzHdHhrZp2fOKaDn/ZmZu7uAKw3cz7bhrsbzGIHjr0ZAPgE0Axwj/9epmPvZtfhmID3XAUwPE4ABnSYDT7d+T8D3BB/aRb7P6ajm6Ebvx/rwuGObsB0oLf47+S5Nav3mQGnbhgTmO4Az703w0Scq0/ADB67g9d+zA6PfTSDuQNbMxjfC7h3M8CA63BY/MqvE9ZbnI0FfX26o5nprEx7HrEPdwBNJDNgTk+amhnG9Fizw3qL9d181uDdSB/E73vDQnMnzWO9Y+oBQfMZZ29bg884Nzumuy18tDUAFr9vfE8z4HI49t7sOifc4UYaAwayY/CuFc31erFvfCZedZ2OZrH+MWGwOPfrdGyUhzgLh5PGrRkgGTJg34Lmwx2GIExvwJw6HyfNzZx8Srmyg8Q1M5vu2HswRvCTe+P+rgdgzczgfsw6E27Hh/PMgtbmHr+f09EoW+JVM+Ajn7j86PbaJ/s3v+Vsz5kBsXTgIPOUQMfPmy1CxYOYAE6LsO89Do7KBjuFJ4hgaC2e4RSerRkOj3c7CbWZYaOQaR0eSgY8LLRGAnooHKwMzX/3Fut+nJ4EN4v1iZDroQz+0N3RrMEAXD2UmfM9RhGjwOKuN1ymp1KItxt6QxJx8sy6AZcRZ9ubzjY+d53x73NvVI5Gpl53VETv3IeeKyGREm9cz3U4NiqkZsDDiP0k11AVHh7PkeKf/EQzk8An40w3nHool2MG0x2h1ADEv0VjKcxjep51b0VHh2F60Ls3w6qY3OOcdDbdANO5lUAHHUlPKZxLKMhUBtfZqMRi19ZCMY+JVLCN/HLMWLMUm0ihz5w3w4XnOBbN2M1g3Psgz7VmuA5Ha/F7R/HedcQ+T5slXZOFrZRus+Kp6wge7D3eI0O1tXjXmB5r6wYqVjxeZ8iC5fbDGFDJawfaa6PiEt81A8Y8ffN2R6bWByeJ1QAc3JisotGKGoDJF28wDAcanMrEqXBiAxaWOjQtCbEy5JXEkmClNZxBjMm1GYABT4YGgMcx07IfDjTzfN5wR6cAiaGnA50n1RuFd5agmRWzDndMHuoxPYQjfIvQ8mFJaUmQn520LMbnODwZ+zJK6IY7zIqgZlKcjk7FuXgs2Gixg8hBG3kZV6/zg3kw6qSXAccxLQWsWXgzlzGpqGKNnfuf4d2FYjQLulIxT1rCzTw9o0ZBMwsjszfL701y4HWUAEwP6yXlfUxPC3cdYWymS1AcoMLQ3h+vjt7p1dI4hQIGxgB68zRcGy18oyT2FkJ5HSEM4d2sAqH3ODAN+xaGA+LNVudPTwpAnFmnYMioUtZwPYrmB70S6d6gOfIMZAQGPyAec8R+ykOoM9V7Hmfwfxg7YAwPd4x8eKKCg6e+COVocRZx5qFEmxvloWi7dWAT0WXMNjJFM8PGXWpBYMggZXBQMWwWC+pkGDPgxH9f6J5JQTSU9pSnskm7zXKjt2ap4buVBZa1kgV1KpzW6pnyTrS3jQpxp7u492I+A9LKN5R1cxeDBPHuuuEyS8E0KysZz/Fct1FJXCuEolW0xdrF+u46QzmzG2s56Z11Yyjm3A+CWQzx+cMd5x7PPaY8H7myxn1L6cX79Dl5VGL83gyzlfegPxKyw+lB0MpJsR/uaAgPs1sw5d5k7WlgbNmb15lDZ0HBP2jtZN20ikkh7i2Y4MpQTzT35JlgeFlS/WzvNDyk+aYvWykBLIrgmMCTzfA46HkOh/HAJNh6XqdnMP3WwwphJB34szkd552enrwMHsycjg0v87zScynvZkzgvNNwKSTkejr/of0d+b6gkbVQgGca4taAja9wX+SUHsYxIO/JNwMsYy0FaSSRfiaCGT/X+BMJ75AVyO/Fvw9asvsxM647p7aMjStMmU4XbYLuXRFQTDbS4pT21hrcw+JPD8u5auvpSEXWjO4nmW0nPiDvxLVvPrkhQqCD1nB4KSQ9d41TpxZjuLFumCFYc4YiNjLdI93lwbV1a8koQAmBPKbAcIzM4TfeSLrBk14SLZ+socIDKUi5sSKmc/2rQgeQXmHS3B1zGtDiTOBIWg9MNDPcH87wI+gxJxAIiWHv8XM91xnqjXn7HilUeSJNZ5nroDcAUNHEf/VMyOulsM5Bw9HlQVY4MxeDI2GRsp+u8/RUqjrPDGm5quss70gPnzSgEX4aLsctLwX+UTTXO670mFIBWWBYWweO4Yn7xBqdysQXo1rnajC0HvtUGCpAbogn5TRwDa73ktc3R4BCEyhiUfDExMaDe7I1LtxTUES5h+GMk29fHESJD0oZSTCvNO9SM81utX+nxbgC2BCCPQgcAQW0Aki3aUvLHT/fuJCV4YvhpKhClqcD1znprocCeBihktqyH7fQ4GbA/THRmuFyTAphMHQ3xvu+xuKB/4ihLqMYtvPMtPdw0cFQr6yZI4FIiLRS6AqH5MF1Kmj9EVNPlFW8TuEWpUgatcUxHU82Wjm+sytmMuDhKCC3NYWrloCymaG3eLYUx1gVDwWowMAIfz09B8PegOHl7enz4BmZEaOxwp7irCiwUgZi7CXUGiToZZS30xvweI2jNRHDi4+bOR6unuGM2UpzesHEsNxLwR0D2LunF+ySHxMnlpyJj0x8s/CzhFehYXpgOgviGuB2p1Wo6TTI11EGdh6xhm7xncMdd3sLXSA5i7DPtlBEBT5poQI5D3dsBvTeCEiWCy9B7Ysgn+j+jYVhNgviywvpLQ5gp4vqYjAobotDO5H6+vl0T+E/4GTMINxmhkHOuAwPrACAL8AjvBhKB6PDNzAzkYxRno/ZbdgywkDCl++IYc2KcGeeiQRWGYebzxY/Mm6uzIRZCbawGcjaQQqBTIRgeinGrRnGcBzueb76zkSBosIqFBJqf5uFK2tAYkf6n2guD27vy/cptB0Erj2wpp3K01rRQLE7UEx+2kRzeWpWmMYsELYxFNIzHg9PAXCUQpHA6j1jgJkNhto9XG23JZzphWVovwLpIZrPUA6K+5XVONPDkXcoo9IJQBJWoOIXbuVUrMmmqbzMDAcB0kHaK2xvBlwIWE2uexzE6KSUZ3kawsDEg+U1Fdi58ecb9+iuLI1j2xu8meFs5XqlbLnSfZY4wfRyX6+Lhd95unuTd+CM+z0xgxsNiVIwElRZ9MND+EuIQiPWOsgY5snMaQSkdWHp0chDWhkCQLqLpy2YwRerB5QgiVk8fxbnpJhdmIBSyUC4x5kWRllvA3DuApLpQjPsAhxj+blR6JxrmzCChnWeyhAFNhB7FMjoC1hqVNCHhxJzBHPZosjFqFJU5DXS3SsDA6B1w95CCZ2Iu3TIOwP2Lm+xzjNdbr7sbiPNXSB0fViA+svDT9F5VZKOyny1xVrre1IqrVnRnOcmI5DvbWWclMHpFPLIMhTvOJbMAQUuhNZu1mwwnLdbkHTriFAOpRjkkYn+7iDtkaGElLG8zk73e++VAettVTbBi6e+nJNVogH4ve8V2Dn584OA8Ka04lyIIWY0pggv/IyIeKKQ77LaYnordF/PW+PCrSEVwcU96xQcgWs0WD7LEMqoQaFNRN8Hn3X1QN7jrMKLUNysWEshlPZ3E6PyVLpZpD4p6FtbrMkMhaSDbFaejBi/m6VSUBi34gITXqkvKioJ4GYWYQ+/I4smxTFnuacijCyWlOv08B6aKzY2HHCcln2IIZz7fxy+CHgdOGUswoAlXjWTF1EKFqSLrGwz4CIltigEAcTCrK5LZur+OlmDIM4zZgws6dXJ7EB8d2+WYd2cwnoMq5qXB6PsTWJkspAtvDCFRjc058IbPaESwAL+JYxKnToKc2it1g4rbE0CCAssYsx6hiy7+FLeqf5cCa6euoTYUjERmsH1CK9s6gfwm7Tw4xEp2kHMw3Vui3zEe+KdhnjfMR2nDTCDt+nAwyyQTbHd8HIrpaz3Jf4PjAMpHMf0dOuHV9ZEFneniyOrJlfcwe9Ja6Ks975YjyvfqVDp1CoTEkqC7uqipJpJ2eBGaXS6fiqGMpTbOGnl9GKlivdFGSgjcOWep5cVAoibkEi79t4CgOzcQFjYSqvqPdqHQNDhnqk0AHWuXmtWtgkU1I3vIG+mKOo9Dscj6z2Gewp2gInJo7HvXtZP1na6Y1DZKx24psrd4wx2ruXEZwgT0NolEMJXzMpiS0gkeAYjzaOOYBAX2Fopik5FYobMJjX+fWt1lsqyHCMOZqblRj4HCO9I6VSFAMdwgrM6i6JLGJPYQ9K8Ldm2VmlheUFmorkVzect4KnCK/E7sGRzSNOdHk/Q3JPm8rBDYXhmOETnMf1m7wYjDTxBfMqDbXcs0RteVhvLZoqZSXCE5eoIgMhJbDFx8PW6kUVDTs/QQ27amfFu8mh+39M9CtzD0ssANb6yG4EzROYii7VQnoXcdbdIV02P4qepdaAUiiypCNrz+RVr7rKcbvTAkIxijENZhZexrgQTUHqOAFfGvFgyGHX+kZLmfhj7H1bYkta1WcTx1pQaLfxA5JDgnczwSOt25JriQ2scq5BNFYSd5yMgc+tBK2VyxKwCY8WMEtSDlv20GU6LgtMe9H2lmfdetIDJpbb0BPS9fcUkZNVhDEeRaekz06cHPRVl03TeczmzieIBR3kR+s76OR2x1qPwpryiyow1KkTRPF8umjNslYIJj9Ngs7xZGYGtWWZwDnoF4kVY4CVKp/bN8HiQ5srAzSXLRGWo8+78GStVAQCbXPAGS0S0USPLNQ0GCnBRbuLOgxoIV/Y6wyU9KIBnC8aduGXAwwNIEYM5KvSR5yB8oKEwD6AUz95YWZkhRKxZHo0KnsR8GU5kaozWAQW2ZrGXyfMQzkAsOS0cLc/MsnIEhAg8zonNAsEPy06lh1VxEZkGoOIlgY9GV1uej5FxwOzT3i0ZeDoyc9Ap1cMB49k5f3cdt3UEAIFCMm4nkdsNrRXGVXVma8SjWhU8XabjxHTcnI7z1mCt9jYhr61Ki5s0LtfnojmLjKzRE+hxfqcexmnvxmrUCKOEaSk2z4Ilj3DrOh3by/hYJdaqhWmLkGfFJiVXP9f3O9e9L4oXYIVsC8XZVu2DCotTka58tjxD3lnwWGXFpseZax1RhWs8x9inBFnrng5MplwVV7pFmLIaqKhZqfoPawKpg+/GEABs8O7oDb51Mzs1w0GxmO54JB5hkAWNh1ylLYfDW1iby3Q0C4XzOBwXCvHjrBqFK8G+EJQQn75aYwvmkrvtCEup8AIQyBUC9/QILbpT0C4O7GTSTKt5FWFFfC9FWJ6LQpm5uFwwwJpnmbaZs5q0QL4JxwMzLp0a/nGEaBweL4/yac9Ub2vGGpLAE1Tz1OipybKJuQaVASyEozd5A54MpBTsMatACfkMwzSVdldfQoR7fgMuC8fYewB5KukfGWYYrofDGcNeZwDRvYW10vk8HosB8JmGguyYGQH38viuU8JUNSNSKNMdF6Ynn10mn2WJo4XyjBher9l7PPPcC6tIiwnHeaufizZmyKI34WPXwezCBHqPFKQyLt3C2l+OAJSvPLBjegKeKeCIz+4LgST4oCyIXmvG5XLofCe9i4ixLwdxIypskirbC9ZWAq3HrMJT8bh77Gdn/CsvY60UvQ5PPnu4wjYVZKnqUC8/PATuoICcmqXwNRI13F+6Vi1qErpVX4c0+t6Awy0VhDSY4vywrKz0dL2fyLLJC4mDOTdaeqvDlicACtmg8lBsmsU0LxMoKYq05Py+4vnLjDqDJ5tRGRYSrTr/E03y9ECcgXKl+6LZlXJeq/Muw7Ooa6fJcb9N00nJSbg7vQt5OvroQUbvUAZB1spvalEckQpXDJ6enVUFaHh/FXtfp9+se2P6c29Va6E4n48K5Y9KAysMk4sOMERhaAB6rcND4MV3DifmUc+XJ6A9rB6DQq0p2sr6cI15dguPDnpGxvTt3d5wt7PmYoSRUxHU9GgEE9Zx2piWdtXWhHfkqPX0FilbWCgBvVs9R46iubKITsV3THqXqDBSIfoxPUNa80pLFy5SNTkqdEyeWbwao+exdcNpa6FwB9C3bELE1oBtunuzxr6LIGiUggaTPWktMYY5q3RbZalV0Vh1GU2ani6hwRIrkFBm3QAiJdjFBHaL6NJPyLJd9VeMSZfVV6CIzwBBV3c86S0PRGfEOqHQ6qhqTlmNiVJs00Oz3vXK98Pk8VRBkZjYxRxeoGUQhX9fYsNTl6IULuGZSdEfuaWrYvXld8Oj3NsB+KTHIdfYCqRWxsVy/Uonxlmeu5g+SsIF+q0YRAB2lf2Q5zA8zjTDACkUFKA3l6xShjgCPpfvFV600ryUi0IxWBRIyYg0eqbDgSd7lbTrrOTyy+IH37CYLdOKSED0cOBut6xHkFHUs/RcpTalTEVHc2QF5mQbQ9Bc/U4qXS8lvNJc3k2dS3ymMeQ6s/pQ5eDXMbHB0DM7xToVVg7DC38TDqGaljEdd6cGd08QX4p17+ENbh3ehldqVNVj6uKMmguJq/5oY2F5Q1gcF25YjCaGAICHMfFAl1aWf9CFqDqGcg13Mvp6hMpaROalcskuRuDPx5TlX7Iefpvl0J5UUai/i1mnR/+H9iyrrs81Ay5jwr32pJoDMfv08lIeR7jqSqEFk4HgYBBcrc9PttuT9mWPa5epo0rQL7OyFGaVWbiM2rvc65nPQu7HlveojsKBJa1ZtLgcM0O2y1hozu8ptHk4HA+HzqfOafURxJjCY8SgRfPgs0kmVum8uypB7eb5kXFSNoFp5ZcJ4sFQDjy/wtTCEEWYZmmJzeqMLsPz3ENxKVRd1jWj2e3xCGEXv8v1l9ens+8W9SaiwXrW8h4MSGM3RqzlOjyzRVHJSZofnhiS5NAXehkK4JSXdYziAVWX1noi3IqUq5UwNGN+PT6TAiDXG0D2SUiw5CoqJRppIE8N1szgDTjxmRtjqmfhN1ep8mLt1JPyJNNoBDwb4LMQaMdtbApU09jkM8VAjnL1VAm4E+hRtsO9UP8Vq1qt/SRDFNhqGW4BpfRkpZT26i08kzGr58BYVLbOxHDEmvcWtShyZiKTU9kXc9a7gC5wK2AVfMZGZaxaACnErS3VfGDZPcOXleYS5g2yfgY1kbkjPZpmakAs4HRDKRvR4Nkx4cxmGJTpqdRlN8OTHek5yIWHV5jorgInT7HSXmXh9x6M7YuBuBL3UWp2LJKpCtzotKWgIQBLYWnWKiu14g/dKs2pvUdFa5yTKiHDna/yALQFtCSesPXqB4EVhmWmk1ffiSf43MlfCOsf52XETWaFfVG0pSrQADCtBWNX3UWVQwAVokiu2tUL6W+LgIpxVxBSymSiUNpMvdFSXpiHDqGM36n8YVIYs+nIg1GN1nK1uumxjIljsp6CQq7nDZpDDY6h3Ob/FEcruyKrark2MpuFdZSy0jpkcYTBJGq97se1V/ZZOLIbVwoIKM9o9ZDEKGucqXffj8niKE8FLqUnZaOU8anbjTJLxYuq5XBXDt9TaSgsuGN8NehJKpyIMvCgaYUjjmOU8jGENTtG0GstalppWcVWtR81tmndasQLHopnSXjEhwqNKiZfUs9Y6zjq3TpTAXYS7LtNpfxO5VGl/XurEDSbBFE1NRKmg9b9GGX9gTgnvXcFjIPmFH1fPGMDHq6TPP97953pTvJyzMCougx9djpYrJZQTeyDP2hU3HdM68wpj+JWzh9p9YSrXCewGcw0vMXcwR6aEhxiFxupoZJfKYIsuzUko01UqlW/MwrUJmKRu9c40JZ/qwnqzBeo78NRlv/EGFoWQASiYQI8Bt8IFJKVBq30dbG01xGl1irdFpHV4akKRhFAf3ROYnx15RqK6aI0vOLFOeI92USFIrYwoA3lCqe3YmUFzz1+l6MiLIRsZxgjARcDa4aFvMjLQJarz8MXZmPogkoNAyxAWyyovKlJRpNQquxafw6PFKZZYEnA7awEKaw4S9J8Mzgsmxmhc/PYR8TlEkopWtW3SJmyroY8qHdI0W09skvTywuR4MmaapCTOlhFUwHqqUSo9JPmvWZsZFPZkMdR4XN4ZEFDGTelYJWpEV/1ZpnVWz3py1E0f1QzDjXeibUVMnaPR8wCmUCuWUZ70AlQyX1HhToIb8m2RG0XQdRCpGXU1BOWMtKqEjRNWGpQFV/Er3ur3gwdbmMqEYtisAVMlAJRCkugUrjLoQx2AkkNSlnqXczgcC3DgUf3G49Fzwr+i+dPlKu6L0xsKEFXEU+3Elyh36tgGCqksCbm8szhy62XByQBaVZK1xcrIYFsqO5Z9cgIwF3LhddSbIFcQLnKa9aoU7AkiPlHWSsUOOmouRCyrHK5hcYPCrIETaMBO9eKhQawZd9d642zihDJUrHq3QJVt04B6AVqBq8asSZOf3KHm6Z5eaZshXsIC9iSdwKv2DtwjMKStG9AmYeiuP4WVZoVIk5UwZx4a62faC2URM5OmZVK1jNU9OaOLDYcVEy9IUcRbJ3t/wynZRh7Mxzj1mPPLCXi3A0MvSTDVlPRpPTKc3LflBYVmAOU0jgWjSrvwswY44Zl17xJ9dzfVFVSXV8mPRNgSeN4uaiLpgUPS2Cr0pPspMXjdaYgKe5UOnd1aUVECb7CATFso+UWNqEUZRSoxWGokErfUSpWViDlCwV8aj273U4BoxxmeBK/W3puZoUtiZb36id5UOt8IzOYmLGYZExnmlarFACHGyXVzKrOwsT2SnOWQhO2Y4uSPG9MIy77U7GQlIgj0PkuzMmrL8hpxQYLzdosAVGaTqGVeErpWYfCFscxrIyPlUdQLezl5sswhbJhdmIVnEXQ5bGIxuIp9YkkLV3zWmKPl8PpvXnO3DRqexmgMSoTJp6S4VnXop/fX+m1mMGaJ/3GNBzLvBCAVZ4uzAWYjThEC6xDHbaSB/3pzTCtvHHNuzArbPJM4d1OZh4WkfgBqBCm6iioPCCFsAyEoaKINFd87nGGq9u8Nt5IYPNC6mVpcvair/MMQxFdFuuYQsp/a9iprK8Kgwp/KWbICVmtUmlnfm8zZCMZ4FXj4OV5qFS56UCBLPqCzm5WLYeQaTVZwRRfhyDIUzy18pyUrXCLwqgrrewxqho1B8FKmfCMcqamVZOTShPkrUnozXATXoSwLdkwW6sGnfU2EgDLtKxZVWU+zihDd3lVBgyyZDO9O7SeI0IwWf8BJAZx6lHMJ68n3hhj/IDCNaRxs7YCVY2oVOZpC2aPvQSxzz2wgq2zxkXFSxRihZPCotS/ogbCeC57mxCKQSUDKuE+b1JydqMYaH+Y9anakPA4QtCPoYpZz/BXxYDTLQFcVbLG6YRRiUG7pDUxLAHMqsS0sIo3odYgf0UoRgXE82iUiSvPanPAnh6ezT5XMocsh7dqNIqO0aW2gcsVoDe8WsuVD1+HnYRFX7QzyipPdwxUIVbEc+XFTFTI4oj+BgGWg8w8PRq31gzHZqxObEjBcq9sjdy8Z8fkcJ8CMQHP6kkh4iK6piQ1K2ZX9kUelhLPOhMx+eS7syBmVgXn6sqrIlIhmbpbJ5WvxglIQW4LEm5NZe5yWQP/GQTzHg7PztVBI9DNEqAc8gLclzDAKtVNiza94twTZ1bKOovm61g50V0ekTCSwIpYW0FXaXJznZZ6b6rYRAqHMAdAoQzD08XS73TV5fXK2j+7OJ47WdI8PBRjUR75WeXr5OkAHitVurH+xsxq6Ezue9kzw9YxSxHBw3jsXWGn39KcSkDDdx3CXBzO4df7Vh5UN62vPAxNEp8zaL5vlucHIDMwjviZ5DGa6KQ0ADOz7eru6tVwIIejaMZm9+p425lyu3gNpxEBJPhSIEJo142U0CPnMjiWONbLBVNqaKegyfsRI8MCLJ2G9O+FU6hUXSXjZqEEJxwqZ5RxHTOeIe/D4Yny925pGZtScR5VgWJ0xdflzbBIKy06iWnVLj3jBwnUZpOeFa4RAGZNHQOE2yyYhleYo2xD71QYXhkR8HePY2Kdt6lQUSj6QQ9qBa13eiuPnMV4WtYVJKzuzsJJbrGZ6Z4YCIpchVuJfygY2Wg1K65XmleNVi4PZgZYK29JGEMzLHUITpqXew2EQFwOz5Q5HGi9QpDOtScuM0vRF7ZEfvQlpOT5JQ28wqfeLGeWpHXn98/bqpSFb1QquzXDYVULIotfWZFScuZhJFQ2LuM4qHXo6OE6IqNT3mkUC8b0twB3961hzIltM+RczAs9ClnCE+oBArcmCAS2SGAKBAtPIA5KFlfujoBICWlWF6IGv8jyhjtbaP7KXI7bgiSHcJNydxWTaQAOluY4vU+fUWONLHvLMIWNNmZovcqUz91g6+RjCpnccRkWhVnyHoQHdSv3buP6VIFXMMM6dcrSc1jBqXXwjoqVVjC59WLyJ1uM7xOOYXzPxjM8OD17IwPuzkE6KMuv0f9iMPhSX0Hh1ewRMWw3zhdF7GNr6j4twFLh2YkhrIqeKFcA9x/CaUlz1RpEw2PQSiEzxL9WAqs2dimBZtWT0loZuYmqDZpevTcKJ5pFJuvGm1lwPdFJIaneZ1Z1NvqcQNBgcE+wVlWnNzSnPGxap1d6HOJjytGYjic7FUkvLCb4suE6HWNVDi08QkOB2lIoqs2g5+zbRN0l4R5W1qfX6DUgh8mUe46MnRXrdaifhBOb0msIwuYofgsP5XEaY2IBdGxBJ7ahwToTAkJppVulnkJwFiXB9Qpz0YTp6cAV8W+5mEDkxuUxZzhghSscCJsh2gMAACAASURBVIorG6FwI84oGPoGKLMlv71Ydz1fFwqhyVWvcw58wUpYUM1twSARa2cJ8RLvprJFWU1ZpgcCYarSlaJLMHKJh6fPFL4QQMvhzJMLq72pXwQ5hWuR8RJSKs2d+Iq8AdWYAOVt1uh7T2tc8zTLY1trNkRz4OVXCdS09cuYqUyVCnUeksIKJy3kVUrAQ3DjxarXkcCmpzAlC8r6VZbsvDF1jvIaw+jFJ0Km1rJ0z8lbUkrXg5msBURXiBB/Lw/dofDVeMcIoLGJ1znLUyOfjFGJAG1OILqjvCkzoF0n7CCBRGTwQMSE3eqAdAjurHNAZFMu/F7ObFiYqnRv/HkYlbtu/D4gK1UuGAw5NEd/NLot8AuWuM7q7kxX3quDTt6P6iCmq9RbVnrp3UB5SjoHLEpS1vXcq1dEabhMq871/Grnl+HpxQj32ExeEd0R/olW9/IypDz1LGUf1np+KQEROQSmUr+D3kYWznkxuDarKkYx/FxWJRCyU/HJW1TWIt3ghXn1vYejrG2zGtaiClft3qxKv5PmizEQL165B6cR0TujeM+z2GiSB+QdToYta7jiuMXhdBiu0MLiLM9bdY+qolXv1Rmusz3MQnA18NhQQ3GavSxlDdVZaGDPmhat81RFZmVtiDl4FaJpeM7698uogjl5N+vfDaEkhP3pz/RQeL3FwN4bRSDmXHEI5wPXzYmAEw6fIcRqJHOUe9Ys3BtlGdabr+Lflf9XIUs24+A2lDGoZ6OerfUrZ6y7DwRiwgo3SSHWwbvqNqo4JohW1aJzOUwdruLzOhdLhlGWQt9JgHc5X7mhaU1mZB5Uo/E4fAmvorz5qhQMbrGL6ZWDXy2vFH2NoSdjWAnl8FuaC1+RYArPkMC8fN9ZozA46s1jiXVGhT+tXqnSzKJ5hhAupROfU/m6whmgUpVKO08PTzj5dJa3IS9w5e/Da9BwDHiJZ2nsX9ZoLEQ3WE6YuvUMqhq22sWlQIIXZdnhNJzrlRA885go7mjCLJrhzHH/KW+Z6Vs6WScwNZWbBjP6jarIDqK7DAMPQvRZM2xaY803rRaFMd03s7hLUZqd/JYvVfZAbpFTUXSr2QMCFXXZ0ORTzj1cTz1X8yMyfjTEEFov4QUijTRpTS9ORQQKJV3Qq9dNW6ded00CEiBlS4IBBI6G9SEYuLiCM/fNYhcyt0BSB3I6ts5KrvKZhUThZsdh3l5th7QsDsXacQqaIxAgm6enlR4eaXNiu7JS1mEJLHGRU1rKVZGwAtbKdVffTe7bV5pTgao+wgo5j4t/xMw1C6GbwXoJzLnXUF+XwKMUxVrt2VDhkJSn7lLZGGK1hgRoVQYOQ2U6qAUVllUlKVJpgzTfeoSPKmxTPwTIyxutmPYpxdkW3lH25sx4Pslr5c47UHfrSMiZMQGERy1e/OR8zMXaG3QXirJUDAUa8SaP7ygsdRRucWJBiEKVScMnUDjOxAL4XbwYgbQZ9hPTCxqx70oWVKDHpEDnuDKrqUfS0geYnrTCBh6oVPS5Z4emXHGGgleH5kEXWYqkMT6OEMFp5Vk9R2GXFYrXLIU0jt8jAGsxjYRbJeQpNK2+s47iU61AzrlYnjttLQAKsHcdaAzIk6mqvAkpoNjv1ZX281S+V3KZhEpFTKcFbNsW5tf7qy26QhPtR+XiqnOoi6Q0xIcMIEsMZOgjZVj0D6st6yiQ8TFd2wgJnx0z6zQEaAZ2wDBw+NKiben9HHSXYQ0aP9AWmmeYQObSKP5bmnv+W3TQGcmSCgQVfc3CY5ChUTq2rkcIVSqr3VpMibsMh/EKAQmYO3LilPh4p/K+HsV3oFEdDIumlI2pEpbh8gBrKGrN+l7s8TaREEaKoHevvhHd4pb/TcsZClMgLux2SJSLLs6zC7oazjSZ4ZrGAal6MMt2kxGLcOn+o5jSV6Vh0pVx2MoIuAAuL2BvFX4pJVnJNTzSAQQjoMqCKQhAeDEPBCuk9NLlbQEYSqh2Qw6PgSFxE6MAAp5FXXLhpOQUM4vQwAKaQi5oKSAJu/AVCYKEbXilvlI4gLxn1VBMrhBIYZ2hmF7KJeNcFIAoJXmm8hFOgfxdff6RAGnR01IBYllLgmBexkLCWkaGHgqFaj2jQQygLhwq4dlaWVBZfXkNWhvAnozDs9ERuL2IOu7ytMzi5MBke9lZ878HhQ6io2gOequtQqY1K6KzXOfS6rs3w5R5AObIOp6UL/Aw1zM0pDckGppFvwectS/0qNQDs3dNV4+X7Vt5X5JfhTjiDaVbwXdK3jeBg+Y16NURDKS5iOF5yOaBzAi6+TMtkvNIxLjTJQi+HGh84tQND2mV/EbgFG+5qwisLjzWmk6oRjDnzg+XdXbGzhVzV/cgsnEnMikxLpBhJRqitFp9HzqsROodrEMpT6uqB5Ft9E5FtjVPz0At3UBZwtW7magUsJSkQFozRDNSI3I/C3u4ksgKEV6uYKevgF41YRmWZ6MsPKw6LSVA7uUZ6gxO2o/jhuZrdiaHwprh1Fvc8CZl0DTgJv59aurfCKG452SyB15Q03oJgVMCD/YBeDBY8itQbenKjAgMDOUzKQxBZ92oJ0UR8Xr1nigtCVOVqkNzLDqth2p0NoaXOaSGT8yajb7QnPwu3mzGpkaXia2wcCwgfKRGy3AqrAtjylCsI2sxRFfRRArLEXM3xMc1VZwFWqyvebxG6rZcMC5eE5ZywC0q7XmVSuLP1ysFB4Vt7byUJzABnFrFa5dUFMV8zh9wT6n5NA1Ksx/JnzllWy618V2y8AJOBVxK+4uw0vKb8WKcFp89MYbezVJJKnOiBihVik5Ky2AdwL54UY6aIXGXeflaS18EuLw4ZPigGgrd3yCPJgu1rGJLkcVz3xzxvoRXsu5mZXmlpDrNXE/TWPiUPDJ5F1Ik8KohmV4xsdz3qbNMmpeicO7PqWiFnUt4hzvutureFAOv5d2TljTBXajcvQYBya0WzbNEn2e/C/PZCqOTvExnq3hbqpJR4dmYMmLiZaPCiPXccZpVKhwCu8fwRUFQEVL41By21qzICIk2quhVb4+81FQotPhKtU7+bB3+KwOi6mcdsSMK+668xUihz9bNtr3FrMQNpdnEACV0Swxrlm69ekkklHd8lsFyTJsbqAHVO1GbVLu6btGaVHWn3tLSXUiZh6GrES0n/mi9smriixXBjynPVC5mWdGpW9br4KpGorXIP7dWdRCO22sLZKkElikE0yU4FTJVvURZrbr28K43qK5Dg3wUyik0ml5gV3C9pWVY9w9UbUMaCFR3pRq1lGnpyzNW2sOrIWwSX1EIVl2U8V0NwB0eBWAKHbsHL8hbUhpZnZQwusgk2t5aerQXljw/HHU1oozLhMDJUjrUY3m+GrbrXm3mCj2E8bgjvRqnAZkzjIVoOh04b63wKhQAqOIuswJ6Nct2+lKfICUIXfLjObdT5+eQhxjZCmWc1PWZYQsPPY0jn10Deklxehkq5bblrOXB2LLeGt4TK10ne5tlr4hvoZVjKpOYLoA13BBEDDI9AL2MF7EyWl2/J2Dt8Mo9u9fvBPzIm1CFaDNkma1Sh03cwHdJWWm9Y1mfYj41fj0h0KOMhrIck1Zct5rLA8hb1iKYqfAAGkV3W4ItZtUadMO4vKfEE9LqV5wf7/C8HastZ6HSakdkW9TXIqur9GkphbIcjkprTn5eeIS8Q33XXek4DUzmLIhYXipEVVcWKLl4jb6Ara3amo2YVPVwLFgPRHOWiFtlGnTHp64pkBVcFaOUjArHWpMlNtztKkLyDGuACiMPWlOFNOv09+CjKrHWPAfxFcSzKK8lvOpQJBcVOEqp8Xl1AVNsQsVg8qiOEc87cd5EXX1Q/GsontVaNOHcvZoyVfQGr6yQ+laECTXzookMmVte8TmdpfCAqo2tCUlfJ0rvVnHvGj9LQXQrq5TNOeuGqCCuLIZR9aMG5yTDG5VTxrXxrsBROCAmCVMu7to9elCLGoVQ6wSqFiRnblgBQ82Q1wLo/RoaDAkb/y5LuLV6dyizGseu4qjp4XFpfxIkCbXixBIYEpnMrXBjxWx05WPdBVpKQT9S1+/qwQReUVceqGcmPC/LOZxAeRJtOcN8tllaUs0djd/JM6iKSyn9tQNYBW+yaGZVaap9XpfvZSiy8MXesdD8dlaH1iW6ao1xCU8NQ74xJrS4WfNjlRmSUKkbU96a5rsqw7d6EMcgfkBMaM2kKf4XX+a80AbecFa1MFL0Y/mM9i3wXjysdOd0ZBpX5x/dsVXWrXtPr3mTmOqDqr9EJQ36ncb0Ta1Zg09tEa5sFOJhNtx6GcIvgEBtVQADW8AtKRkSd037He44t8bLiGW9FLPXrIYLteNYvu+IZjFZTXkK7izPXoiivaSSMkvAMbV0Ml54RTYtp0TJik2PzMEjwSLNhawLi7lhvj8YvQhkqLBOxJB1l2CuMz2CCePDmmfguO05mF6Y0vSq2Yhzr0KbHBDUV+XAfUPCWgxrKDxDOJBc8Bxh5yGQYl6H4vYKD46JHGzjpIMuI4Yzy+Tg/atFc1lAZUHEE2OI10pBA5bA3S3NC9Vf78uwuf6++GYynXvq5VE4BSyu/FNFaVUEw1chFn2X6wAMcRfJ4gWou1M9SOryTAM7pfCX1PoozGdJX0aY6wobkSCue5z7IztMdd7y0Fqr1O6cM5X31ouu6wBi3TvCylIzWWvF7PqflEcdRjXglAWVAlEmpTyGrAxDKYlYdxA9bkGrEesZc9JyxfVrzFUvz2pao8dlP7lur+eoOUkpydVimpiRPxeTwZFXIhQTxN9VTxBErrqIq4drqV6KLO4yVSouWRS5zqhS7/IVCp9Q2KW1resLSxiey4VMLmXd6AGIboqjcwgvbi16TsvW2XlVcWpNGjCsUOUyPJk8U8VeOJH2qu9HCXIp8WbIrIMERUpCHpXCjjhiZZ3KoDwc8uJi0dH1yjtV/TZL1XR2KKOTZQZe3pjmi6o+Bs4xdfxggJ3k41mKwhavRtkWXa/w8hF428vK2EFekscOlBHW+oAK4zI08FKOZsJPeG6sy8hmO4bY+qwG4OgspRR9IdrgXtdwZE5mQ7Q+xeuK1YW46sFSAnIN1clpJJksVW5WG7Zyj+R1CLDaWXwkXEA5caAyHULWM/OCWNvDVFFKAWFXEmlFflU+nRmBZc26xPjw6mSsc0BaBsXnWQnnrFnQWYhYVKq6BEn71J/h0fUnBFr9GjURWuBoZVuM56RajxVkvI5lFsn0vNe1hsxSCLwK18Q4hvJadL2jRuSJwxs1X4Z5MgxWacO2bHHK5JolLcQzUm66ZFrekd4B0MvIjIZlZarRo3g4ihbRFVkdymrIasZ5FltUPjZ5k+kx3NafONckT5OJAGjidwm4p7csWXAUcKpzVayfZ+KR/l0xPilxhcaZ+eDvzQu3iCRE0e06gH0L2boeQG/yoApQzxJ4q5VEuB5dye6OKzuOJWNSHg0MyVoA1a3Hzjej0F/pljoCUNMAXE2LAi3nQACPewM6OIIOVaqdhVlAtDlTsBU7mxXTK6zpfBZfc0OI3RAX26K03/S4i2Qicto1SKbStcIkHMj3qr28obwXFUC512j9eE54NALSusU1g9OrICzc6+oxyc7atuIkVEJNsyzK84gdG/aNysmQ5bW6j1NhX2SoIqTQBCijYnscbJ+3KhCDAWPW5CqFUCob7qYxdrGQUy8AUQDdijnona0hLpGyQt91HkDQcZLZlAYGkP03RXNeLEVCqylPgqt9yxOcDtwfK5DH2hmuUWcH8p4mnkuRN6taHRWA6XM58t6rM1jFSg+jaKoCLd0Edt4svYgS+OADFQsOL6xBXq65Y7OWQHpvUS+is3LyutKg0YyGrLTcDLhcHee92t9lxDBrWNCFFaDpTbbbqwZOW01WK0+OZzuizkqDefZu2B6G+/2cGYaU5fXsQ1AtgAogpsvFrlulhV3AEbePAdmGnFezUXWputC86g2k/4Y7Nl9qNOTGkRnlXRyumQuF7KtSzcH4FGIKT65UHmW6ytErx3wVgamVn46ZAiQ8RKk2rTeHujqyBt94DgeA3aq8+fFQibMDk/81ZWI4bxHlUkqp6WpDMb7Wm9bagUt6IVG7MBQ2WYHRqWiZmtxbhUYZLgG8katibfGEFLLi2nBTPYlTSD33ZNXYp+Igxc7VsKUwwXIdqstJy03X2hcF7/zf46yycSlzCZz+6LLoOR3PLipyik9ExqqyYU+vZTQVhSi7o8NQ2KLCq/SmaTh0RmMaHo6ZGQ2gzjRDFA85kstvFu/TxO4Gy9vRdUoq2nocs67opMGEKROzhn+Ox2vI4tbLQMadvsKsWP/RLIq0jOE2wmu5HO7bWWDWYtGvXgwvlxOIdOqEZZooNlPfC6Ep0CaKm9j4NasG/tQt6yq6282wXQ2nUX4evhSPmLIsuthXigA59zNdObGDl8cBeiinZpxxabk/o2DJAisOV0jTDFSAt30gGvq7hqKNFrSjsIoGy/ZuM6N3FmPuYIWNrN26wFIlyX1VyrCAY3C/GVJN4UbqRTB0ztAQ4q+afw3RUT5evGAmd9TyvVpjpY6rK9G5Jo1TbBYA9SDj7t1yypb4Y8oLsFswWrw2NE1sItOIavACn9lmuMtad8r0Qo/pINhXWZry7Ni4Ri9AQqsQJwxjzbwQTXRGdFKCXu32isNmUafBXr7wznphg7stWJbVmjTnkyJYigoCji2mxAFovbComlsRa1JNxTqAN9scEOFMy/Cjvp8XNKXSoWd1mW6GVmCmlYstJk5AiFZ6MKRQmbQs4zFUxGQ5rDbG3lUbcrg5VZQir0KEU2zdbREMILsZ9XsJ72bVq6ApRRtddBEzi0/4vAtBJbUDi0FyzxBIeFtToeKVEJ742zWzFWSkFp7B/TFT0BRySQE5wprEf8tKwqJjUAq3WdVkCPvIuz5o3aQcPUEsw10vAV5xJxUVaWBQtwKO9RwJWk4ag84qhuDWfRg8Ey83/dRqvoNzLdm9S8Ohda/41USFojIaZpGBWmt6FG6YlSJXa/nWkci+6jWEbQCRMpS1l/AuzgIB0RIM0Vxp9ZzAbRECrJPjd17480gvYnrdTi7F6agsyA2/oeZkSmCFbVxH/Ez3tEjZi4dmFhjFRVE1SWzJrNBLuB630+Jl4KQ4sUyAC37klZF74D/qTPUT40ttLk8QyCYrCa9+/UAw7Zp1AlUXsDfOeySipMozHbYAx0lOlIIJNy6sERwZewNRwTlmleuqpkNKRoCYZmIaKpujTIiwFE3SPnfj9X/In2+L8srRddy0872b396qZebpAcGAh6MmMxmKqaS4kiiQta+7UB7nTAUVN9N7psV0qa5B3y+QTswfN1oVCTuxD/D9miC2lhovkUQqt/VKB31O2YELrXzGu6L50oAkRtTeJUhStFIwADLswCIYQLjwmj+BTEPGTmVxo1xZSsGzVF5nrLB0ODgnYmkgQ8XoAtjNCteQwshb5IcaES15T8N7gubIvatwbjrTvlYYnbIyws0uB/KWsmjem7m/vAgat2lueSL683jUensDrEsuaoJYf1kmRHt1r0rXDQV2AjFnw4PmtumOSrMCY046DCumEfMByOnbhxMMRaRRBVKKfbux5Dc10Co4xeQNxqGr8d0c7oLqBtXQlmZKV5Zl6CSgJmALSKzBOdS0qektp5TrwHQdQOAC8VyBctUTYrhrOuClPmNWoYyUk8CtKLYqr0rnGFWsek95LMnABtwfMxWclNhNepXnfV7c4itTlQLuRCeXFWy2XH4b9JGCEKPfxOEoZRsDYDwGt/Jz8jpVwqGzljCmq45bD0re0k21I4HTMZXFQWI1umaziq+osKyUQXgUnuGTplkphs9RfIi9XEd5WGrA02VMaxbsbmvJ++IN4XFS0Pl8VF3PjYcOYWrVM7SeiVr2H64zBXid7RqXC5UcnbcyipqUpfkWGnLjqNAw1wLRw7GzZ13VrErLyxhZi9vfmHHzLcKDEpLwDqr3Y1804oHKEGSFpRkexozMiFWMpQyEiB1nVlYBBnQvd2giQEtD9aiYWYBaPDR5I8JCtHF9XnF6VpiiSrS7EbH26kRU8Y5TM63DWtW8JsxC+73OUGJPtpbX3526JRgm6yThNETNhyzXim8Ekxfo2iw8HcXwwlLWWpStDpPYjt2ESk+YDJfwTo8mtpr1QPSfSr6j4lpAcXUJ+TErva0UtRmxnUUAxaz6I11m+XdL4ZORmLPiYrWd670qfNNN5WvVboaWqBAwaNfS29JZhUccVjXCKatwBoXhKCw4MyRQnYIazsyi9yVpvi1ZBqsaE+OGM6uyGDmhXZFt8bLsfMZI41VZLIOqV/WOUgIC0wNA1aiI4O27vVWhnQGDNQ4yngoHHcRyerVQCFvRjfN7j4zdNtztcc5cpAG4X3oaBCBKQz7MKFyRAEVmQhmQINy51SVF6mqL28k946XQXqEBH4iBNEP2RxgFSTUEQuen4+beUxFiOjhQp0pthQyrx+CBQJbavgNzWIaSwHDvMxWkui0PjxTy/SFrczt/MqwsL3uRIEhIFsFRGKb/PlDDnHudvZqbVFa/WmUN3l2rWZvdDt+Rm6xQS+lWnaVKyn1ZX2uG++tcMhTGdcZ+Hw5khaOAtINFO4MZsg6VUFsy2PRS2hoMbDyr69DlvrfgsFKSUZEqQ1LnkOEKaWazMI81rFKF5sMRHsgxSolMR4KXQF3ao/oM7aG3+L4E9vFghjBpX+3f4kEDcpobzANLWn53f2Vj17YYAKsycmulZLTO6wBDiEpnX49Ke4diLJzGmuHxOjGk1IanlyWj0izuTVFviORb4cn9JeRcSvEYwHZqLasdtamzMAyUa3zqUQR16oB7oa4DdZVAM7BN3WiNPDMPhsoaKMzRsNy7JYS4Tl41YMaLdG+VghB+eRtiKDFJCKqzci9WL08orRyqByFjN1ZRaXiwAXkVoFp8T73urFCKMC8FaqXtFX6oDFuzLLZW+eyDngvAydcjGPFklV0yWgkY0sLpqklALvnS1BbLyJhTIKxoqPtihebn2Xp1j8JsoXnD45iRkeG6JoXuvFWGKj27VlZ5HVLbDdiIKuouUo1pW2Pq8JBKO64eT77DkVc/pFJe1iBB08VVMjywygroszGThJ4UFkueGZMYDyAPWSHMKW9fDzxoZxpVYYgqOfce/RU5JWzW7eUb7ywBqt5hxSAcyPqhnZdDrbKwNvtp37CqHE2aW2SdzttiQHm2Z/aPrMps68GLJ44UsxZA6piw9jCmlyW0XJCKgDZTjOXssY+HSptSZjN2FZrf6EVcHTezMaNknK3nJNCpVfNYg0KLAPYOrxvbJ78LqFKzEH65tzokAaBKU8l1vcwSELl9An3W+Hqd3wgUyKm/y1WUKygloz95k7eXizk8zjEu+2GDFj0eeSJrM54GEwGK4z33LZBQ2k9WXFY49w1PHEfentKk08uTE/BmKG9ADVv6+ZVAnWiurJMyX1LQutckzj/oeh2eowVCIAOnEvBYNA/eUh+LlIlBNSU1Q0TnKzrJ7b6tvan7SPRvnS9IRynJvvCCQ9mvMjhmyIpTA4VtAc9iTgXrUHgWqsXQxLGtxTMEHBqqIld7rfkXPI9R9SjiT8ATK5FyUAm8e4R4el6zZTzhXEoFxNdmye91URG9avbXmEUBZLnOvoxr5/8cSJxCYNCVD3IyljTyZpyNYcD9UAVjfE4otL4vBeIIAQaKcS9TN18V4cQQV4+GJPXIxYwKVpouWra3KrJyD4V0dSOIWopBZbSrpZUbr6KlAP88QVJ4AZbNlrgTAmSRnba6WMasYt8TgaULCdNA8HDGRudyNtq7LLVAqLUQqAbplPKQxc9U69Qc1FIOZgVqD9Q1DKEIbj2GdaKW0s1mVaXYW4Rp26I05cEINFX2wxelr48/Hk4eET2cXuRaN1L0UZigJjSlwXMAsMIuWni57zVKj6Cw65kEnam4lOVQs6POJGhe+JzePR3ERaqtfFXMCqcvbExTivQYngJoPJuJ8KBUHCUscT2/Qd46knF18xgnfkHfWdocRHMZ31mlAwAy7av9Kfujd29nMvVAMXYhzJ7AXFlsT6xC9RDhVke1lzYtT0Pu/1o7r+fEFKVaoFFZnBn7SwAVvpjFfArngwy6x7QYVKXPEtSsAPWaNC3rpguCFOsBVAJe4+bis9UQNKcThFQoVUKtPaxejtzDUxPzAHvXJLE4S+GCApzEnDVkF3kjuWpLdEeEbvZeQT1hTIOuQ/aKQEBwTeKSRVGxktYrgrsBPuOzCq80oVu4hegqRSHmBOd6qHXgmAT+4JijirwMMVVqej1LlaxmASZLwTerIirR8fHwtPJSJLKaNUNT9LV01WO5hQGtrfcNyLS6lMGJ05rW4cotjQESR1Jtx4k4yCWyCfFsq9QpQAFF8FxafCdgS1pOCn3WGXFKuXhAFakxSyX4mn0c8XmzHEA1XPgOvWerWhIZEPUkKZTLlvjphU+kEFnFnJMPb9QCmXpCFUPJLZQVLKaR1WL8TWGTN6Kqzry7YwEzVTAUmYAKUR4nU6smryZStBcPy4lWSgcoj2QaEntY3U19VArRUV5GqaASiukct+dKYa6t7OXhaAjulTG8XOGMX72spVmlKhWPT37WeB8H4Ylwsa0qT2NtJXRicgmIrKeuXyzwrJqiPEOGUoi67Ca9bFOmp2Le9bz2PJ8FxPZyn6Xsdf/oxrWoZkFg4ZyL4hLNh/8e67oR59maxT2yBqh7T3TVzMtmVfxXHaIyBmUsgdtQPIyeYXKC/ZwLRqKzk4DR7bcmDCbqJxzIytODz0vFJ55zFC1F81nNb3lfiZfSk0GClaLSnzmB2aict0oDz/VdjA7yygMoRKruXkMVJU4HthSYZFgvK2VqMJOFEAC6XBq0HKqjGL20reUwnVQQLfpCQhgYdrTbacvmt70JYmYNgSlrDlzmU7MZeQAAIABJREFUJNBo2FFl0AIWNVxX1qZr/Y5sSdf1eiujGIl3w5g8L1WzmkX6UWcjZjIP5tXNWzmLgh6C3HcpNsXZGgYDWoSMHbkXjT+s9Wo4i2eIECFHfDZvXFuESMy9utPqjZBXKQ8Ey7ultIT1aLKWhgjrzIDykgyeE8OiqzVeoG7ZVaC1tluaewLDUkynhrTWhgBPY/w9ynvxEiINMg6LzxCmB23k6uudCvU0XaozbQl49T6l4kTVg1jtXR6sum41dS4H4loYW52nMjPhNVh6XZPnrrLtU6+ainUeaG+Aj/AeNKS3Rcy1KJGglTqLo8gtfhPXDTAk0dqH47QXlgRQWURMX26g/qiN9uqeo+kPl6gg29MVy9ayUqIStxDjC5F2nTC/uQKIcHoCDmhAr0ICCVJoQt1pWmk6xZipmSHgDfRiFgAMIRCbCcwDx9CxIMZ1GxZj6bkqnbpJDagwqmJ+403zLd1bKcQ19elA3sgthZMXy8idR+Xtmyn2LmHPYb6OBL2keIUX6No9Q3lO+5L10h8popovoRDHEjyUUCVdFqsOVLl+oPmGvYXkSsHLiAwegJg+/s7UbdJ8aXDzKulPmreitVx2fVdezt6trjNcBCZTs17ejpPm5429FKgaCr1fgh3NkNU4plBh30Urx6m37EoWvQFgLGHYSnN5AY61VqMGFNfFzjW2Tx6HQqZIbXviLooI4JGynVNxwK0neSWYqawW3PNiZADegrglpZcZIKKERhOVokfBsh7CLNzxnN6M21jdUC6jyoez2EQCJyKj0n36d/0cWQgj70LofuIgqHLz4bVWWcmJ6nyNbEy57J0SfszwcK6Tg1XISDHnwCulSgF6wqo+1e6vYY3CnLte4YoG3urSZiAEW+hz3ZNaTKD7PNfzuM4a9iPBlELQ+et8mxiIZ/tIV0ZWDmS06+C+3UvJtErnZbyNEDzVUMj6O4W8GQjeUeHMMhSNnDlnDa1Zr0IU44KK+XG5G1VnqHtLZcbX/WmGqXjZHXltxEG6SrEpUxP1HrrgqDIBUubnrTzq1mK2p+X51bqAakq82y2zEdEf4inc2uuY4jnypJQ9vbCbeZlg09/0xCWUaKiqSylgCbc6Wh0PC+rdlxmoxwivSlkTeV/iC90360lzYmsa/GEIF+9wyylSslJlN6jtUdZLMaZirIb47pUbe6CVGqfn0N70eeivewv251+Ntm0Y10fgUx/D+O33Ax/9AI7HRxZwUesu7m0h5aVIhof5lEWVdVczFnJfhoP/3qw6ZHeTBxDZEnkwYhhlH/CyNT2OUKL7c6/GPJ7Br5cMxaSgRGizuuwmPQyeY4KwXtcxNlSqb8VXBATL+hyu81mo4+CouvLqlGKUogdusx0nhmryCFqris9UPHShhwM+a/pW/9yvx/zIL2LePw2hGCxb5s3lAuVyNN3pFRg+gMt9emFKr2qtGkgrADiEv9KDK2htNAwRfyOxHbMlXic9ewMwLcMVXcCTBXFdmayK71egXpmMjVkPeRe+0Mu9UrjR81EKt0BoKc0lm8GDXhURYAvN4zP6XpNQoDyLBKDNYE21FC29zl2eCtS8FmHWelEUIE8ReQfOCMVrGwx2nSpyYh09yu0Xo4ppDFWnv46gK0WCVCT6TXvjF+D8B/4o7DWvxfzw+zA/+gG0j70f18sjbDsBL7wOd1/5HfDXfwZOH/8gHn/u3fD3//0gktKfiIPNpitqcjH4dUbo4gvSbcthKhadbuhf8g24vufHYWD1o1V8ve5GfSrByDWUNtrBDfbG34fnvv3PYDx+Ag8/8JcwdDU5KrW79roIwRdjhQJaLapSohXbCq/IwcpLyKFu1kL/Q+gVy0txFS09J3wpVpelXG9hk/u+hpcCJt3LTcb5Rdx9w5/Gs//159NDWQ4vIxPF+Kfn34j+bX8BZo6n7/qP0R8+vcyToNeDyrqE4IVFXKskVaNyjbgr6aIz0h6aBfg9+3PYP+vtePyNn2V2gsJ2K6c3Lr14Zs4yiqpwBUrR6uzRKs24ckANOma4/7nfCH//TzBsqgE3hspEBc0Zgns1ssErnEz8yArINADeX43n3vkv4tlPfm+E31yoY0nbAotxLUWhvetciubx700f0E3nW4vMAiayUcZADwMVp2sCFhDhyBUeFZfheRWx3vkvYfuSd+Dyf34frh94HzqCKYQMq6X8asBAg7/0Ntx97R9B+4Z/Hg/v/h+Bj34Ee4sS9NVzkLXQ3upS2ttUaqwbecBAw/Y1/yyOX/3xxFRmqgawAlFKu/7fkxmV9gS2L/82PL77e9Df/i9g/8zPAf7h+zC86kni0C3BQMXICmXoFCUarRSnY7X48cbTP/XnsL/5TXj6v/3lsOLL2tSfoXBHjKwliPHHRNYVGBVVZKHYAj+jcUgKoZnOI6y9cvkAi9C+7rtg89PA/X16fuuMSf1N1Yb+eX8Q41d+EANvxN0XfDWOX/qxBP1OjE/dAWvBE/cc2BI9M8GxuibAUV7XRFUFA+C1mBIqh51fRP+CbwR+/WcBC89hoJTCdXgKG3V1XnTVG+AzKkuFoRgq5IuKXU+jtvKdBuQ4s4mtGU5f8p24fuj/Atj2vabF3WId8sY831/7Em90MLULZFjYDLDteeD8PI2EBvY6vbBScBpoDD5LekCKY+/APILfFY425VSvVB/PGCSbAfdzZhwvgOeeKcDVOj5j3JezByyyC/sXfhP2z38rHr/vPwE++N7shJPQD3f08/PYv/3Pwl75Ssw5gY/8Gi5//Xtw/2M/hPM/9+/juXd8BV3qajLT5b5yR4/FNVVvRf5O3oCXpYLN3I8KwjSuzuil3I8omhLWoWsNAhdxDDT017+Ex4/8Fq6/+2HghTekAOYYP6u6/yyWscWraCtG41lABq8iHjiwv/lLsb1i4PFXfhHb27600pkoXEmudM6b4F6V7hOKDpRLr+sfn13LxN5fZ8bNes/9VeoUGZ48vvSV6K9/E/zZ76TrHHGuGFuAaAlPf8Pn4frhX4N/8sNoz78xAce8i4QGSlO2NcMibnHXOcVKVprv9DZVF6QxgMLEDo85bpPnHKB14CJS4NfheLh6/sxRmJEjBHvOwBQuxDoUDvbGsn8ZBq2HgKTAfbn2c5Z3snorayOeBHT1eMQbcwL2mi/G3Zd8OwzRz5L4Tdvh40gluHpC06sa9F6MD8f9hfs69Nn4GaBkQXywZV3AwoCyEmqokvY8vNzE0OjlMgo4UqffdKB93T+Nh3d9L3AMWr1cH+Okhu2f+W7Yx34F9ulPoxtne5rDPvTLuH7/X4a/80/i9LYvTmQ+L+OBsJECrDSgViZGiDGgEAbovI1ZVl2f05QgR93OvabAxKBXmulhO8wOGJXrruoc3GIrgYSXkpASEVsI+Dx3W86xCLE1YPvcr8Z470/BPv0x2PMv5lnIq1J4IGUZY9ci7aZ08DotSWBcTsdOi1LZKg0OVtPZWnI82hPcff0fx8Pf+QHg4Sk09HWSkQeZSaFSTo5+8irY/SfS9dZdp5qpqaE0EjLtU3d/pKGx27qXnCzvKrmu5+zNsPUO98EjtaI5ykMQqCxFlVcSTM86hxw+w3NXn4cMiNajIbtSDLFeek5W4wDOu6WntDhkWafUifM0IA2NGeD9Fbh7559Bf91XYnvD57CmgxjF+QS/HnwOvYuh6sxFzhcvQkp5a3F+2u91IBX6mMCmQcSdViCYdmm/RcX+HREX92Toqgo8ZoQpbS7x45Md/olPViYD6hYMRbO/+ffjdPcUz37mb+cBqvagARhPfwf4a/8FTn/8u7H/1n+A4/4xOkfNYATYLjPKv5uVV+GQVQ8/07C6amyncpY4WwFDuhYOKOEWgbTunf8+tjvYuI9Tv3sBl4++J/PWvjwDqNp/d8TcjvXCnFkptwAhxXDAkz2E/fz6z8DT9/w1bC+9Adu8UkEE4fZuGBQA/XxNqYpWmtOgbE/Q3FKpNHpUCkn1J1PeBFccQP/qP4n5D96F+ewe4/KMGav5slR2CU9rwPAGnIIDtycvYDx8Mt8h/hBIKYxKTXePh5eQ8mzkeVWVboSHmgEBnY07WuuYtLaTxkAhkwrBFH4IaG1W9TjFm571F+68sNkK2zNUH4Xu63ALQVZdhBRvDMUNJX/ibIrrcDw5tfz8/ZUp98/7wzh/7j8Byjhsfx7t+Rcx91egfdWfxfbs4xVC7c+jPf8q9Oeex3j26eQDDWpWvcnd1nKdK06hu3UUngZfBQKzNcC6IbspW7r6mp4TC1SLeAMxCndmLcRUyHtAoo7BgdmAvaNfDjQznKxa1w1Ae/s/iesv/kgSQodptMATQP/4B3D8f38X9uXfiOMn352xqYqfTlZZi8ML5RcDddTU7enAaasgUHhFN7u5DNqs5nnKM7g/HK/YIk9xONC254DxNIq2XvdmjF/7SIHAdosLaHpT/vFb8FDly+GJVPwojwd3z6PdfxzbCy9ifup9UQx1eh6zOXB5WsCfAQPVbm9221ZuBnTn/gC0t3wFTm98PY5feHdmtXJojJUQRRcxaffS78f5za/H/Q/9VfSXvhI2HvjexV0GPQN6CscErG1oOAB3bK/5DMyP/0J6LTorUNltUPrPcr7GOrjmJHC7WSkXYkU+w6jlTXET2LcN3cKzSKyhlaKp5rBKQ8e1A44nJ0sBX+N9hy/3z5ZBVbe0JnxLCaWg84xyqphV6b5Z9ZJowHEzYP6jn8fjR34K83qJlPzv+1Pwf/CD8P5m9PMjHn71x+I8uqG99h24e9uXYTz7dHpg06vYqi3rcSpM7SPDW6uwUiBnIw3cUd2OkUKLLz2MiNnVESo3+irBduWAWZvhUY5tiG7Tx1/+OZy+6TtxeDz3YVQx1NUBvOmz8fj+92Iwjjw8YqdDz3XH1YH7X/wR9C/8WoBZhcMDTG2oasJUarMORfUBapM2i7Sw+bgpQjMUxmGIas3oDg3360p3VpcqDXdgu8O8PuLwDe1VL+DhYx/Ltag7UsIQ8yRUax/e0CNrG2KvjgeOe7/yHJQifDgA3wBcB+w1nwH/nQ8A1nD61j+HJ9/672D2VjUaHpZqa5ZDhoMfq3hH1hSnF3D3Tf8Krr/202lN3cF1xLyJwVDFQLe8P4fzN/wpfPpH/3scx8ThHeO4BAZAQwAKlJ6hGpmJaGh4PBz++s/B9SPvyzO48J2aon2dtQ79uY6lk5Xh5UHsQRmJZsb28SWEMeDwDvOjhh+TzmOh/2XEfS6Xw3P9Wxf2UdkHTcHWWU0q38uxdIjC+bt4zpyBhTwegMbiqRP1GJ78Noi13F+XO3ZOr8WTd/7rOH/Fn8A8HmHzEe2512J84gOw0wvwZx+FH4/ofsHmFzQ02HiQTWJ6tzJFEQLWFDUAeLhOjv6vGqOkOR80J6wl2Gb5czwOT23vRS9q/gINwxrHru6aLiYqYA8/9b+gv/gOPPcv/7vY3vCWTEEZAGsntFds2J4+xWa6mb1u1Do15AXId08/DOwv4rlTQwdwbi3LsOVpKI5UbcFGJbHOXDQAG5PHGTdzX8NVsHWbdl3njg7XzFHDbDt8DJxf9zb4J96Hzu+1J6/Bk7e/E/srX8LdF3114ivV+htMvbdo/9+sbmcHQtDP1PbdovirNcfWOtprXo/9Ex+FwWG/8yHg0x8GxsyUrDwDSYBG3AeuU12K04H20hdhfOjn4Z/6JNzr4uMC1VRwxKYxd/Sv+S4c7/k/cP3dfwyD4bQFcCgh1l2wG/8XljieBQv0dju/Cv3OgU9/MpW5Lu89bZaTuJ7sDVszPNk5zpDDYjQlHCicQfiGzkEj55yC3NuGOQ42TBk0XWswJLvy54k5zRV4jjPbm+XPT5tmk8gjcf7M2FOjoi9U/UND9ttsLeZLiFT7snft+bzFs/p8Bjw+Az7xDzkd3mDnF2CXp7AX3gL71G/lpCwzYNvOGNeHBFb7su44s6BHhMTL5UuLwdGah+5vZejSdIXecJVyC/UOCzhRWQGhyeB/LxQcCaqQYD2k+SPmD/4lzF/6WdiLb8CpVRESnns98PAxXEfNsgCQ1WeHI2/7uswBPyYuchM9tN+FFkBxsWLLDAdQ1lzrm9YSDOyod0s56J6Uy1BFYwmY6jfuD0fbOmxObG//Boz3/ESCmEc7ob/yRWynO/RXvjpBuf351+PuD/3pROakwOR1lDIury28qAkfDXj+jbDjY3h8OMJS/dT/hIe/9X3sQVkAVKhGwTN7I6GVd9gNmJ/4ELa3fBn8/CS9PVU0CqRTpmU60N/6B7C90nH/yz+ZQgKfaPsTnF73Vmxv/Uqcv+gb0VvhCQ5mSMxiipo72md9DY7f/GlmEwrtX7tYZdWUuYg6mljPhd6I6KlBNe30Ak5f86+i7TutOZUFALQOnxWGXF8mJGN7NdpnfxUuozxaCZiKmB6Opa8CJeS6HjAEUyGRp2croBdArunxWnNKRHOI5l50cAd8POD+p/4rPPvld2eGx3sL3nv1a3D93Y8CqMzaaCdgXCjwVZUrHGjMzG5wf47rUTQvXkd6iddBQ6Qyom7Im8NkleRtWCuXThVz4VoWcas4SqWrzI/PCfv7P5lpU/fwAvpbPh/zw+/LGBSojlIJ+9UFNJ1gG9DmJMYAuDWYz1R0YwLn7sArX8Jx6hgf/RAgZkIJiTgk52u0hm6ev9+4P0d1QgLICVXGZ7TeAHuC9taXMP+fv5oVm/uzf4Tx/7479v4LH8yCsdPX/gm0z3obzm/8mzg+8hGoC/euFyhb8z9D1KJN24HrFfsX/wEcv/Fzhc28+FkYDx/D5enTsFhQKGUYBBsVTo6JHKn3RAj+pz6Ix5/+YTz/x/5zXH/j72B88D3AJz+C+eyTwLjEfRwGtO2E9tq34e5bvgvH3/0hvOLr/zX0V70EPP862N0r0U4bZnsR7enHgE9+KC44mhxf6JWtaM1gbji//Rtw/6P/WSqUx9mwv/oNmJ/4CCLjZOkJOeqahuzWRHiMc6KurYDD3/5HYW/+Uhy/+X8DH34fHDPxKG8dRiAx+isaevNMV2+v+0Kcv/w74L/5cwHm0sXQiH5rBhs1dd3Avo0nrwMun8TpuKT3GYJr6cI7UKAr13u3E9C2uNFPQusA5+E2uM/ESE4vfSEeP/ZeNMys9sVzb4U/ez/GMZiNCUBybxv8OKDRhsdwPNlbrk/Zl0nL0pvBW/Gf6WdgndTyu80BU7l3pC4LNAqw13BORcEvAnCzm9mP0ozrpTerlWwWYFNea/e5X4bx638zP69UfzNWSKJKkO2lL4B/4jeB6fD9eezf9m+hveFNgAGP7/ovYR96fzDX/irc/bG/CNsOPH7vv4fx5PXYv/3fxP7x92L86P9MgQ7uO9Bx/tZ/G+2zPx/zt38V44f/u8jnn5/H9p3/IfDCq3D52/8D7H2/FIdsyGv75Mr0t30dxo//N3CO/rftDqfv/At4/N//U8ztVehf+vXwn/nh2NjlKdoLL+H07f8RzgY8fv+fhz9c0vPROdY9r4a7L/oW9K/6Nvj+BPaOP4jLD/z5tMbtS78T9hvvgv/m++q77/gjePJV34r5j/8e7v/Gf53PVYu8cIkJNpH9+k/g8sGfRX/rV6B95pejv/olzLsX0Led9HTYkxeB3TD/3t9CuzzF8dvvxeU9H4V/6mPYXnwb9q/6Qzh+5L8N3ji9Gnd/+Lvx9F3fg/HCZ+L8mZ+N+1/5iQjbzGCv+QLgfe9Cv39KZQw8+dp/A3df/E48/Rt/Efjoh2Cf/804v/QmPP7M9wPHxPb534L/n603D7btvOoDf+v79j7n3vuepifJmi1ZkgdZniRZErbxKPCI2wk2YNNxgBSpIqE7kK6mu5oEQhdUupymuitJpemhAnS3gThOt8EG0vFEPCbYGDcasC3ZlmxZ8zy8d+85e+9v9R9r/db6zqNvlfTeu/fcPXxr/q2pXHAZjr70u5DtkbfwF+zf8gsYzr8U7WsfwXTrpzC0Q5Rj5+PgtT9neNsf/iLk8BmvoxCgNSzD2dh/038BOX422l0fw3z7JwzYHSvK8QsxrCqwXWI+xHDiaqxv+ilgtQc9egybP/l1zJut/fzMq3Fwy3+J9tB/xOHnfwvljEsxXvt2HH3z4yiP3wM547nYf8nbMd/3BUz33hYDb+y9BetX/C2Ml78cevJ7OPXp/948aqyw97r/CnLWhZi+9nvY3vVFQAT1up8G/v0vYd5szKPbHGF8/i1Y7v1CKLVRvf+pjsCyxaoWbF3BEcuK/b8lS7/Z7CcAhgGRRk9FzcFHTQeribDMBtOWDYDO8JkRBiZuGjtQEx/oXd9ta5HqaqqoqwOsXvujKFe+GCoCffIBtDv/DMvX/xSl7KM+7wqc+sTXsUbuQx08Pbnyl6oWnWN18zuBv/gYAMH49r+H5VufxPajX0I5fi6W5Sjy3Puv/Gtot30Uw8vehiYDxnf+PPDVD6G++qcwl38FaYo6DFYheMO7IcsDOPzf/jn2/uavYxpGtKMt5MVvwXTvFzF9617s3/waHN75F1hQMTznYiwP3+vWQlFRoCfvx+FXPwc0QETRrvw+rJ78FpapoZ59EeSCS6Jp7Ohzv4Vy+bU4/Nf/Ndbv+G+BvRX0aGvEPucS6PIscPKpAN7Wz3sNyouvx+G/+SXsveLHgEtOoD39THiB9YwTOHr2qYg/y/75OLjh9Tj63Z/D6j2/jmG9ArZbtBNXYHnyu+CKPIKZ9GDmzSmUu76Adufnd0DQUgC96DocvOH9OPXRD6A9/qArc6+bEMH22Wdx5vpYhAj71/4glgdvM2Nx1pXQs8+NmL9IBWSLZ7/0+xhd347nXInxwvOw+caXMB6cCb3yGoxXvwRtu8Zw0ZXAwTUYrn4hpkcex3D1TZju+Kwx/CWvguijePojv4kz3vF3Mdz+abTbP4zlsusx/ftfRb3hZ1GOHcd88hnDCNZroClWr/lZtDv/bxx99zs49kM/j+1ffNxqQa56E+aH74W84HXQ2z9t+M36Aoyv/hmc+sw/wfLkQ8CZl0K2k4OXwP71fwNHX/ltDFfejKUex/7r/z6mOz+BvZe+Cyc//3/gjB/4BWz//INYX/fjOPruf4NpUqxGk8Z6xZtRjwOnPvpz2Hvjr2J15lnYPPkk1pe/Fnp4Nw6/9L9j/zU/ju03vwhoBcY1yjL5oBpgdfIh1Kteis2Xf8P7X4C2Phe1TqjDAG0nAwQujlOxPWLxmDPxpDRS6sDnUDNUoXJZGlDCUiGt2+CexNhZIhazjJIFMYENiP2LueUqgvHNPwOdH8XR//nL2P7mL2L67B+gnv1c7P3UB7D347+I5f/9GMpMt8o8CyqaWTOcqS9+M+Rgg6Nv3A7ZPx/DiTXKX34ZIgWrH/kF1M0pSxEOa5RrbsL89T/HsjToNW+FPHEbtnfeAdQWYRAuvwGyOobxmpfh6LO/j/Elb4M+8x2U7RbDuIfhhreiPfgdrF/6RkzfudVCixe+CavrXhcTrYwIAr3nq2jTbLMxtWD/hndgc/ethhUcOwfD5iRYdSoXvhxl8yBkO6GesY928ijKz+ubfw66v2/ZkOZt1de9DdtP/y9op05i2jsD+uQDAXqWg/NRnnsNyjx52CZY3fBu6DMPop11NdCeRNtO0LqP9dv+PnQogeQL+uxB1lQMHn8Pxdz2+vIfwbHXvgfbP/41lCcfQr9HJGh+9Bh07xzzKAUoF74Qm7u/CgWwPusEcPRsAGvDpTdCn/gm5ORTQfPykndh+fongLqHJiusrn8btp/5X6GnnoKuzsX4iluw/ZN/ATn5BKo0DwEr9m54D5ZH7sbeC9+I5X5XTieuheBxbJ55BvX4WWinnnYsRlCe/4MoZ78ABY/i6J6vYf+V78X221+w7MmZl2E4cQZOfuqfYnzB2/0FBavr3ge973PA0w9DzrwKx65/O+Bhr5z1fAz7gs0jj0HaBnsvey+2d/0Btvd9DbUUrF/xfhzd8a9w+J3bACym3AtQr7gFMhSsr3kDDv/0dyAXvxp1PMTmqacAqVhf80NYHrsH9XlvgD5ymwH9F16Hur+HAvUaiIJy3lWYH/gqpC3YzoZv7F3/tzGc9RwsJx/B8vSD2cjIjNHS0dxJyUVRQ03cCN3P6GWIG5FSBUrMgI1J/fLdodiwG4I5DEWqAFvNMup9B7JW1TyEesbZkHv/EmW7QdUZ+vC3sfzFnwBPPgk99Tjqy38I65vfjLJ/gCqCY9VLxD3WruvjGF73ExhvuBHzH/xPVr++fwZw+LQppYtfgXLZC1HOPGbZlFf/p5Bv/jvoqQkY1th/1Q9g/tzvo5YSy4WW/fMxvu6HIee/AMv37sD6vb+KeuIAyx/+BoCC4fU/DcxPY/WDfxfQh4HbvojV/tlYv/rtmP/DH1hR1mn1EJaRKdi/6b0YL70cdTmFVSkYn38jcMZ5BnyOBzh44/swfe53nAAFBVZctr7xx1CfuBX10QdtEzrMssvxA+DZpzCedTHGSy6DXPwKoBYoCsr3/yTQjoBhMEDxopdgeO7zgHNfiL1b3o/tx/+F1VG88scxfe0PsWxsrXM967kYXvQqDLVEQ9JQ0/WUUjFecROOvfsfY33mgM1HfgX69OOhJFg81tQ4cb8cAbqP9bqashlWqLpBkYLh8hsgZ5xn8freuVjd9NcBbZHtGq94Ldbn7UO/9WXU8QCra96G+RsfQzs6BQxrrF72Lix3/F9oh4eQcR9tOrQajBf/dZS6xfrlP4rhgvPQvvpRaFljffP7sPnSBy1FWAZI8zLEq96O+pyLUS55GfSxB3Hwjl+GPnk79I5PQOo+Vt//d7D5ygdR5meAtsa4Kti77CasX3Az9PBJtKbYu/r1KOdeZRZc1jj2qp/E9JXfxrg+gKxOYLjoMrRvfh7DuAaOXYi9i56D6a4votY9SNsYDnBwAfZe+hbIwWUoT3wNx275ZexdeiW2n/kfAAXW174XMixYvfz9GM/EnCYMAAAgAElEQVQ5wOaOj0OGA4wv/xHoPEMdIB6vegfK4bcwnHgJyv5xiAjWl7waw8GC5aFvYr7/i5ge+LoZR+WcFcusMK3MrW+90a/FskgcIgU3CASEAchARoj0nccvjG+aKjZReyFQFXD/B0epUYFw/mMVYPr4v8T4134W63YEPTrEcOwERI+w+fyHUb51G3BwDsp1b8H6b/wasHka7ZF7UZ99CqWO0HMvw3DeBdje+knMv/tB6GI1iuWp+9AOLsXqlvdDnvcKbD/9YQw/9POQp56FrhtOfeS3gdWF2LvgCix/8j8Dh0eGUTz+NNY/+JMol70M0+d/F6t3/meYb/8sVpffADz1CFbPuwF67S1oT96F5V//DoYf+2Xg0QehV78aw80/DP3ib2F++tno3RjcZQO82Oim92G49EJsP/rPML7qJ1Bf8Ch0vQDjZRjf+DcxPufFmG/7CJaH7rMw79u3Y3zrf442FZR9wfZj/9QFMCcwT/d/F6s3/W3gnKswf+Y3gAtfheHtP4+6rKGn7sX02a9h9X3vg97zNcgr3oJTf/QBlBe9C+M5I4Zznov68vcAZ66x/eNPJVB9+BjKJe/B6qVvw/ztL2P/yfshbcG8dw7kOVdj75Jr0B69E9On/0fMjz+YvSrIArbIODF8ffg+1AuvQLvvbsz3fBnja/4O6kahz96FevH3Ye/7gHrpdZi/8kEM195insxVt2D9ijfh5L/9x8DcUMcR5eyzcPjxz/lOzX2Ugz2c+toXUAXYPPwtHNz4DtQLbkY5tsLhH/4jrN/2K2iP3I120XXYu/adWO75BJaH77Ps2d1/hr3X/T20k6eAM87E9Gcfxnj9WzDd/03sXXEjyvYI66teD3nhmzF944+xd+PPYLz2cUh7HPKiH0W56EpsPv7fYfWq92PvjOejnH0e2uNP4Pj3/zTkjCvQvvdJTA98G8NFN6JefB2OPvVLaEtDKfso574AR5/6h1btvDyFJudifd37MFxyPQ7/w2/g2Ns+gFN3fRoHN78U81MPAOe9BPuXvw7QJ/HM//OPcPzNvwI88R0MF9+I4YXvxHT3x6BnXY/h2ncBU8Fw6TWYPvtPMJ94JfZf9w9QHvw66oXX4vCzv2YG/4ofgJz8JqZHvxMeIDehQQ2YrcXa50UM71BF1IKwqU2wW71bikJ+593ff/LyvXJA1LN1MS3dC36PLgmQxVDpzmaqjKmtRQEcPwfDeg9y+DRkcwqcusyehSKC+di5kPMuQTk4A6VN0Mfvx/LY/ZH94Cp5c8HPBi57EZbv3Q499SzKJS8GBqB872s+OKZAr3gZ9Lu3WaIYgK6Po1zxEshD34CePMT4su/H5s8/CTnjfKxf+nroWDHf9adoD9wDCND2T2D1sjcCqwHtG5/H9PB9MeUKsGrFcsn12H/DuyBtxPLQrdAv/Bss0wJccDVkfw9H99yOYXUc6ytegvbYt7E88VBM/F5QUC57CUqZceqeOzD6edv2LQdRyxr63JdifuJeiIcB5ZJr0XSD7ffuxFgq8MI3Yn3ibEy3fwL67NNoKKhXvRrDRc9De+xbmL/xH9HasmMpBEA79hwMl78M4zkXQqWgHT4JPHY3tvfdCUwbOwNapc4gZJt4bg+Ts6/EsA9MD3zbFPOF1wKYgAe/gXJwAqtLXojpoa9jbBXyn/xDtMceAvAMjj7zL9GODi0deeJ5wPI02lOPQQpQL70R8+YRzA/ek/e54FqgAvP9d5jFHI9h/5pboPvHsXzvy9jef5e/nzFqueAa6FCAB/4ScnAhhvMvwObuP0c5cTXWV96ENp/E9K3PQ599HOXgXJQrX4NycCaWR76B+btfQVsW7J17BdrxE1juvxWtFYyXvhzLs/ejPH2/DbdZ7UPPuwLzg8Z7bTgb6+ffBLnrk9E4Nhw7D+U5V2N68HZgcwqrF70Vz9zxRxj3z8Z45RtQ9/cx3fcV6CN3mczU46hXvhF1/xjafX8KfexuTLKH8QVvRZUjHN35KawwW2h7/GKUsy/B/NCt0O2R9dBc8mq0k/dgefI+p1sO+ikCn7HJlLqclsLNalZmQObFUsbfe6Idyofe89qTF63lwAay5GANAmFAhh1MX/EGXB6k8J2nYtfoh/umO5Nl5Nyv2ZSDRrKyjp+ne9QDqVRE4ofAUXjS/c7c7IW5lYzj6ZjxYYENqw15MKzFsP988G5nUVdFcnCsAMtF1+PMn/gVbP/tB9Bu/cL/7/M3ZeFQt09COI/DP8MDjmfJdGEHEwRhOQ909GzV0Cl5IPsqxM+CnYwxrs2BzYYcTcfUJvtU+EhFsLM/FumSmlWqWXhVxH7O+hDpzrYAaOvzsP+3fhPTbb+H+Qu/F7Mb+Kzxrk5081wkDAvpTPru0ly92azrRfHeBlWfqD4gyqrTMDqO5bgcVxayrHkc4Eum7SlZgzDWLCfnM5NXeX0WYpGOPCMOynGM2ORHEM/en0MBRwhwaxpXIIjzlxtcZjnE+2aGXVmI1Kzm0JumzIQgOl8VbO5DpGjVr/PgU+2wkDEbMrMhSCDT/u6VY64A7DOCdSkYitUKJHiSewrI5DFhig8kWWpd6DHIbm0HSURMhM85SI72W5WYDxiCvschIErvRqMyk3MaJs1ZmlNLV7sg08ck1lgkZniyboHYTPv2l7C6/oeh63V2XSqimo6VhfDnYNs2n5UdhVEJKHx2+Hkhcu9Arnik4otiOGTlKn+Px8iReQpjJCCLkZTPKxl68vdGV7jSMbEAvllNfPS+g72SmTQgDQuQiHstQHv06yjPeSWGE+fvdDrGPgz/H9/bFLUpRlZ2jq4AqGiaAntjSWEFMSUrJqLiYhsAz8TOWHLOhDOeQEIJ0nACEr1SK4/rwwMHoodGgGgkAxBFZpayTt4vwntIyBjfuTWOebB3XA15b9KKNKyOI8J/j2p+uyStt94LkCnUlCcgK2ZFuvYIf16I4RfcwFZmVex5UU8ytl1okCyNPVp0Z/r12uukY3aAIno8NK6RVWRb/8bRkhvGqqSXUrAbvpCR2bMxuaZjr8rUPYuh/BJpOh9jEpaNAkgFNUrGZetgkkwjDZ2C43s3twgEYGcFlie+g82tX8J4wy2xOY2CxcnO25YVcRvvA+A5Q9OLU7fwfC/uUoUruugrWWibcmJ43+PA/xMN53vSknD717pjDNJchFWJ9vmjpcUWMf6O0dyqLWmx/irN7fvcgnW0mOBi+xSmL30Y9Yb3mGBJVlOyrT16b5CZobkh+kfsSKyPAeSJ1k2Cd0VItceyfo5+FDEgj1+keQ2Fbb0SLIVWNQ+FG+RjHoZ7C6w05bmoZm+QwnpNOFKR5Im0peZZAVxnKMHTvPZ2yY11rHzl7+R7d3NgiX25J8pW+fVIxZB4JJCt7E2tXyWeQzXOamlAWRd7Da6qV3/pSRWbpjhcmlUMSnoEiwLPzlkCzh0YdNmkexD4i5N5VzUzHv1sAbqaqqmFuRWMDL9tGu6aAr7wyJ6hVzQUOIZIBGt5sLRa7LCscXj2u5vFBp2y1Hh0rTM1axDi8BRVxfbWf4d69eu8c1RcUaSAqWarOPtAQEFpuw169AgYKoV34P/m4mcqRZ5RCJSXqFPRFb8nv8JrqCnUOzRfzCiwQWrovIamimenlvMtnOZUanzfpHk+37pKzAZp9/8ZcMbVWFbrHSGiYmuaS5UpHAwbVOHNVvnMvWABPXaGKLvmFztNuR3NWgvsvTezvfeRb1Ub3Y2cFsVmMgHivVwesZm9L6fzXEjzxUvAB3otksqRJeVhwUlzNipBY3pXNrFpKCOW4M/NnpvDpRVeaUkXuCP66IwQoY4C09y9+9RcuSBqMloDTm5aNM4VVXvc2lnTGMQCS5tGHApko5PQTQfWtXR4Rn52ccUydszCxh0AEQszVUv3iNciQ7fu+739ZBUtBbGgt5SKo6XFQqDiyolNTyQU00h046lY1o4a76RIq0SYU6AYSsE4P4V2coacdZa5tv4fW/oHVst1VlOQFo+KtUg28/GcGhArDyI+DQMlcR4xOMZffrPYJLCh5CDmIhmbQjtMonQ097CI+zyoYEljps/HIsEjQFpJAbuQDcQeHMhYGhW4QNuM+b5vYrzoyvDmxPmPgrM0xJTzUPCOj/UeBGtDyAdL863p7Bfxd4tskPMY/21DfFMxrN3lJzYxVAsD1t4dySa2zBSmW2+T2jM84DBg9pnQCEQ7g+Zn+WxsuiPu0VryNwWCA4IYgvA8Nt7lylEHppy8w9ifkZ4sca61N+sVhtUtn4upVsuEmLIps7KpSWMiNkUyeyHS6vbj7Kih1N3tKuni8wAGt6DbJX+Ptsg0L8LF55dIAov8oiKgy9uQigRIz6J13xMgGuHocXDZ8LZ5KNGshZjvyv8WV2JAeiuCXDDLPXFTUyyPPoT1eRck8wuCKbYeelCYere4t8YsmKLwUplR0BclE2sITwM7J7OgrXPosvVZ6b7aYuV+1CCxHJ4XPQY4Q3P0Xuz87BQavUHz/rpR+8XmoHBilwLQZihLLQCe+B5w9sX+rBrvG/MSYIqPGNiG496gYVWhGaawKU+RE7O28b4aIYWFc+nNcS+L+Mv3y464doDeTUEas8np0I/B47wQfn47Z+jQ3HCwjok0ZJXk0CkME1afC9PgbePpWdGL3FmCjKTfdslWc4YsHHgUct55gwCH8di/FInpLK4N7blUBwIsVAiCFFKGBTEaHY4NIAWzB7cUCPQ6lUKCaJXMJIjZlgQ1F8AncSVQypH9zCIU15yLpnvNkfTc31mdeSFWLs7PAHaPVdmd5kT3v2l6KmzKiuEo0oNdLvSbDbBe20suW9RxDQTyjADg1N8RkkAe3eBaBMuSey/ts0BzJcphPvxqyDkN6mGKSoaQDIMIWPIcFfZ5yvogqaQaMoY1mnP+pYTLW4SLaRALkRbHiTjpiQIZ58N42IWoYAbKaFmKNkGHdSgEZg7MQOS0KxH45joOwbFzWtU+a6c7g3akMAwRP2uNIU5cNhQ092wB+ZBZs1wkvDu93hb1SDB2CeH3bBNSoP/KLNKW5dfLstudXWt64Ev/uwCadF5jyS5iyqphLQLh74jGFDlOZ6Yn0lw5k9aqdpPiCqwvn6gFmGYjgm9el4EWVMGDcc2LXttrMDIXI/cuM+PpQdj8lUIhxTrrGEtSOcxu3W1cl00XokKilaiS+IMuuSGL1mDS9EBEEBOS4tHIgEo32cEwmAZeVwmLSOXDjWsRGoFAbFpZASDPPgyceaHFeOdcgOnOR0NQ0D1nIN5i78732S6Ksbt2YgPp2Si451PinYFdz4mMTpDK3kdCIVCZiHZYT2Pqz/p+eOaxo4UKBhpeAmd3gmft6claObU8hUJKZs8UHiK2I2jZxwRBPX4h5OnbwxgBHnrAlCPnS1jKOa8t6Mbi79AccSC9YDS1Z2EYsJ3dG/Az7hUKXEFCTCFyEztBfXpNQ4GNYyzpGVCp8Tk5kZyhEj3LbVOMEHDqFzOHbbHvsQyf+0b6MCPLEJJuLMluagaS+2OV56mZgbSeDyuqFElFq438mqFnKYmtDNXlT1UHABIZCUmtQ+GOHZzowpKOaQWw7ekKzLCmMMbsMXhU3CPpXFxiBNILDJivz10L4gzL/R78DGdvcH8EFZ1qhjtcN89Bq9tG5eFzKjSVAZAt8cysLHBLQSPQaXVsHodO+6g3/zDkzAH6yEM5WUjcMoNLmzItC/dsuOpeO++Bi41sRkLuF7W9oAUcSDw3Q6mbK3XGt9xl2YOekHzufqUhH5XAmNFcdhQHAW0niQm12u4RLgJGSy9ibon50Itc4EyvM/DIfTh2849ieO5LMf3Rh+L+Ejzh3o97XaEoxcJbgoi1AG1xYFo6A+Me2+JueHVBpeAvSnwlsSpO4IK4O99yqhi/KEgQ+CRtCfd7WjJ0Jxawql7M5JjBCGBaJMoR6LmZkSL4nouiGT7VCtvz4iBn0FxdMfiLi+RcW1M43F3aec2SGRQOxKEoB81D+efoy5BzEanvfvHl/+CgyCjovQn7k24wc8M9YEQLWGQXWKTgc7x7CAE0hJNCScFQ12yD35jMGdvUYR4KGYrx4X41RcFc8eJUo0WjwLAqLZ7bTRBDKsD2c1RaTM1wid4M342aVwG0796Ocvb5mL/4IZTtEQjw0BOgMgyLrp1XIMmIPFsqaBKwOEAY5+wPMgag7HX+2oHfwvfWULpS0vUu/lCmLCQALb9VWKB+ujaQKVcpWRtAl7+fhSmO1bBOgNZyagp98A7gzAsx3/oRLM88EdOj6CuKexXcOUrMqJ9svTcUmw/iGrb3spLmWdNCgxE2zs8HbskrQwNloxYiPBKnC3ssKORxJpI3FucnPqcZrJxVEp/n+5Tkj57mYYyFU8Sc5kPO0aQh4herMllbQW+WtRW873Ka8eB1Fi/8ogGr/mJBcwFObnSSD73ntaeu2C/73BuSgiGxGo+doH3xTKSfgNiSbszYKxK7WCwdpjfQWVtqVRKcLuSkGq40sxLVX3RBZkeahzicxNwLY29FC3afbW5WKxIhV3fwAJfdcmgumSE/XwQxyYvDasMbElOQmcJNRuDfeU8yx1hMaVohkVuvTtnwPQQZZ5NexJiWZl5QDIsFdio1ySgKVrFi593oZZDZFwqdPzMXQqkraAMXsVOp2DOmT9JzBmdYmszKew0u0NOSadMiGS41ILZ8M+ykImP4wvOP33VDQ+UpYs+/Huiqc8FzDgni7yfNs1SaP6dHQO+tF6ix+IY75yb+DnlR3Tth2M8waIfmwbu5qhIioTTg9Oe5xkrEyuHBkulnf4qm9jDDIBGGh3IreT5LO03OlTQAvvdkOzWMRXQsBgZmvKxBALggqh8Ckddhh2ElUoVUAjZqLJnNB/BHOWnrCk0YVogzhcKuEZOzNJWEgXm2NY2Wf1ZAHPwEsoeBDLdy14qEqGLr6Ydi8TQzFPQAyJwW11LAElvolH9IPwWHDMdCIQoGmZI/U+SoegW6gjcTws1iS3ZZB9IXobU5kfWtu9sscDPmllAkRSRoSaB6qCW8KFUT4H5JsWIXoaeiCTzIz5Ye4uzgHXENCggVWZFM//ZKhVaXrnwVm6jNcA3ILFAVwxxqYUyd1zXlpGg9zQcJhSliv7NXxIcZO58yTu/4C06XpDmXPyW+xZNRcLG1KdCpSXggPIPavXcDukHRnKZl12lq57AePISpTnNXMiz3LgJMUxbYzR5aMwSuFT6hP8u3xQ1IcdmjXPezOVVN4Wjr9umCBVseZgmswo7anTen5u01z7YpVnwYmPZbFYn4lkQrxUfl0XoghYKaGgIHhZKROemaglDRp9ISIBV4ilazYIVCUsQ8Bk4UZwxIwbGDoWuccfLRbO/Gzd9UKozfWTvQe02CRMwbQadCt9Yo0NxKMzxTZz4oooAqtpcj5zrmsuBuHSI6Za45u1McWOH06qnlfpYqHQiMZIxNc0C65VYufg2SNQ/bxd67j3+JnxCXmB2QG2txZWm/2zR5h8pT3JgQq5k17wHZrYkgrUaPc0fny57JZ7fAq2F3Cxj5OLw5F1ZiGFDg1NRsxN2SRo0ZsOb0oeIQBxwh6e22BWH8ipTgcab1B0klXFzLsmeFszCbKsaB+0uMrqUY5pARWpZqc+GV+NyF9eAVn4thHMRq6KGLGJajmsp29vsWMhSyjwawVDUHCpNnxwEYZlXM6mPVBSFExZlydIIw3l0UOLW0qIBkmrSKhpva1MBOeiJ0DQnmjEXw7JzVmEW6TIPfF+rZAygWzT0R4tp+7IUSWRBmRklQwSXK7pJCMM0Na1pM58bDRUPgWVlH646iODmpC6HEWPtSqNzozrdonmOVXbjjagVPXDHYgKj2NLKzRsXnaDbF7EqH1Ys0tCxlZyp41j48MoVRvXO1FutNoNWGn7/4Peem7g06s2l6BxRC1+lG861N8R6qYDu3wJnmJYFQNI0N7nFO/u5jETw7tRC4AtI893HALXEMC3bATTtlLeAGerf8TQ0QdaGSIcvRtVhV8XroirkAr1ZMD6W5YqewnNy2UF7bWSPUYgp3qJL1NmCDmoan2TTDHXpXXJQE9+BZ9s93VxfYaQFqyTDICrkQS4oaw5wwIglwW4o7h/2KAEXNWIuaQuFCbMCzicU+DymY5izEW5rxfi2Gl0wzZBDhli1z7TnK34Z62p9rZyim1vZd/dMVZdqRef5s63HkVzINVfzFuHmr5Efd1TEi0Wpy1L/U9DIACUYbaUFLxqrqYQWBp5U//14XfwvcqygaBCySbmJzq358NHPICc50qwGYdu+emYbAeS8UJCdDi7JSM4cMbReNQjYzeKnMWC0KOAJeOmXDc2q5eX1q5ulVQdQTRB2KezNqGioUDhU8sNs0xoFIVBj7Y4n6gamrE2Bo4pewd0cCxcvCVgAT9r4mh1+xGdwVVTaNZfOUaCq+oXiKvuTmNaYE4cKxHuzZD2ycaAhBdQtvhpmLfLKbughwfGXx7KIWDpA3eA2+N+kkMKyIi45LsW1iVQRN0ksVGB22Cz0WKuu08nsDOqWTGbLNpGH9F7VwA7AzGUUi3JGCqFoOIFS7cxaW0AsGMAS1d2DDmIWzgv2V/R6B9VKCxVNgFZ6ec0m2PafagYvMFSM6MsnWg2s8pvhYV0EGEpARmWIz78MKsFLA3FBY6lAVp+asqCP5BQnuESsBslSdpcmAA5ximRQSTjuXuAg6ZWRg1dw09rmenjbuGYffEGQ6lkAW1+VRQHlvwJiV7zzWzJtTaBdVHHovStzG/9pOe38gwyxId63uOcm0/Yi8/hVsQnoqCTavESCO/RGym3rrXXe6/xQuYjxUCOQDMyLZuGaGJkO7aVGc2uaqRWIIdo1cLkRwPAqZxCw0lR7/I++RbqqZLUiaexs68r13aAzEM/bKzpSVBjYSQu4gJpcc9wqAZzJ6WC8e+i1qS4ZYtdrfK8KKjhH6dv2xJm9FJglpSOHv3Ru1ebEGs6R59p8UKiELIXWYmsqmGbP2FZQKxGb1BOmyfFth3gEcj8ht4zkYFjCGn9S03baxmk69OS3rJ3JPSKa6VAnKJbikcWgSKDy5kABXf7BHXbgTB5zSigUaY/4VCDDV11gmQCd5mATxouALu9kKxqucf8Gvpob7cFWinPYzjoUXUMGK4yiZkeHUI9UMxxbVCPEI7rIk2Sxb4jb8ilBOEttQZDgIdIIoCcCywc2K1MwCbZcu5ew/a41utcYaPHqA05KfK359KgUrzNpdEmTnk17Z0nmtbBZTTZozNl8YryA9AMAU3mrMrAiBTj5/LyjcEkaaF9LcsQVtRi/DCro6DNj32TVK7Ew6L7R197Nz9toc0tyfe1kyncyaoaYWosEVay0Sy5GBlEF6lAyRV7UEH3EOxsxQVRGVoP06g9Hxi0KhrpCos+ChA3TXUxs1Nas7Ci01rVVakRBo/zvdbFZkkkkAxFRvWiOCeQQZAewME6bFZbGVwsA6Q5TVBSEFU5Bgpymb1Nj2HNna21se6d6Hqr0IvOoz3fhA/5GxOp+VJd0KCqLuZEbY/Ibu3jFXgZYAqZQ4e8NwBV+Bt1h3YPRuxPsniBuAJ2NoTVyFtOifu0jWydBwsDGMIRTdd9JJnelptdnMRaaLkDPOJetammb9Qumeofjh9wt/iGcdzdlyAM1x99PiNF+6DJvS883dL1HEhqzpMM8g6yjgmADbtOmtMbNAQWcHqbiQWUlBtqhnvYiEJ9l/rQbDYsjvljVEZEhU7X0Ao/12zhAv0uaqwcdzsx6gmMpdxJvSEqgW5wM+iiC9L3o5tiEtsmqGWYh4mlKS2QqQC31wuhsIT4+6N6HpUk6Osi4whbI443MN/Sge32nfyi5RUUksg/emW7t2P3NqVtk4A2GhD4Zc06edYmgtcZEq+bzMuKg7tH3KE8jMQeuEAJAoma4lG9qm1sL9E1dkxAAAjaEkPaBp2ArCetLi8n0pcOrvKIw9A/Cz51hXhGvLWR9S0tuhQhAg2u3ZlVmk83zC8/AqW2eh1hG9IZdI8QxtaAwCNFs0J8IbOGfrIcYhq09pjJortFm7Lle1WJyWcuWYjWXhuBTKFMOxlWcxxEIy7ufkdUuxFoLZvYvN3HZqOKjYYqyc9koPURMBRVSGWpu6Rp8Jf94Uma0CMQDptpDTQ8g6HWIKOzQHw7QUajSg+L2aWlGaItPcrBRtDfF9FsZtJzuHo6kFnmiej4fMLZV16d4dmu0dxZX93FQHAXR0hoG7ZFIMUSBx+cIsrTWLk7UVLE5iOq2pjdnjQ9AFtg5QBIjKQzTX0w45BouoKYXJLzItLZ4DsHvbFnfxoih7sqG4lEtaN9eMcTBUGgVdAxJ/rVMaPLAZWSPBJUl89gFs2rHf4WBUkV1rSmGl98SUtHkpXKMo8YbMTDQ3tU3pUoqDhRamBChYOGvEFGHUUEhHK+S1aCRAhVIIbuXQICoNRVp6KlZWIAajUehbhkvEBLZLMisNjtFHYiaDuNDsiWD2MIVd0IC5x9OSqfneeBFr4Pmr07V07zg19xw0C95K9zykoXlFOWKwqYUAbKSjV6Uw48D7q79TH9JtJt9sLkk/dwoxFvHO2DyPItkBqkueO2CKaqwClfSoVwMgLdOxQymhcCJccu6mciSYy7SsCLKEwfk2SNSdHyEIMcbw4h+6ZrDiFYGDaILwGkzhaSgNge5UWNr1EMuD0mrnaLjDpWEIhaFYmldjOmMTVORBrkQC52B9B2sXRBI0NdddMUpudGdb0uGMGEfXkLE/5ymK5nyNCC0AjJ4NifeQzuNy4RuocUyeU6j4vL6yni554CjgZyWANXs/V0aFVj5xgYMxc+icQZEFbvYuTO0VFUxoGWYIaeafLznLVLWblOVHT7detb+HXYioOa1cFcQM1iKIFQw2rk1wOLc4awAxK4SKkbMheY6r6g2KVbB4CjS9Aonp8gzX2LRFr3IospMO1Ja0HppoerEAACAASURBVF3pi6aAiyA8s5VXRDIrSAFTmMQsTb1UnV+Kph5Oe8aP9RPEEmKeiLAoLL3o1jRG7Q2dJ1H8XQ5WJbCU4pO7KDvEJTjVzGSVCjDrpQQZXi8tK03HmqFZldxOT7qKy8zgvL1jfRiDbVrQIi2rMO9tykAXRaxGU7hXYrciMEdmVz+UodomdLqAjHGbSigaChljq0nFMxOaxHTBKhCPTzWet+lftdx0TQvcq0Baej5fkQSX4IfML0E2sHE4DVuwyeOCrGgEkiGsyUpT0dCiOwGnlt8nwGcxZxZfUalQoS/uOrAxSv135qZezp4hS/yc1sLPmPUN7BtYFleB4pW2HlYxu8V3WZwGtMi0gNMCCJlPnQ7NQp8otXZFN3Y0F8FOatVS7QzTLMxg4ZV250zhoEIjzVeuOKjUi7sRvYfE4TIiGV4BeVb8Gb23aUkj02N6dm5AcRPNcHRZmAZmF7CPWnDBnZp2GE0O4+U58/40MpQFBYAFXlPjHkmz51wNWcCVe0rzQYW0RrasL3PyeHUaWDu/+swX64QdrPjGcq69wCwhwAZQTh5i9AqFQJ3SugBxUCKIQiPWy1N7w3+/702YGjrC0xU+bWLzkkJJy0f9SOE2TW1FWARK6S1QW9J6mUDaoTDrkSyTXYS8F9+DuEOVzDKoSgCJVBI7k4/I0HDCkulAK5j9Lwyt6Cq21m22RrY2F/cRuei2wWJ0K2lOF76v/uyvAX83DYbjFHTxVvG0+lISCCYdI0bWLiR1j4gdo7UY3gEQdExFrK0LeSS9oqwa9pURTq8c/OOCCfIShUPj/hxxQKqzfD9pnrhBPwKSuAa/6FmRByvy56qsOVGneSoz1Sy1bppKv4rGmbNexMI68fkaCZwqaV5SJsOZ8bA9MK9q2AaVNz/XG85aFFAfORGGxcu8NRVVFSQe5MxfCjAwTMhhNIg/KWSLCwcVQhWLj0j4JvaEtJQqXhgiWVpLxVAprMj+ktb9/XTrt3FBKZr5adZUpMZECIOouZt8D05zas4kTDMKEvQs/ly89lhYVttpbhjjsZKO1l4EMRVLRGLytog17tBi9QBSLxgAHH9wQFjTStNtNyucnxexcYeGnVAROJYxJDPTa4gQxmmwdnO7dM8mSI8mRtmT5oqYnzA1NtmZEEfBDlLQqqfUZ02+WFxJZViV5eIWlmXownmXAF1kCW9Ner6RXW+OqUcr3+ZZewl4pYdsmAjXRTA8YUqfPMjnEiDA1V6JpHfWF48Z5rJDc0Wkd0MJIisyx5LyhbILRg7VDJM7euYp+vWYftkuLQDkMISaipCe2mqQMJBA0m0oZoxYTxHK0/mwDqFAbCMZm5Gcnok/wDR0eOKSmoohgrh2YLw7Q2MgicCqQgFj7r5XIzoVnYDUokUyrqSblhOg8nfs58novUew7lDv4TRsYxAekmDTmgtDWlkRFlYRcOQ7pkvau6CqCNSb691WNd12TuZyhR9hR3WFNBbBxgHAUiSyCbNqxPp0MyGIknDWT6SnlmlXCmc0REkW5rBAbBvClZ3FMbehScTEfE96NixK4pmPhRkriRUKjJ0t7rfPcFAOBa4fkhzYjGZNCekkkBAwzioRf3eApewSIVERowetZIEpbYV9P0b0ddkTkQyx+t2/lMmp9V4cvALZI34XOmZ0mN3hwBvKDOuCWHeymdnDAYwwfmEYIbCz4vg70j9kDiaoTXMvTHWFuvJO6gpvOddOic4tlATxuegMJl93grSofY7nPQCQsXRFScWYni6SIoWUxAir6odOJty6JAvygEkMFtWwi6/A0m5N4QrFfpHeC2d6siiHikyoDJApIN6D3lDTHmDM0KVfmEOsg64YP2Mb3BVbzQ7L7YJo+2aZsDiBaY1Ns9tqx77+np4Ln5FeAQRA0ejJsPdTNFDR7SoCEW4sM7e/ym4dAZV7KGBa8OTnqFdZXLH3TU7VmZkdq7yuOqM3WjhkqlcgMemcnk2lOy35XAxpi1CoTKHEoZvGxtYtPhUF34VWtenuOwgY5tj5NyWg7ooD0m0Et3CbXh09BZEcKrMsKTBbL4Tqe2X4NXrDlj82OGSnBM0R/TJFLAyjUCuY7vSLKboRBx3NG2lu1xkUO4VdxJJY9WmG0SEB1cBFeB/WTXCAkLhnRVxMXeHEsCtXig2IyVnDrKrNY072RbDggw1TVBjCF+rUD5XH0n2GqHkom9AFPqTDrQ3LmPlwigSzaLWpPISCr11uXDIsmt2CUmD4p2EY9rvM1xMYa0E4Wg2xAi8HbClgZLAqrvCQVYwx7sy5nqlHemc8C4YDTYFJMmVGnqGCFb+XteoTZNwlnp1thgtknCmwF/4+lVlmLaIcXRlyOWCthilU6bJDksJa1Pop+G9776yq7betkab919Ssh2GeeyFDWFSubSRpqUeKn+HcnRc9pblZ9yUxANVUGvDn3C609EZwVTdkJa935IdCT8ywCVeigTvYE/XX53Oy2I21J/RI4D+zIblZUMafAa4gJUNk0VT0nJ6lToxI5wb+4ddvJvyG3Vj3aWPaD6bonVxYWj+LxISDTXKqDI+1U1z2wEMRDGwYsoGl1No5MIXpL3Gi9fGYCSKZw7sm1ZiCX30WhXX3AkDQTcHqmMPO03CFBe56xdVcOwfDazw7kMVkRRDpxFm9iMvfrR/+MQCYkM8QrfMds6fScS8AifF0xgbC4aiya81Zjk3icIGReDpWuvvRcipoOY2ZBEArOYaPoBgHv+bnc9gtwUkjl+y0qBsmo271NZiadSlU0DziuVNi/ZRv9edtmr0fQFeVKTkOX7qfUVm07rxE2b2aFp836Z+Ff2fakhkGDoSe1RTxasi2ASoaw8IEbcmuTNKAtOaXeXD57nTz+8/wEel5EzQea4LbrIGwRkKvIaFR9bOkjNGTakuG+NHk1rIfhnMnqLRGjy2JxRCUjE5YP69cgWjfW9QXIbvMxbtpdsVa2GVdysNsQHcIVzywwmdApnfArEBJvgCzHH0jl8Jipkkz7YemsRuVh8sMi4IWU+JwKBi0lFH56OBlrdKV/OZSHr4Dsw+rIjsMwc+w889xH2x5wMj+B6ZJIey5kM5b6CZT9+4B4JWOVLrpJhuBAHXUiQqXTG0VfX0Hql+PIQWtQstUJ0vI6TmVztWmUusH2Wybhusc3g5SmMNVdXeQcy365jN7RwJzxqgK80K3LRv+FClszgKRHmya4RwzatWlj7E5XACnZv00SXP1LMRuSDEUM1j9HEl/CwttF42GvSKILXmq2XE5NzXkFIilwFRiAs8gLIlT8Ysby2YFtO56IOkdKNinE6Fz6UBiSc+qeobCpl4VtEXDQ7TCrZRTuGwwE8TKTBKVJeNstgNxCpf1sQu3qJD5bL0XNVSBCiS8CWXMYL8aDUopBFmMZUS2n4oLzehvTEwByOpCgmOLu72BauuugNP6LJqoP8HG0d0tEjo8oO46FB44w7JCbXY1niFVfiaAUKQ3sNd5BUMVHC0Nq1JQoDkR3ok+dNfiM6ycOtY6bIh1D6ABif8YRpThWR9PhjIUE+SpJbaCzhqbB2fvxrQvBwgxzKTLK4JoSgMEWlKhcpu7CYFEVS3pTmZavIGMvT/0JtQZkEV2pDHLtQVwQSBAnROc+mHEPBuubQia16Q5611oBRP/cUWzWAl8AbzRMD1J27PKNQMmZOuBRVg2G+RoVqxGC8NoLFGyhJ9Ft5wncTDYxZdmhogepSUKpBNweKOaKULiPcXPgIahqSuhZuAnlYlhGhayD16dxroYVu9ayFFCHvppZjxHApz9mZZi1af01qp4b9BmUbFsCHDUNA+RREZ248GJsmlWIcmY2ZjeHryepgQUhn8orO9DkTMUOD9RJMEbBVCbBHpPzIHxbBDMv2hZN/Q43NIUTSVn4JwJBU1eTAtyAVqcc+0+GhgCFQAB26MotSYwau/dnNCMhRc19Jmp1FGy+9D6JByIErExgf7uc0vvanGpLNjtH6DSriU7BhNcYydquuhVEDM+Zh/mMjjzUBHQKlPoSfPFFcDGy40ZVsKFnb0G/UwKBWJsIsPcpHkqiX7qNiDd9xLUPd1FNg8BUQvAPgriBqzxMUwzGVdhZ8VdIfRuBR0QDzZseZGeX/No3o3z7Wc5CIlZqbkppimB6NE9obEmngAk/pbLfDo8Dpl9sIFUOcphmrMWgspGPfwYqj075aMWYJ5NoXBREUcSkma1WLsCZZVeYHOv7WiyfhoONB5KgbKIiWDm0oBZvG+uI1o04ngMTAoOApTqzOaupH2/A9yU+0w9V043VhGKg3lvClvxgx0lKzDplhYhzmJ2gvMn6Ov0w3uNbzTcvVqAop17KTmGrKliylcL4WShFMBZi5lFQKe14Qw0illnliBPvbD7vfrS5wGsBNUo2IGk0IgrIt0Jh7ruRA8vRO2sWic8KAhrwy5Zu657js7oMzpcoPcKkbEr4gy7jtPunPlOvAfT3/QYzY/NUISFW6aYkkZj8Tmb7qazjHvVCQtDJnUJ6SsfeXZRN+Q8xloHKibbnZGLp/nVe6cAFRM86yChIGgQqXCbv2dbNAqbFAk079C8ZNqafMkwhQpDJJUWC8I4jY7KRtUWAi3gxDeTCZZD1I7mBR5CuZLiiEaTc5dbZt3AdQPG+APBkOYaXDpVzIIs4gxumyEenjQXpq17CCNTLCVTjRYX5/wKFSv1FmS6jtO6Myxm3iQt3P5QDCxzoRhLFmyxj4IVbMRBIGkp2cKuTlmz2kYkan0Sn3sqk3H6/pZMB5oFcqZBi1oTSyPaGLro0ZAUcjJjP8yVmYFBci+qZSYQfTbRWQsWHkksjiZSnkii0xUZojS3WqG4FJihEUrxuTgGIlx79WcLcExjHF2MmiuWpsyp4h52+IXXNc+u1OK7THuaI6woddL+KD6XNY0VN5+NlQpbQyCotJjdCb5WM1wcPUiaQ1mNzNksCb4WDwObawOGDORnU56OcXnPymY2wJCl2SLpbQoslOlnmVLoGUo3daNdJa6f2brEIrIOCTtV0dzAB2HdUs5xDa9BJVNqQWfZ8Ug4tAmwMCZ2v4pARmGXohMr6ZcpRCExTWtxB0YwGWitJFI60ml3LkYWJCCZbr4Bew0arn11zcTD4I5KxvpUPuLMHVOW/R4EdOgZrbzilJazSP6+ABB/nt7i9ZgLh7+07h1YySigB8J3T6UrLiCUTjJiv7czvBJJAJBKxVxTJJLtocu6mqfDgq+CBFH7iVMcCc/zoVdGD0NDQEiL02meCvv04b6FguNMFqFAs/j89AnhTO9qy3b0ppk5yPkovB9iSAvQYSzu5Ww75SktlQa9Kg7d4TkWkSgWJMA8txxGlMrLlPDUKRzD4cCNgEnzkinMUNQugPwMf0GRCqbH/5aF1t/fzYliQ3glQierzk3sJkIpyqH/m7Us9Eo5X5cKlgqR5lCR0EENxstQaFEQG/Hx4i0FgKPSCdpNatZFRMMi2aGyZoIvmQN7j5riwNDTCEPCykvGfFQ2ZGIyHst3dwSm2ai/cKP9ZUUyg2GeDtNMJsxrt0hctmPLZRCAJte40Q3jc9DCnVoce2iZr56auZHMjvA5Nh5nMm7lNOUiGt5IccLyHhpxqinOfhzh3BxzCUvQYR4uYPR0eMbaMj3cYxf0jDg9fe5oMLg3RavFYrK+KI7nTfyhVwKL2rsfDFyalJ7Y3CmiKLcXi7FJE7rPBEjVlcO2AXsleYg4hCCVGsRSzEBiCnujRGxOga8dL9rAoMSYWADIIbiHHU5BoWIoQh4PmnuLPUM2eiHkUyoPQH3PiPnwqVA0lKIAUUdRhELr6VDJPiNmfBY/kogQpatVouKBRGepDVDS+N6i9FTUMY88s4QgfBWB0wXrItiSsSDYL5b6bLABvU2t0nKUBCoh9jluJu83qB/4vHvpmKy6Nm9AzAYUmELpwT/xuDzG7oFhTmIazFz1TExGX5XeQ2Ipc4YPNiWabr+9x+Fi72YEz2xNMQkO4HBwBjnD4+Vw//2L4/gZFxujeKpSFarcHG/X3rZm6wCRnsro+E+UGWsqQ1PK2WjHCeNDyRF5jI3pdVCwF2RczWedXGEUsD/CznRvyFZ3ex57mcHfhZPO2bMisCFEFKCgudcXuOPUbRJ3mgPxs+LvsZkb1JXbypnc8KtUXE5as4iunHuLyfMnVrAq6dqTT45ma02wmgxPTRfZUdpDkTCaq7VERy89XwodQJryvd0zJQ04dV3ghVgJ9CqyVJ84h/g1aACbn09kOQSoHNfveAsHBzVFtLlLs1UDlOvVYPgGPVoLHU0J7Y3GG9wJW9xlqQU4vue8T+vDuNosQBdDN404luPy4YSfmsZgFxZR7Q8lrIR1I1Jbsa06CbqoRoclmUmd4bhkWSTdP36RKIzvieSTwOLX3DoDFGRTGVH5pbsma/23Td1VTdeb2622xEhqEo3jy6ZmVlU7l3NpFn6xOIn34n0pqBaiSVeRSUHInhsKBydIs3aDrn4M9AnLl/0ZDTYpas99zc3ig4hbplG1e65+AK8A4YpCcmjLdkn6qjq+4DE1p6K5ftwBDunSsj9oh+aknytz6TJaihQsxuNUYFlzYQplchqOpcRYuyEsscYy4JVjA9vZ79lhAxyyYxiJT+qCeSPzoiiDZScOVl3BmyLmbxRgl+buuXPORKzULJwSZ8/JJEKE7a4MuEaR3iqfk7Iw1IQB1q44N7MtqlK1UKc1jalfRRPPAdIboqc5LRpAKzMtDAHDZaXrs7jry85SpsyoUPphu6zbJ1Fp0RYnGvGGVUlXcBckhNcApIXtFHeAc2s/WN5JkfGfWSuNmDliaGeujbvoo2Sffu3e2XLt9CL8e/6ZokTVJboXt+79rCrArsKppdIy5udMBsXewPF9DKM0hJ1WxZjSgFx6KHMnaXRBIcRuJNPJrkjCbfX3iiyJSFRjFiHe1E+ESm+AQ1/ovdCyD4X1LeK1EBo0ZxzN+DsUYc3RBFwxiQa0ENZMIUMyLFWlF7jLl/YzjcxZ34ciSB5QcOiMtzE0jSlUDBHmRaNng4AxMaEmLIZTVI9VWPVKIJ18A1eKUAurOHCH9SKRqm3iHjSiZkLVl2I1wTgkjajAGT6Z4shD6LfoNRiPqhuuaDrzcyTgShxvXojn6U4mSQQxSIf04iBgEciggLIIab9KzOKktabQDCI4CoAu89mZs7eH3nMrQWXCHDoFU7CLVosIDhxFn5TLZBBhAq3ArJZmDW3KeoamUGINSMXXI/68rhTLIY+F4UfiEyUUnlsit6BcJBy7WTWR/gwNmNKyZ2rIWJHkZcs7cZ5aLMND5UqhHVw5HM2aOx1cWOnhUJgmzREArSVepH4N9t60TtEw1crP7tfiBUE9yOcDUDwkYDZsbqlg7N1NYey5UES2onWgpyvpoolbFQEOxuKKrJkHRpp36Pq8dEg+hUXoAZkbFFO/JKeNm8XM+qANvEbEPZZSM/XNZ6qFyhC+2Qtd01Z6ikPtwkvkAml6384OO0IKFSzuiR24qz8tWSEK9+Y3U0NMYveb5N+zJsM8MvcSqjimIIAo5sl5UA0brC1T9WN1GV3lBHRTZvbA5rUIljnpRA9rXqDD0aJBUKYipXtpgUSdA2M3IBmrz8SkO6k4dEYlUaiA+nJmKzO25iteb/R4mPsr0kMhwmuMyvoK2rZB+g5XWhmEVzRUiSVHAQphdwqUuft0n1mK7uGZCx3dQr6rwvATutSM+RU5Pp7vwTixudATDafwUgHw95gtGmR312nMofBzVE2QkVZOkNeM9Q1qYPV2MQFX/3uDxsIkCVpm0ZM7VTvAa8TANcPGw7mF4Ibl1xSuYCx/B2Z+xmrMux52G/TGmlWvK98ByhAPyNRzgJ/IuhlxrGE7+1SxltPQmO7lHlwaiKSPK6GCuP685C5dVXod6bITK+HyZj4j339xHsk5KZztmaP8+0Y8XpfeQXMhk1ByiK7YlBTEIqKK9DBU/Xy90nM7n3ZNmCIuPc1dBuZmyrMWyLBPxNcFAoLOCzht0Ksz6KSG5nLSdoQgHpMVSdepIRULAc5t872eHT7S8xPjOAXdX/ccJP/OYSlALryhwhslU3BNk2Dr2oU6kOjApKLj/QsyFmdBDL2FuXt2CpbCc+Lo0fw+ZEqr25fb8two9AQ9GQbFWkAkKKeae2SzB0OjcYznRFCWhF/XPpzoWpWRoRGxkoVaEImIR5jh4RqrKnkmFlpS2A3nGTsLTi+N6WyGQUnzxMn47up0RrV7x/YwQXgv0FwNWBwwz/BIHKizu9A7Yp3E4BOPmHrkGsKY4KUdzd37UResUNpuudUBy9Y0wpSxmnc3L1nh2tyC9XNKS0lvghXIAgcpnUc5Qb4PS8NzIc3FV15WO4f1mPw5rDpFBMTKx0b+VY0qX84JndxVmmZ7RvOypYu9/HIEyRSJUVia1V4Imk1agCmAw046qAQauJ0sATTWEdCdpzViCfIgrJrsQK3k33CroUYMpnopDEXys72GnxpiKEk0BoF1EQiGZBUlK/b4ztZ3Ib44ONN0h7MX/EBCOZmgaSDNMcdD6CJnsRbne9ByxeZqyWfh8iOew7RQJbkgoPOGqAH93Zqf07KjILryXgqPCzIBOLrmjF+BbDpS2FluONVKEO/JazA1S2tOhcT8f7y75M9Jd2rGpF92+XLSNbEVPl9fK0IBmBaNtYf0NG3eJcJqs6CLo+VK92z0rIaaRqGp4mhq4cn1TWNN6WmwrF66LAYQHbKe5WH3LEF5Cj+9ddIfmvUVNAo7z4/8mhd7l82cG91Ami9ZUAYPozj1rBYL1Yaa6W+juYdM1pik4AIZFj0FSOmHCKTFECBKw8kAqyLYq1nkREGHIkb/A65pG0u78rqMlflFgRQgaitIjB4j4TYxMtq6lmBOeiZksl6JMIsydRYQSGCNG+UpsH33ZLiDLpEHg+wQu7pCECrXYlqaxG55GX/HfG9aZ54pU36WIs3wig1gBMCGIiFw0l2L70vlQ6XNArRKK66stUmB570IFNOA0ONZV4mJ2/QOyMgsMlJoeFTxHMgCLlppSIZNArhHIEGT6kLWkJO3+fwcN5fFZFnNGcrT7zk7PmTAK7VS8kPfrcpJW/0Xz3FvLEEPkbwnsxylWLYkcKNQ4Gndg9cJgKop41XNhrK+niVStB7CDNX5Li6mkSmJ8KLkAOBpMYxjcA8P8H4ZTTkXvz4H9LD0u1ivISL7QCSZQ2uKiC0TFgq0hOtLEIeWQ5F9ABQ0xn5klObCySo02kXWEtgQX7dajdYakbKkZaBwBUoMVoka48auVGfwdc2dp0yLUtFR4Mi0VJDrWrwOIXEGehsAgbt8VjIkS9shGU9yk3vT9GwoBMUt06IaSoorDOi5EGhjapLe4OmWmeg1MQMKUnHFRs+LfFvQxdSaIOiaLq/ueiA8t5xhYnQkJmBMqeGp0ppzdSGnY8XZKzxLkYAgaT5FetetaRRv2X2ZrbFdou6VSQrfesgKUv5JniYvhhX351gPJqgUFDY6xogA8jq9B55Hp2Q4Rj/PI0f5qWvFXgm3ZkK8mfP3Fs2sFeeHWsHW7viBWuxnvfdXCxV4KnGBRDhJpcQCtOYexcotOr21fpctPdqB4FY/ZDWtrxMciFb1tfuIfHBmNkiI5j8lXgAAB0OJgS2DqzwWNCXbSbjHAMOSrmZdrF+kuRYocezq8yJlpwaEA3jpIk6aTWwb1ejBMEFDJ9gaByma11g72FZ575J7MNm5Sg+NTLTnVmKzeOUp0nI3zkxQDbCUgsy1CnTXV6etTaiSgswYlz0oUK+ToGfYMoXJzlFab7qZ/XSrRTODw7Zxru8Tsf0tDB8Bz6640uRSbIFlO9gbkoOWtUvlZhAVU6vEU9sdzeGIPTQzV0CCiEzL8zr0dDmdis83z9nzkzTP9xfxs0ICs0x90nPgZ+hxFpGYkRE0H4vhUw7YElDvwwFFYhikGelC5W3PmsqIPEpPtSmiK3UBKzpdHt17XA2Co8nSw7x/DIoizV1RaufZADnbUwCUARiKyGCzMHlA2VjDuRGsPJTuRbPNK8HJHiyhawtkByhBM3okjA+paCZVDGCWg4whkRKrRaPbtYotNFZXZrWz+ABDkxzuWpzJea+BDOwhSCzlVQcV0TOmHRmtGU+BDEqrxuIvqw3IGhRWOgLEWtIqEkSlkmMpMGtR6CIW0eidAYCNmrXcLFxe1Ck0eCmzu9qsr2gt4+8qiGKs8P40p6NRkKg06An0cXkRTkZzQRV3gVvWhxBboltPK8Yxb1Mzd5quOj0mkZx7Sq+neRqZPEg8QF3gOJ1qUbblC6Qm1hHbzCFRwMR36cMrw14kBIkkJ+ZgNPdakoXKN4fwCrK+QwHfqZrKJXevZJ9NQ3qI05KYkYseIILt3CyjN7Nt3Hhtb0gPJRYfFTOWrHMS0Osw6efYykW77IkfNGlFelBRL021KCDUaIJc2AtkaS5rx6lpyAQxXVuoPen2pLXpmYyfK2I7GwniCAyXUGhsMGPqjXHbuqSmY9qOGRHODiWTsr6DAt90l/BAejX8k+9a/P0F5qqxBsViUgs8uEmL2EXsE1EydzI/8Zi0aJJb1CGepcjYlLNE6BnsuTsd2Qdkum8kg3XvkgwtoYgaD87/oPdImjN0U2WYlr0tggxXeA96f1zyZO+anZNUQixWs2pLRLoWbgTWg9O85CwL4iqM3ck3PFtiYRzPT1pul1RiJgjpIdNXoqVe3KqNNfmX9y5OAxZ7qSZYq27tRAgwm+oin6ab76nYRuBaompYgEgRM3xgWwE9nb1RdkKn1rJ4bKiZ4lR4da0TihPZOTBJSHB6TW40xI1FAOoedo4++CflDAHSlyJSeoxiq2YNLEVKpvZ0n0gwvnpcHtbChZaMrugawyQLt+i+EX9gZZ+AeAPrNBK0ERfejVuqsSQTU7moMzSQ+Autc7/1O0BXpMKjouxrHizzwSpEX64UmeP2EAAAIABJREFUrmoCZhQk81SSKAwVbHFSvkvniYbGB6xln1+xlBhZOMVdHRxQY55QAoB0LXlePFMRlpu7AVCmJn0OBBBDdzhhqa9BYIqVwtqHNsxYDc50jOPpvbDjlfUhPeZjfCGxro8KRkDAFzE9qml2UdJQedtRAKiCXfyG2SW+j7jUGG0S0LM6hhxr0Feexp4VJE2pdliMlQN/7OxryfH9tNC90oouXEk3v+dZKmtmccT5SgSxRd1oLh3/pJKjoqQXVT1Wo+LjszGTtjgeFzT3tOuypJKfWyqggTFS02zVBRKkpEBTUZD4JBB/Rsuj6GoNNBmVsR+zKKzfV2f2jV+AGpcTwNelYAGHuShmTZS9B6t614nhRmZbnNlDKPwhChWj/d7GawGmppiF6HqGEQESoa9FQQwCqgWx8ZzeChmeyD09HlpKhiYULiqifQepjpYWwlcjDOtCBH8mDkbhkB9aUAo6gFD66tdgn0lvcS3LkDzArlnekMp3UZ67zfSIEQfO8FoSJIuCs8Y1i/aM3EpOr4J9IadP1IoSdfIcWMPSddc22PRxf85FrSGxtXS3+RUT0iDR1zQ5CE2B7mtkSPPwFOGdq/7cZqk0wpGtW3uO7WNanSP6aSyJEfBW+6MZ3aM5MRR6lRkWZ/9GQSrhJokf0uhxJysLBktJ/s/QW3E0seOVk8SYyLDvFfFsCAWX2pbIPkGmqSG0C1H9WROH4ExICiwVAtOb25aCrKC1tbBj6qx0z8RUGIJ06ceSnY/8TB93NqR3wO9RaYA/CwtvmAdjxwbgyE+5H6y7WdKDsqYxjWq9zZIZDMb7YeH8+fp70kNbRXhg96NXwGY3IL0fVqsO/u6nW1/A3pvNTvQqZmW1pVuR/r2cSbbuNTEDZddKy0PQc+rSjUTpWbvA0fYU9qB5l/Hh9US8y3Vh2jxxpqhlKLuFRwyz+s80VxKqZhkn7qCAv0/LLEU/SZudmU3pHaoJ5Wl8ZLUJ6UlNi4U4qo5FtDSkuzS3vzM84XVzpqiGAJpDQkwpBZl8t5MG7wwDJL1hLlsmze1Z7Zy2S3rwQIbo7DbleykyRJ8Xz0qBf/dxfKq+vR62rCmAHZgQs5tU/AFpEY3IEtqdA1lTw9lF2LRFy8BDKEj3bFJ1nCLvQWkhM7HTdeC9SqazNAC2bqWAZMUjrzOIbUljxgIR6riXIznujAi7K+WI6azPRMJ7gGTotFnS4wqrhgQxeQbiLEQruV+ZLUB0by68vivh9ZDpV3WrJv6enPRcCy1qzl4gNmLpM+/cLeIT2vsdoARGc7dpML97BgS3zcXthuxKKuQKTw8KAVzEtXsFN/kmdOI91mWJHcUSVlPEB+yyuMs+RM+RaXMbk5cXUDjdWhY+AbmCohZBUY39sv30L8XuLFFKKflA4G0D8y7NGcoSC2juVXAd6+Q9LuOYIK+Fk/x34kFG83wZ4hwiGU70+E5zhhXJ4TYMqbh1jPfkRvWmRgd6cxzay0pSGn1xPiEQWzwtHE1YQFpzChAPiulQVtmxrZuVl+pxBItZGLoArINILRnaEpwYpeHakinMVc9eEoKRRMkVuzlnHhQPtHTvIpKhD98xFctuqpfvx4PtpyYPgQEY0zOeNrdeY4ZGf2asAbERgmzU03gOVnmSDjyfAKnAMyXwlasHq8DXHCYWwNeiEuzPlC46z2Sn7gCI1X/a/Zw4QcbpbKDi03U0b+ktVTc80tGQVs6YOGPiXZojXO/oj6m7ypexdnHshgVwPVAoQHSaCtKj8LA/3HGRrFOh8FeRyCBR8Q7OdNwna0B0Ghi7J4cIS1yTckA6WF/MLvBv4WRiMzwjEcT0KoYw7FROmqcsLc1xh6Y71+6VDjGcgAb8OaEa8sT71AKsBhpeV+xkUBKClW/9wxf4vEv/zuTamULOMnCmRIGsB6DgFSdU0wwbVPLvC1hfoUEBBV3knOpVCsITgDMCFUhTxts54zAyGkivgJ8NyyFsyNIdxmaszpH0zIaInwnnZzK1Gh4Admd3AlZHwDV9JmSM5e33pzkVBGczhCA5o7FYjLUiPFf+HHCX0b/f98DQZaZnkjRH5O/75y2CnaVRnFURW8j9Rzw3RbZyc0wjP7NoKkAFsPXn24ZCJj0lsBx1Idku6YUFTyh2vBgqbUBitH/JR496A9X0IFi3QM+XSozgIlOL3PBGutbSe04Sz0paRGm9K+yYywlgxm7DFtdd8t1zhmfeezXabA6mtekhKrJehKXjBZm0EKSij6yJX7u6q68tsY9Qdj7bFMqpcGKLkTOTYIxV4Sgxuviv5fLk2rmjTBtSIUxOsAUaOyuhiAnS7G5Dp4RMEDO3TwZVJIg4dBpPJXdJkAlFEmcZi1jxkBNq0RSQKoLGKUUl3z0tRCotCynsAIGsB+BrsQjLeg00hIbKJS18ptN6CyswwadSAyxc6AWHgCLvmdPAkEpLUulVKglY16Sdv0YIGHURVEnSjcnTBC3V34n1MwMkwDFOL6PCI3DJrWaUT/INGZbMy/cyQ8MemRw+HCGrh44MIZjOtTPNTAYkG61UU3lHy7kAizB9LSGYbOrSJUvqg5/cGrSZIpyY21CyulIljQ0nh0MS9ygFkNaNfZCsOm20/hXBpwx7pHtOdlQzLCVAvDigGq3mHZ9wKZb4WZFPSBtmRiASGSJ+v9L4Fw1lPy2KgcqAwInA0pTGJHa4vVXmYaZllS5PbDMxuNeSlprFR1ycw01fAuIhubE8axTs38yehFbvLIn4VYp0Gj6eEjHMhmXso+S7ugxFEY/4NWkR+HwsTGPowFmRdEv3qm2KX5cEklhiHbMJgCiC4ti04i7W1qsMGRatK6IoqAg4jHqHYe0cxN3GtEr0+GKordr9VkOfwkyB05ZNYJtZd8bk0zvi/SKWdWXKQr65WWFQAH5Ocy7/OX35rlk0V66+PHVpAHwsflg8pwdEYlcuvVwIYmFPvntiCopM/8Xofb4zFAtnf8LuvUB3+IsDchlWhXIXC6VXg1n/9cBCP40eGT5nEfX5ohI0Z6EiZ3nSK1yXlCfxrFKny8OrZvhQC4LfSaNVtYdfVGMsHj2OpSlK5d/togrgaNIdJU6PKmmO8OxEgKG3BDx4tl/TppJw0XNBKy7pujHnTu08K2LAZ4EEQSIN51/0CgDOzLB/UCB5GNz85OdtnayqKLAXbA1YVY1wJsaUOXA3uOBVmGJhSnhqSZW+vJwYiskkU0vpGYTbrxqpYfWzKAg5MMI4I/Qj4pdO2dE1XhVxz663kO42u+UpMHCYJNZO2c1emkcPwBgNkR6klRprur5UsIO3NbOYjlEg4/ucZG5EX9SHCJV0uWflHNYEewHdyUooMn6GZKUmkGlJ8ffnefKrada70Igxw0LFVSQ7Upkiz74SV9i8eCiTzAAG2KmCUg0k5CPwLJr2wCjid3tj5g5GbESTTgFD2A6PCJdqYR2KRJaJowALsvYFyJS4CLDMdq+NAqVqnN1mZiRgxoMpXdKhAZGNoQExQ2openUZCSxNgKF3T0xz7i5jUQANYgNyJWNApk+BDplGMti6ZBqMv0Mh5WGy0Ct2PpQsO+/3UVD4eH24sgpl0rluFIq15LwKAqsQpqY6z6h7JkBiGLE6UThgZV0FW69L2HTWJms+EAOAWbadE7Lt8zEoJt6dmI+db3MGM6HiOrsE0aR7TtKLKw/tUO0D1S05z3Vds8x49A3bVBSArVmkh0W3nu8GpOtuqXPEPQjK0cNhd/Dk3hLvsdO8V+DAofNXRYRxFPJBPITSXcynx7xUkzcYDq19QI6C2SCnefNBM5p8Tu9LAJRSIqPCYrSm5kFw3YCNlusUIdJg8F5Wdu2hNhB7Xcj7A/JZFgVQNEqvKcA2HzNDkmhH72R01uQlhuJWe+KzNFr2gyz+WWZSmNVbj4jt65Rz5WrP7r/Y/g57fukXv0YFWxMf5mKPwtZ0YhKqyQCMcwXEJgCR/LdtZLZrcHcpYBWj3DClbrX7HY87vhgyRg/XKA7LK+/8o6sip2U+ECHPIObpbDXXAZAJGS4xNUdNu6jXYSBdYTbtKPLz4bb54U7q+1GWHPOuMEtRSsbUvDfz632XLp+Nmr/PME2uzAiWeaLCLVXiIMQN1l1FJd/bvKvsQYnFQJJMYuW+yC/15UoAGPhxRBw9lcMZUdBlGSM7uGVhi7mdBRQRe0cI2Fm/ftpTn9UwRlbrm+49SNf8Rks/Z1rQlpWwPNepqQtx4irNeeDI08GcKMV+D2i2ITBDV1wm5gaMg3m41RUvDUQt1lbODeUz07dld2paa0Cp6eXEwF7AB+dyGn4qE46/41KkxV1/m+ad/TLETagEKthcJ6GE6U0ICWHPpYZZaC/09rVpmUMuYhvQD7jcVzs32U+Cqwk5C5LXKUCUg/PORHRZBBYaHkCTflKU4yPu6dAjABLM5GyF3lJo3CnR/yC0M5KQK5ENTwDHzMHqOJyZ0MVxfF9WLB7NWfUpyFBsrIJR89kUPC+CoYJlSUXAVCzHBZKZaNmpCNBy9gYrhllDwufj38dqYCRxFnUsih6Xws6WuEhsFfd4fWqK/UEwkzcU0eELzWnp+Y7qZy6oovEnBWXSrlXdX0dcyrJUXCLFWYQYRHZkihDwy2wCLb0g+ZLFb+TvPpwx5tcYVssCJ/VnJy2zdsV+yOrTI6+zYKUlS8O5aLiXAXqmSwNEFcucKVDKj3b34+jAohx0nJ4FIBAPNaoQ90ovUASoPqLQPB3FvEhgRM09xR5zZPObFuuynptif1Wiv4RhXBGRQQ34DutI4Q4N5HFo5M4lBYZ9AxWsyDR3nRgFkKEBBZRFPGToSubz72nL1YQrdzNRIvwNq8AuQVrawT0XpmGJ8DJtCv99ChpgDEmtYjiE+DKl/MzgqRsq0yL/X1lnk+VIDhvhAJlS9fhcPrZ9Hq/8nlfdpVKS8AL4AKpHm5mqLklMEgQCgb+G4lJY6+A27MjxiA94WEReulkvro8Vh2I8d+7tqSjPKXH4225dqKXcPxTkO/0YBJeeEGTYnsouwmufeSlnKjepynXm+R2BUsK1YO7Ic1pegHaPvqbp7e2rd9u9nrPix36y3utqvoxJ7lSF7tVcBYVQ5CtAqIau7UgDiMQ/Lr9KNh8jQpkVOVLnD7lApSlbaUCJSlTyk7VcPUYYvCrFV5/xVetQdj7zGhY0TAcyUxkXs0giI2EqzrwF9J3oZ+2orKZ3iBZI+8jhsUSjFgIw8u5aKpZrWITclUhmd1W0u+t6phX5jww90WjmzDNnc5daS7NehPA5opVOkYSONeqKyvMSsnnVeWuQExHt86/jj/vorNKXTbDEqRB0IKF82DE6YYp5JSP/aCtHGEj6ZaSsx+d1Fye+ta0NF+vMHCULEUHeUtWyBKqiCjAbtuR6T1RRxKL4fGn6CW/p26HPTD6jvXx8jyygJyGxqeh38Eyl0m6B9M+ldC2P2p7Wq7EXBwqBM9oefR+YkP6YrZADRv+7+xgKKs48vpdWdfR/OC8B+yAFEkF+3JsHwd9HuMnDOEPmfA7PRgv+MZrHCVfDI8tV/fzv3TKDUiMxiUgbWcVxLl5oYuhAv8ldrNWo4joMQazRimdC9Fe6864kha3zYhhnCYn5fCSqOXiex2h37ZlK4J8c6vq+/V8kcqH2vP/wmUokcv1enUhTeQDHYXkKE5tY8zy9Y/BmnUyVe1/CF1YwVkGhGmnStLKnDkNqboFFx6btFAYvRQTfEdbYk+Vu5LNSOrhsPE81c83vvEZMI2NKGFESLpZbhD4hqthAc6pbQzgff3ENPAtcDtmwsTavafPLd1nsyMprrqHyGazrIoDwNGY5E6FQbd/LKychLtKRoGQBnx+zrQzP1M/WOS9ccj5jDpPlv5EhWvxVChnP4OyP+syL1N0Bl2WJynBdvREMlts9DMN7RYhwDKsIC1EPrO6dStgxHNYcmaub+/68m2QNOW5CPspNukx8589E3s5xCtUgahN+7f28rBO+1gKfNkdHR3kut6k7eo/RSAhy9etSuROuLlOXIgz6fHS69jCUTWS30gTnfXe4NO4G7Re6UpwzuYZq0LmZ/JKCvPuamXrsyonTbV14PcyqAAslEhV4ncBB+A2CkFh7+ZUGzCVExHVq1wTkYPnAWCMgszxGKt6OwMfvH9auEfkZlgoNBfhOiP7aO8J0TlqxUthyfdauAUL/ytDTTnLuJ99jQzU4Wd6hQFADo+rMIupRijZJOE9lUntwIg4/DlbRE4ICPAiqE44/Ri469wnUw0yLWJfrdWdPiO1FrtLqPw4hThMliPVEmEmF5vR2CricJLjDzzYGKn0iFZl9nPnI/27HLWmX1WX655ERmd0NghgLgXDDa3D2prgEj8v0enfYFUXDOYUMcwbx3zmOlnhSXVyfzWdhHOnEvZWRuWNk4xygwc9O+DX57nT/7HO+inv0tyDU2u4nuSr53aMNOgEC8osgLV+Vf5EcyoAfPGp41AECcp9+Ijxr1z+ZAbPVLgGXBKGdOnwzD2Vg6hZr8zh0LuY5jEbWwk2jmnc+wJymR8hYv/KwILnMTF+Hb64SxIBp+NOmbAzjCJ0XhEJbQJL+yq5SQFUO1uwIBVuHd3FnXM3m7xQ8XK2AtOFuVLZoHXynBHdYrOtcYJ5BQangiwPhLMzCVYu96E2bI7IsadBKRTbPxUWaZrquQBe4N5TVnw1XmpRuziIQVpK2k3PuaNMwkrNi8S4V6truNVPlOUPBcpbyPk8uCZYUJcmLEDlKVOow4vnivKRGJ19Xl+6jlOrME7IPWblVKBDchihi9MpAZl+QFQoBtzcfw+WuNADrUCtKzeszrJQHiWmePyvXx7mioFg/4WqeXcdZ0SXrlUQuqCy61eV+7h7VIOvnHuomQdeftXU9x0f+w1STNlQAA/fIh6erNr01UQyEH5+ksMpLwQwL4vLkMPBnXQeBmE9ryrBaXnCE7jGCWY/5o3mh6oJ+ClddziOmTD/DgMefCOK0UHHRP5NyuETb2goEevGA/+mfotF5oYjHsc9AW2C2ScXXQOLFPnkhLD7xVHJXmqAg+LwsHBfjbOQic73WUTwk5aT7Ftb47gxFqpPTfl1H39EU0Ofs7MynRcu6k0swdZjvtF68ViLDKO22UvJXwowxm4O4M/PxlQjIFPI5ju8qvzuFiXOIEHN8Nsql+pqk0oYg/awzabIX2UNmcQujhX4jAXQ4PMM4nrtcbKnmdBB2RpmDsiCqMRK7ni2iHhgXulvBQUCYxgyfdDEW/TVUbwxeL9cgutD38CMz01f2UpXJr+cwe5hVN6btrtfeNcjmJDlhmOl1uIWf49VZ6uZgDsf9dq/LED6kl3DWRTxuN5aamg429yfh5+8c7SdRrWpSukE1PNa61P5rdh6JCvpFBIfEMngO19b2TOjKdbzds9OXZ1FO8B38+5U/Y/Hufc5S9brQ5IHQVQtfn9+f8J3kLDNmo2RTFe+wHDUdwHIsAenp2t08BUtnKbC8L/8s+nkOFJHLIO0USq3asjkDjeIzflY3KnrvT1lxtYKAeKv6iePcsa5YavIpbnd55uj8ee80LlYkKjkVJz/2TC6GVGxThxjNookyoy3X8kIG2+04q86wZNTk3H3mc1qdBxb6vZugXMnNRAJcuki51jKO8D7bi58wbyP5eofr9HPvzN2ItIUYWNSdzMiRmHnx3UNx+YFeQ+Fl2v1qRfd6749uXyP3HwO4VleD/7xlFwx+df1VCzZkkxQ+PMihBM0YaBxf9L1I/mgtJ9H81wq2wmvU/JC/1tDVlKGEgHBbRzz/L22NwG3P0KZ/XthATP0aahiKizBNWrKsmjT9eIeFac8G1A5iL1FPbv7XaN+WPZE6pOpquOpqn7KiByKacDzPPuoKLFNxj9+DzqofZm5+oTTv+g+s40lQe54zKEmycjmu0ZzFGcWgLuSyGLA01Iofw/pAOVq7KFuqKVcgmA7PZng0z//slP4gfTjXJW9yUorPRYkWkvJPV0SswVth7uSQaGN3TdOdt+ZrxqXTOqIPI1y/7sTtOafGy2UeFouc7IkdZ865DCtlFx3OusHvGYWYyQE9L5WiQabojbkSMcf7O5MUpcQz81+K7KR2NT5c3Gk1NX1endD3nPLL3d1sJCmZPRrQMEpSM7XL2l5RAZhqajDqYruXFeFFVQUKaKgzxqRgn4FLNrp+5LRsc0Tct8bo/QUJnY3wPpzlritb+FsdmDSr/LbXXkKtEKJhAavdo5kPXAYbPhKmVLjMWlHMkaX547MyFpg6TAU1cRd4hZLt35yNixGmZjRUBU2S5NuKh8DV22pm/M7PbWvfa3pkAdtyVVEc3bFOV42u0uwxLg7fw7HDQXA5UZSQv1RFeu75Oeog1mWV2fi61bkACctnfurZjZ305jlN+0B6nAnnw+VARs9qYEKrr+X6ZYy7UPXT8GON9BQJ17YNKMe3vCNDIJzh+giT55Vo42qqu8Fksb1NNvrs7hWRD0lZQZ2Dk/K9oJm9XXfeQAwLSiGUMKjC9SsjKTeoaGSgIl0wDWksp5eEVQMTNM+dgosmnokKeMAe/uOVMkySUghb/N2ftfVnedUWwHVYPtzIDeYwYihQX178TgSwHiYfHLhJ8tF2ZUPZI7Tln2ncwXEQkWhtTLjqvfu7uTw8t4nWcZ5Zian8cj13ruG9g8d4LU92uXNVpPaZEahppl/XqEtnx6WTnclNuZbck/fuRDQzFQoiMQgFxP5yNsq1lq+dgoNQUnvBGlzdRJfn256Qfzdhuj0I1O/3TuvndZG7SU27Di7p6xofEaFWrJacTfcoRTFI3VQZTmdiWSXRNhCkO/L5cFsa2eJKeK3veTUyYm9oF/hOeI5LBZm/PS7y9x0K7mf19/ECEfF8c6jmi4C6y46qOSdkApm/VzdNqsY8it+HAWpiXZw5hnZ3SkHsQ5/FSZqS0P9zR7brNYxqRy9fBuVIR2igdyAgL98UKKq0/LLY7OfwurDDQiv9MkJ7QaT8ztFus1dWioCuVL8SFbjaMuPfs5mgCy7xWbQ089nqgiQM3JKWMjKjDhO7mrBlWVwMSVWVaLMtPtPeEfoahzDi+ylXn2ZlhV8rUmtnWgvWDnE408elHyoC+2G1vcmvaguYXMjKfUFprLxMhIendfalqVPMZZClqvcB8cjcJCFK6mHLUg/J4TklKyVLV6ff945qyHyTySW3dE/izP959EClOvPcfxMoiGhI57BwVnTzwlozGQ9F+zzyU3iBcoZSoShC2qZAyXARkNtfzIo4LrSOM/5KuZ8WKOfeXjklVG6nrktyMz776+oJ5ygwvofExEeSjyC+UYxpjm8YoDAlx9GFdRTqsWbk70qGONbV+0JpvRTRr+t22t3HBjysp5xb3sq7ZUY/G/ckDvNH0oRAUxfWAJi/eExvtwLXGgQTOQ0B2U9eQ9LBO/C3kUJdboZ19WZchIb+JxF4+m5Kt4rpZjReJZORnIQhmHni3PT3iH+ntoBZpjy16zMD1T0EkAYy5BuYgvC71GnrKKlXXh7qJGJOhtUhRvOU4Eu+ZvMFQGKsTyOvTjrSCDKNdIyA+6pmMFZ72JDcRTl1N4aFEzjJbClcBJCD1OiNMoK4WPEGFELtlXr4ztoBBwhLcwFG7WNzAhiRsNxNwhbqE1mwVs88LBWoN9HpZhVtoNgtZMfrzLl89/IK+ePK8WL/LnXE6mz0MwVK6PoWFOmdl+Ux7ejj2VEKl/T1sCPyo+w3alpZZXe2AWDo1JVGHaNanIfa/ccwvTK0Tqbre0VkzL63dGUhSUAXVe1AGqs6UCAX4TSSl0KZdKk2sHqr+YC1pemHjw8cSyE5p5gNC9j3rC+OxUXVZlz0rxH9nuZEMLsrtUuyQ2i41Dvx1lCEluReyogLQfUjfImpSVrXZ6gOi8Ykd8/GG6Z2l2IeaBde3U6+QAvWMFU2K/szLXzV5WfaeluJQElHlyOnYtdLeSnX+DDTa+0S2u9bxWtw4aKIC2tyFK+l8K3ddSG5jbHW0eQkhX3c/9sjdG7WZ82/eZ5JAiUNi72q4UK5NpT8VqOZs0XiOaqAHhI0G6KuxJDpw9L+pBJ7zB4tAMwf6gHMnnLAXkJEX5mPcTZMWjsTwJhOtrp4DyXOsw/Tx2gAkIn52TAq5WiCHJqH8Xwe0PX3UYQ0EtWQsbp2RD/m7IzRSEvvfqCmzkkxg7NyiE8bw0y/Rh8g1mZaNjcxK+JTAvIi5KosRghK+nA+EwZP6yK0Uiw6YsDIo85JZM3AW21tEmTHe+Lixb+dfQOUmpqWahBSyH7IYoQKT4KsR73F/z9Gp2hHJIY96AjLqTBY03PGsz8H1ZHtaZ0XyVPLDmPIUrsbp7U1A6l0bUBk22aDn4pOWB2899urgvTkBCBFzzO/RrLh6dIUMtjqnAzh2zfhy1qfyTXxfi4rr3vrY66ppdx0tWmkoZthMgjzNjSPqtBUgOP0rw/rjPLaLVvU8XA2KGjK16cxBU2FHnHv4qy8eJm68InYoqmt1f7t/akY/n3mKn6gO9P33qA4Lwb21pk3h0FSXIXndxeMyYMOuBezb/LMH6Nd9Pw9bhuNmoMczca/1tW+79v9Gia/RrC0LIz/pZisGpqaaao79nQj3G6LftfP0shkge2d9DLyc8IfhOFPMuqwPMWOK/Ik3CMV+3vtYovLt02kg4EhxEdUAsiHZSPUR2akCfeoK1lDuDOObh1RaOtoZVnR9NyL93LtoQ8rVVxLnhaQj05M5K1QtBaWq5Xdn70LFvruaNLPaqRG4RPhONwwXD9cyZjxYRojhEqW/rHiXIg6cKY8u59nrm5LwGSr92p0uP2z4UwO6S4iGSEch9Jd2xPmc+Yha3Q62/k3svDtawyAffZAxd1I4Cg6nQ3r/q8P+6xfOTu5cUZmndUc7sLRyDnPa6QSf6+o2Yh8IiuFx7wXGYhHiZBVTY9lVp3hS1G79OfdBGY1kTKh8K4UAAAFJklEQVRp341s6Hh21nuwPvdwq1yBMqr/Rco8MrEV+RfXzDwMmeboCfbPy2Qmu4Aww6I4y/Iy3UJ7N+TE9+fgyGiTvDTY9956WCwMQqh6NKj7QwLlyEGQdeQC2EwvBmBaWADLB4zPRAkA7d2DTzFrviO6f3XRE5dLxyVDaMr/VucKuGccfhxIyDp0RuUn3M88LAbNUmfuh7vKNWOPIF9BFvF3nQimdIXiAqBE/40YSLyhH2Zc7jh8n6Aza8Vtn52kSVx7zo4EkHNCByf87+J6LIT6eSCS4K6U35fIxRLyOlaxFT7WGgVFTQwKFkTHL/D1V/rxrg4DVr/VCSKK5w8XRpJ38WEoTum9drkZyNAt1RgBeAnSsN0lG8eZDxPNh9zy2V2dHKc2NJyROwRiZ5P6hqeKs4ozPwj2lI17eVXsXkm2g8RjL9qFk+LcrlS+uBcoNJK6nlejreoZOoLbCuMhv9yl7+2l+csqW/qCo/sxIEA/3oJAhtewjs+GJWlyMRBLl3RPk16rrTSXxdXZjgh/dDLKrE/1YV20QrNWJGv391MCLgUL/zDT79u7bZ438nDP5x6ZgZrrvN315/b2aYvIMz0O5Xn2GbhSmZ2ZoURkUBSM6cMCUF0qU71fUg0wkntB52ktvISfUR6VZCUE1Av6b89paAqG//veBUVpslOdn1BSCPlUZSsS5qVMntEEUiuoc8RlhaoNwtWOfWhCkxqia1gpZhrn4kdfV6IR9QQ2OAKpiVyZ9OcnLtTrrVpf5PN4kZR0m7+TIJS77h3Zopw5TY1N3XODHIY688HnqVAayotz7+rYuEf0oTib+Li6cY1SeZLbFJ3kkjdCWA70mGJZk8WovakEsu3loknNiTyOVoQVWvU882zuk5mhdlWHKy6QIdQRHZhuVZuhRAFvb0ISNjufr2GTNwvN7zwhGvUA5Vsb4n0O+wnlQJdwLBEHUAVa6nUtl15rl9CanUSraiP4Ss/LgM+6/GDsPdJ6nzM7Fo1OQcbdxyJyYU2ZKq3+mQxIGpvI4S68ohDsk4T/qSIqz0YxZLpKoLbjfTuS20JIs+1dIhK5KhOWTRl/oSxPlEZbfxQ2yO9UsH9HMHCZqknu8fytyDsBzo9185lbcYlnIpTKOwBJ5mKx6pSLr7wEjxRc9qgqUPUZ5QHtAd27dib3dWa4O79DovlvG7a6D2ojhYsXSMhKrtg7lAgGEIUgV/Erz+PM2W+zJl+ZPsehRre5Vhg1SCiRWCto6d7ZoEhe/6Y8l2rLmHs+PVEsd8xM27df//v9/q+v+fzP7a6Xy64P1BUedVySFg4Tm+CV1EOEYE7pvdxCFqOGY0p6rW2uGJV4FO3YNeTE8109uDcKxTiUSPDOZB5P8skUB+PL3UJhmXcRUisLjDU+IXCbOpX3PlBbXn5PtOSSbXe/vQvZUn/526O6s9ubtSaC+HqvHYrKPmPskRORkQz/bIobUZFQb25xtbJBjrubvffWNaKSwJV7CI+UpNjeuziGn+0FiXFkEPL3drsGKizOHOhI5i4uWwjQtnvLx3ER0pXLM095MNNruZnib6+RCWm1Xsc4JkQmJNzZjS6zGeXTnhnEFq6Al/IxyVeiIsvnO5WZpyILOeikw/cK3WEZm/z7zJe7c3Hz88zkTpUu3ONdzlISjvOzzwSoYXnmJMkrWgihXjU+yQURkE2F5y5ZVpXmbZA9phxX70mbf2/X5OdOd8/QSSPla+tesmuyxLzmfyJ8ds6iifXHz//zfz///f8AmCMQS/tDDwAAAABJRU5ErkJggg=="}
]}</content></body><script>
var SLIDES='<div class="slides">{0}</div>';var SLIDE_STYLE="background: {1}, {0};";var SLIDE='<div class="slide slide-{2}" style=\'{1}\'>{0}</div>';var TEXT_STYLE="color: {0}; font-family: {1}; font-size: {2}px; {3}; justify-content: {4}; text-align: {5}; font-weight: {6}";var TEXT_ITEM='<text-item class="canvas-item" style="{1}"><span>{0}</span></text-item>';var COLOR_STYLE="background: {0}; {1}";var COLOR_ITEM='<color-item class="canvas-item" style="{0}"></color-item>';var IMAGE_STYLE="background: url(data:image/{1};base64,{0}) no-repeat center; background-size: contain; {2}";var IMAGE_ITEM='<image-item class="canvas-item" style="{0}"></image-item>';var POSITION_STYLE="left: {0}px; top: {1}px; min-width: {2}px; max-width: {2}px; min-height: {3}px; max-height: {3}px;";function setAspectRatio(aspectRatio){switch(aspectRatio){case 1:SCREEN_W=1920;SCREEN_H=1440;X_OFFSET=280;Y_OFFSET=20;MAX_WIDTH=1800+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=4.8;break;case 2:SCREEN_W=1920;SCREEN_H=1080;X_OFFSET=631;Y_OFFSET=20;MAX_WIDTH=2150+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET;SLIDE_RATIO="16-9"
FONT_SCALE=3.8;break;case 3:SCREEN_W=1920;SCREEN_H=1200;X_OFFSET=540;Y_OFFSET=12;MAX_WIDTH=2065+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET
SLIDE_RATIO="16-10"
FONT_SCALE=3.9;break;case 4:SCREEN_W=1920;SCREEN_H=1280;X_OFFSET=400;Y_OFFSET=20;MAX_WIDTH=1920+X_OFFSET;MAX_HEIGHT=1350+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=4.4;break;case 5:SCREEN_W=2100;SCREEN_H=1280;X_OFFSET=210;Y_OFFSET=20;MAX_WIDTH=1920+X_OFFSET;MAX_HEIGHT=1350+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=5.2;break}}
function getPosition(item){var w_scale=SCREEN_W/MAX_WIDTH;var h_scale=SCREEN_H/MAX_HEIGHT;var x=(item.x+X_OFFSET)*w_scale;var y=(item.y+Y_OFFSET)*h_scale;var w=item.w*w_scale;var h=item.h*h_scale;return String.build(POSITION_STYLE,x,y,w,h)}
function renderSlides(file){let root_object=JSON.parse(file);let content="";for(var id in root_object.slides){setAspectRatio(root_object["aspect-ratio"]);let slide=root_object.slides[id];let slide_content="";for(var object_id in slide.items){let item=slide.items[object_id];var pos=getPosition(item);let style="";switch(item.type){case "text":let text=base64Decode(item['text-data']);let justification;let text_align="";switch(item.justification){case 0:justification="flex-start";text_align="left";break;case 1:justification="center";text_align="center";break;case 2:justification="flex-end";text_align="right";break;case 3:justification="center";text_align="justify";break}
let font_style=item["font-style"];if(font_style.indexOf("italic")!=-1){font_style=font_style.replace(" italic","")}
switch(font_style){case "black":font_style="900";break;case "extrabold":font_style="800";break;case "semibold":font_style="600";break;case "bold":font_style="700";break;case "medium":font_style="500";break;case "regular":font_style="400";break;case "extralight":font_style="300";break;case "light":font_style="200";break;case "thin":font_style="100";break}
style=String.build(TEXT_STYLE,item.color,item.font,item["font-size"]*FONT_SCALE,pos,justification,text_align,font_style);slide_content+=String.build(TEXT_ITEM,text,style);break;case "color":style=String.build(COLOR_STYLE,item.background_color,pos);slide_content+=String.build(COLOR_ITEM,style);break
case "image":style=String.build(IMAGE_STYLE,item["image-data"],item.image,pos);slide_content+=String.build(IMAGE_ITEM,style);break}}
let background_pattern=slide["background-pattern"];if(background_pattern!==""){let pattern=background_pattern.split("/");background_pattern="url(https://raw.githubusercontent.com/Philip-Scott/Spice-up/master/data/assets/patterns/"+pattern[pattern.length-1]+")"}else{background_pattern="none"}
let style=String.build(SLIDE_STYLE,slide["background-color"],background_pattern);content+=String.build(SLIDE,slide_content,style,SLIDE_RATIO);get('body').innerHTML=String.build(SLIDES,content)}}
renderSlides(get('content').innerHTML)
</script></html>
